.subckt aon21bv0x4 a1 a2 b vdd vss z
*   SPICE3 file   created from aon21bv0x4.ext -      technology: scmos
m00 z      an     vdd    vdd p w=26u  l=2.3636u ad=104p     pd=34.6667u as=138.775p ps=49.4u
m01 vdd    b      z      vdd p w=26u  l=2.3636u ad=138.775p pd=49.4u    as=104p     ps=34.6667u
m02 z      b      vdd    vdd p w=22u  l=2.3636u ad=88p      pd=29.3333u as=117.425p ps=41.8u
m03 vdd    an     z      vdd p w=22u  l=2.3636u ad=117.425p pd=41.8u    as=88p      ps=29.3333u
m04 an     a1     vdd    vdd p w=17u  l=2.3636u ad=68p      pd=25.5u    as=90.7375p ps=32.3u
m05 vdd    a2     an     vdd p w=17u  l=2.3636u ad=90.7375p pd=32.3u    as=68p      ps=25.5u
m06 an     a2     vdd    vdd p w=15u  l=2.3636u ad=60p      pd=22.5u    as=80.0625p ps=28.5u
m07 vdd    a1     an     vdd p w=15u  l=2.3636u ad=80.0625p pd=28.5u    as=60p      ps=22.5u
m08 w1     an     vss    vss n w=20u  l=2.3636u ad=50p      pd=25u      as=173.333p ps=52.7273u
m09 z      b      w1     vss n w=20u  l=2.3636u ad=80p      pd=28u      as=50p      ps=25u
m10 w2     b      z      vss n w=20u  l=2.3636u ad=50p      pd=25u      as=80p      ps=28u
m11 vss    an     w2     vss n w=20u  l=2.3636u ad=173.333p pd=52.7273u as=50p      ps=25u
m12 w3     a1     vss    vss n w=15u  l=2.3636u ad=37.5p    pd=20u      as=130p     ps=39.5455u
m13 an     a2     w3     vss n w=15u  l=2.3636u ad=62.3077p pd=26.5385u as=37.5p    ps=20u
m14 w4     a2     an     vss n w=11u  l=2.3636u ad=27.5p    pd=16u      as=45.6923p ps=19.4615u
m15 vss    a1     w4     vss n w=11u  l=2.3636u ad=95.3333p pd=29u      as=27.5p    ps=16u
C0  a1     vdd    0.096f
C1  b      an     0.293f
C2  w1     z      0.010f
C3  an     vdd    0.381f
C4  w3     an     0.016f
C5  vss    a2     0.200f
C6  z      a1     0.003f
C7  vss    b      0.024f
C8  w1     an     0.007f
C9  vss    vdd    0.011f
C10 z      an     0.391f
C11 a2     b      0.024f
C12 a2     vdd    0.027f
C13 a1     an     0.477f
C14 w1     vss    0.005f
C15 b      vdd    0.042f
C16 vss    z      0.200f
C17 vss    a1     0.052f
C18 w2     an     0.007f
C19 a2     a1     0.325f
C20 vss    an     0.267f
C21 z      b      0.169f
C22 a2     an     0.156f
C23 z      vdd    0.463f
C24 a1     b      0.034f
C25 w4     a2     0.011f
C26 w2     vss    0.005f
C28 z      vss    0.008f
C29 a2     vss    0.039f
C30 a1     vss    0.050f
C31 b      vss    0.034f
C32 an     vss    0.047f
.ends
