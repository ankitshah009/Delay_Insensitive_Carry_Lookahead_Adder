magic
tech scmos
timestamp 1185038952
<< checkpaint >>
rect -22 -24 222 124
<< ab >>
rect 0 0 200 100
<< pwell >>
rect -2 -4 202 49
<< nwell >>
rect -2 49 202 104
<< polysilicon >>
rect 81 95 83 98
rect 93 95 95 98
rect 11 83 13 86
rect 23 83 25 86
rect 35 83 37 86
rect 47 83 49 86
rect 57 83 59 86
rect 11 43 13 65
rect 23 43 25 65
rect 35 53 37 65
rect 7 42 13 43
rect 7 38 8 42
rect 12 38 13 42
rect 7 37 13 38
rect 17 42 25 43
rect 17 38 18 42
rect 22 38 25 42
rect 17 37 25 38
rect 33 52 43 53
rect 33 48 38 52
rect 42 48 43 52
rect 33 47 43 48
rect 11 27 13 37
rect 21 29 23 37
rect 33 25 35 47
rect 47 43 49 57
rect 57 53 59 57
rect 121 83 123 86
rect 133 83 135 86
rect 143 83 145 86
rect 155 83 157 86
rect 81 53 83 55
rect 57 52 63 53
rect 57 48 58 52
rect 62 48 63 52
rect 57 47 63 48
rect 81 52 89 53
rect 81 48 84 52
rect 88 48 89 52
rect 81 47 89 48
rect 47 42 53 43
rect 47 39 48 42
rect 45 38 48 39
rect 52 38 53 42
rect 45 37 53 38
rect 45 25 47 37
rect 57 25 59 47
rect 81 25 83 47
rect 93 41 95 55
rect 121 43 123 69
rect 133 67 135 69
rect 143 67 145 69
rect 131 65 135 67
rect 141 65 145 67
rect 167 79 169 82
rect 177 79 179 82
rect 187 79 189 82
rect 131 43 133 65
rect 141 43 143 65
rect 155 63 157 65
rect 153 61 157 63
rect 153 43 155 61
rect 167 53 169 65
rect 177 53 179 65
rect 167 52 173 53
rect 167 49 168 52
rect 107 42 113 43
rect 107 41 108 42
rect 93 39 108 41
rect 93 25 95 39
rect 107 38 108 39
rect 112 38 113 42
rect 107 37 113 38
rect 117 42 123 43
rect 117 38 118 42
rect 122 38 123 42
rect 117 37 123 38
rect 127 42 133 43
rect 127 38 128 42
rect 132 38 133 42
rect 127 37 133 38
rect 137 42 143 43
rect 137 38 138 42
rect 142 38 143 42
rect 137 37 143 38
rect 147 42 155 43
rect 147 38 148 42
rect 152 38 155 42
rect 147 37 155 38
rect 121 25 123 37
rect 131 25 133 37
rect 141 25 143 37
rect 153 27 155 37
rect 165 48 168 49
rect 172 48 173 52
rect 165 47 173 48
rect 177 52 183 53
rect 177 48 178 52
rect 182 48 183 52
rect 177 47 183 48
rect 11 14 13 17
rect 21 14 23 17
rect 33 14 35 17
rect 45 14 47 17
rect 57 14 59 17
rect 165 25 167 47
rect 177 29 179 47
rect 175 27 179 29
rect 187 43 189 65
rect 187 42 193 43
rect 187 38 188 42
rect 192 38 193 42
rect 187 37 193 38
rect 175 25 177 27
rect 187 25 189 37
rect 121 14 123 17
rect 131 14 133 17
rect 141 14 143 17
rect 153 14 155 17
rect 165 14 167 17
rect 175 14 177 17
rect 187 14 189 17
rect 81 2 83 5
rect 93 2 95 5
<< ndiffusion >>
rect 17 27 21 29
rect 3 17 11 27
rect 13 17 21 27
rect 23 25 31 29
rect 149 25 153 27
rect 23 22 33 25
rect 23 18 26 22
rect 30 18 33 22
rect 23 17 33 18
rect 35 22 45 25
rect 35 18 38 22
rect 42 18 45 22
rect 35 17 45 18
rect 47 17 57 25
rect 59 22 67 25
rect 59 18 62 22
rect 66 18 67 22
rect 59 17 67 18
rect 73 22 81 25
rect 73 18 74 22
rect 78 18 81 22
rect 3 12 9 17
rect 3 8 4 12
rect 8 8 9 12
rect 49 12 55 17
rect 3 7 9 8
rect 49 8 50 12
rect 54 8 55 12
rect 49 7 55 8
rect 73 5 81 18
rect 83 12 93 25
rect 83 8 86 12
rect 90 8 93 12
rect 83 5 93 8
rect 95 22 103 25
rect 95 18 98 22
rect 102 18 103 22
rect 95 5 103 18
rect 113 17 121 25
rect 123 17 131 25
rect 133 17 141 25
rect 143 22 153 25
rect 143 18 146 22
rect 150 18 153 22
rect 143 17 153 18
rect 155 25 159 27
rect 155 22 165 25
rect 155 18 158 22
rect 162 18 165 22
rect 155 17 165 18
rect 167 17 175 25
rect 177 22 187 25
rect 177 18 180 22
rect 184 18 187 22
rect 177 17 187 18
rect 189 22 197 25
rect 189 18 192 22
rect 196 18 197 22
rect 189 17 197 18
rect 113 12 119 17
rect 113 8 114 12
rect 118 8 119 12
rect 169 11 173 17
rect 113 7 119 8
rect 168 10 174 11
rect 168 6 169 10
rect 173 6 174 10
rect 168 5 174 6
<< pdiffusion >>
rect 15 92 21 93
rect 15 88 16 92
rect 20 88 21 92
rect 15 83 21 88
rect 3 82 11 83
rect 3 78 4 82
rect 8 78 11 82
rect 3 65 11 78
rect 13 65 23 83
rect 25 82 35 83
rect 25 78 28 82
rect 32 78 35 82
rect 25 65 35 78
rect 37 72 47 83
rect 37 68 40 72
rect 44 68 47 72
rect 37 65 47 68
rect 40 57 47 65
rect 49 57 57 83
rect 59 82 67 83
rect 59 78 62 82
rect 66 78 67 82
rect 59 57 67 78
rect 73 62 81 95
rect 73 58 74 62
rect 78 58 81 62
rect 73 55 81 58
rect 83 92 93 95
rect 83 88 86 92
rect 90 88 93 92
rect 83 55 93 88
rect 95 72 103 95
rect 136 94 142 95
rect 95 68 98 72
rect 102 68 103 72
rect 110 92 118 93
rect 110 88 112 92
rect 116 88 118 92
rect 136 90 137 94
rect 141 90 142 94
rect 136 89 142 90
rect 110 83 118 88
rect 137 83 141 89
rect 110 69 121 83
rect 123 82 133 83
rect 123 78 126 82
rect 130 78 133 82
rect 123 69 133 78
rect 135 69 143 83
rect 145 82 155 83
rect 145 78 148 82
rect 152 78 155 82
rect 145 69 155 78
rect 95 62 103 68
rect 95 58 98 62
rect 102 58 103 62
rect 95 55 103 58
rect 147 65 155 69
rect 157 79 164 83
rect 191 82 197 83
rect 191 79 192 82
rect 157 72 167 79
rect 157 68 160 72
rect 164 68 167 72
rect 157 65 167 68
rect 169 65 177 79
rect 179 65 187 79
rect 189 78 192 79
rect 196 78 197 82
rect 189 65 197 78
<< metal1 >>
rect -2 96 202 101
rect -2 92 30 96
rect 34 92 38 96
rect 42 92 46 96
rect 50 92 54 96
rect 58 92 62 96
rect 66 94 150 96
rect 66 92 137 94
rect -2 88 16 92
rect 20 88 86 92
rect 90 88 112 92
rect 116 90 137 92
rect 141 92 150 94
rect 154 92 158 96
rect 162 92 166 96
rect 170 92 174 96
rect 178 92 182 96
rect 186 92 202 96
rect 141 90 202 92
rect 116 88 202 90
rect -2 87 202 88
rect 3 82 9 83
rect 27 82 33 83
rect 61 82 67 83
rect 125 82 131 83
rect 147 82 153 83
rect 191 82 197 83
rect 3 78 4 82
rect 8 78 28 82
rect 32 78 62 82
rect 66 78 67 82
rect 3 77 9 78
rect 27 77 33 78
rect 61 77 67 78
rect 86 78 114 82
rect 39 72 45 73
rect 86 72 90 78
rect 7 42 13 72
rect 7 38 8 42
rect 12 38 13 42
rect 7 18 13 38
rect 17 42 23 72
rect 17 38 18 42
rect 22 38 23 42
rect 17 28 23 38
rect 28 68 40 72
rect 44 68 90 72
rect 28 23 32 68
rect 39 67 45 68
rect 67 62 79 63
rect 37 52 43 62
rect 37 48 38 52
rect 42 48 43 52
rect 37 28 43 48
rect 47 42 53 62
rect 47 38 48 42
rect 52 38 53 42
rect 47 28 53 38
rect 57 52 63 62
rect 57 48 58 52
rect 62 48 63 52
rect 57 28 63 48
rect 67 58 74 62
rect 78 58 79 62
rect 67 57 79 58
rect 67 33 73 57
rect 86 53 90 68
rect 83 52 90 53
rect 83 48 84 52
rect 88 48 90 52
rect 97 72 103 73
rect 97 68 98 72
rect 102 68 103 72
rect 110 72 114 78
rect 125 78 126 82
rect 130 78 148 82
rect 152 78 192 82
rect 196 78 197 82
rect 125 77 131 78
rect 147 77 153 78
rect 191 77 197 78
rect 158 72 165 73
rect 110 68 152 72
rect 97 62 103 68
rect 97 58 98 62
rect 102 58 103 62
rect 83 47 89 48
rect 67 27 83 33
rect 77 23 83 27
rect 25 22 32 23
rect 25 18 26 22
rect 30 18 32 22
rect 37 22 43 23
rect 61 22 67 23
rect 37 18 38 22
rect 42 18 62 22
rect 66 18 67 22
rect 25 17 31 18
rect 37 17 43 18
rect 61 17 67 18
rect 73 22 83 23
rect 73 18 74 22
rect 78 18 83 22
rect 97 22 103 58
rect 107 42 113 43
rect 107 38 108 42
rect 112 38 113 42
rect 107 37 113 38
rect 117 42 123 62
rect 117 38 118 42
rect 122 38 123 42
rect 97 18 98 22
rect 102 18 103 22
rect 108 22 112 37
rect 117 28 123 38
rect 127 42 133 62
rect 127 38 128 42
rect 132 38 133 42
rect 127 28 133 38
rect 137 42 143 62
rect 148 43 152 68
rect 158 68 160 72
rect 164 68 165 72
rect 158 67 165 68
rect 137 38 138 42
rect 142 38 143 42
rect 137 28 143 38
rect 147 42 153 43
rect 147 38 148 42
rect 152 38 153 42
rect 147 37 153 38
rect 158 32 162 67
rect 148 28 162 32
rect 167 52 173 62
rect 167 48 168 52
rect 172 48 173 52
rect 167 28 173 48
rect 177 52 183 72
rect 177 48 178 52
rect 182 48 183 52
rect 177 28 183 48
rect 187 42 193 72
rect 187 38 188 42
rect 192 38 193 42
rect 187 28 193 38
rect 148 23 152 28
rect 145 22 152 23
rect 108 18 146 22
rect 150 18 152 22
rect 73 17 82 18
rect 97 17 103 18
rect 145 17 152 18
rect 157 22 163 23
rect 179 22 185 23
rect 157 18 158 22
rect 162 18 180 22
rect 184 18 185 22
rect 157 17 163 18
rect 179 17 185 18
rect 191 22 197 23
rect 191 18 192 22
rect 196 18 197 22
rect 191 13 197 18
rect -2 12 202 13
rect -2 8 4 12
rect 8 10 50 12
rect 8 8 18 10
rect -2 6 18 8
rect 22 6 28 10
rect 32 6 38 10
rect 42 8 50 10
rect 54 8 86 12
rect 90 8 114 12
rect 118 10 202 12
rect 118 8 126 10
rect 42 6 126 8
rect 130 6 136 10
rect 140 6 146 10
rect 150 6 157 10
rect 161 6 169 10
rect 173 6 182 10
rect 186 6 190 10
rect 194 6 202 10
rect -2 -1 202 6
<< ntransistor >>
rect 11 17 13 27
rect 21 17 23 29
rect 33 17 35 25
rect 45 17 47 25
rect 57 17 59 25
rect 81 5 83 25
rect 93 5 95 25
rect 121 17 123 25
rect 131 17 133 25
rect 141 17 143 25
rect 153 17 155 27
rect 165 17 167 25
rect 175 17 177 25
rect 187 17 189 25
<< ptransistor >>
rect 11 65 13 83
rect 23 65 25 83
rect 35 65 37 83
rect 47 57 49 83
rect 57 57 59 83
rect 81 55 83 95
rect 93 55 95 95
rect 121 69 123 83
rect 133 69 135 83
rect 143 69 145 83
rect 155 65 157 83
rect 167 65 169 79
rect 177 65 179 79
rect 187 65 189 79
<< polycontact >>
rect 8 38 12 42
rect 18 38 22 42
rect 38 48 42 52
rect 58 48 62 52
rect 84 48 88 52
rect 48 38 52 42
rect 108 38 112 42
rect 118 38 122 42
rect 128 38 132 42
rect 138 38 142 42
rect 148 38 152 42
rect 168 48 172 52
rect 178 48 182 52
rect 188 38 192 42
<< ndcontact >>
rect 26 18 30 22
rect 38 18 42 22
rect 62 18 66 22
rect 74 18 78 22
rect 4 8 8 12
rect 50 8 54 12
rect 86 8 90 12
rect 98 18 102 22
rect 146 18 150 22
rect 158 18 162 22
rect 180 18 184 22
rect 192 18 196 22
rect 114 8 118 12
rect 169 6 173 10
<< pdcontact >>
rect 16 88 20 92
rect 4 78 8 82
rect 28 78 32 82
rect 40 68 44 72
rect 62 78 66 82
rect 74 58 78 62
rect 86 88 90 92
rect 98 68 102 72
rect 112 88 116 92
rect 137 90 141 94
rect 126 78 130 82
rect 148 78 152 82
rect 98 58 102 62
rect 160 68 164 72
rect 192 78 196 82
<< psubstratepcontact >>
rect 18 6 22 10
rect 28 6 32 10
rect 38 6 42 10
rect 126 6 130 10
rect 136 6 140 10
rect 146 6 150 10
rect 157 6 161 10
rect 182 6 186 10
rect 190 6 194 10
<< nsubstratencontact >>
rect 30 92 34 96
rect 38 92 42 96
rect 46 92 50 96
rect 54 92 58 96
rect 62 92 66 96
rect 150 92 154 96
rect 158 92 162 96
rect 166 92 170 96
rect 174 92 178 96
rect 182 92 186 96
<< psubstratepdiff >>
rect 17 10 43 11
rect 17 6 18 10
rect 22 6 28 10
rect 32 6 38 10
rect 42 6 43 10
rect 17 5 43 6
rect 125 10 162 11
rect 125 6 126 10
rect 130 6 136 10
rect 140 6 146 10
rect 150 6 157 10
rect 161 6 162 10
rect 125 5 162 6
rect 181 10 195 11
rect 181 6 182 10
rect 186 6 190 10
rect 194 6 195 10
rect 181 5 195 6
<< nsubstratendiff >>
rect 29 96 67 97
rect 29 92 30 96
rect 34 92 38 96
rect 42 92 46 96
rect 50 92 54 96
rect 58 92 62 96
rect 66 92 67 96
rect 149 96 187 97
rect 29 91 67 92
rect 149 92 150 96
rect 154 92 158 96
rect 162 92 166 96
rect 170 92 174 96
rect 178 92 182 96
rect 186 92 187 96
rect 149 91 187 92
<< labels >>
rlabel metal1 10 45 10 45 6 a1
rlabel metal1 20 50 20 50 6 b1
rlabel metal1 20 50 20 50 6 b1
rlabel metal1 10 45 10 45 6 a1
rlabel metal1 40 45 40 45 6 cin1
rlabel metal1 40 45 40 45 6 cin1
rlabel metal1 70 45 70 45 6 cout
rlabel metal1 60 45 60 45 6 b2
rlabel metal1 50 45 50 45 6 a2
rlabel metal1 70 45 70 45 6 cout
rlabel metal1 50 45 50 45 6 a2
rlabel metal1 60 45 60 45 6 b2
rlabel metal1 100 6 100 6 6 vss
rlabel metal1 100 6 100 6 6 vss
rlabel metal1 80 25 80 25 6 cout
rlabel metal1 80 25 80 25 6 cout
rlabel metal1 100 45 100 45 6 sout
rlabel metal1 100 45 100 45 6 sout
rlabel metal1 100 94 100 94 6 vdd
rlabel metal1 100 94 100 94 6 vdd
rlabel metal1 120 45 120 45 6 a3
rlabel metal1 120 45 120 45 6 a3
rlabel metal1 140 45 140 45 6 cin2
rlabel metal1 130 45 130 45 6 b3
rlabel metal1 140 45 140 45 6 cin2
rlabel metal1 130 45 130 45 6 b3
rlabel polycontact 180 50 180 50 6 a4
rlabel metal1 190 50 190 50 6 b4
rlabel metal1 170 45 170 45 6 cin3
rlabel metal1 190 50 190 50 6 b4
rlabel polycontact 180 50 180 50 6 a4
rlabel metal1 170 45 170 45 6 cin3
<< end >>
