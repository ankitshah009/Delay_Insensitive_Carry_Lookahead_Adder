magic
tech scmos
timestamp 1179387376
<< checkpaint >>
rect -22 -25 70 105
<< ab >>
rect 0 0 48 80
<< pwell >>
rect -4 -7 52 36
<< nwell >>
rect -4 36 52 87
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect -2 68 50 78
rect -2 2 50 12
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
<< psubstratepdiff >>
rect 0 2 48 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 48 2
rect 0 -3 48 -2
<< nsubstratendiff >>
rect 0 82 48 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 48 82
rect 0 77 48 78
<< labels >>
rlabel metal1 24 6 24 6 6 vss
rlabel metal1 24 74 24 74 6 vdd
<< end >>
