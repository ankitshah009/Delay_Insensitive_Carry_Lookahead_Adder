magic
tech scmos
timestamp 1179385235
<< checkpaint >>
rect -22 -25 94 105
<< ab >>
rect 0 0 72 80
<< pwell >>
rect -4 -7 76 36
<< nwell >>
rect -4 36 76 87
<< polysilicon >>
rect 9 63 11 68
rect 21 63 23 68
rect 41 63 43 68
rect 51 63 53 68
rect 61 63 63 68
rect 9 48 11 51
rect 9 47 15 48
rect 9 43 10 47
rect 14 43 15 47
rect 9 42 15 43
rect 9 22 11 42
rect 21 38 23 51
rect 41 39 43 47
rect 51 39 53 47
rect 61 44 63 47
rect 60 43 70 44
rect 60 39 65 43
rect 69 39 70 43
rect 33 38 43 39
rect 16 37 24 38
rect 16 33 17 37
rect 21 33 24 37
rect 33 34 34 38
rect 38 35 43 38
rect 49 38 55 39
rect 38 34 45 35
rect 33 33 45 34
rect 49 34 50 38
rect 54 34 55 38
rect 49 33 55 34
rect 16 32 24 33
rect 22 29 24 32
rect 43 30 45 33
rect 53 30 55 33
rect 60 38 70 39
rect 60 30 62 38
rect 22 18 24 23
rect 9 11 11 16
rect 43 19 45 24
rect 53 18 55 23
rect 60 18 62 23
<< ndiffusion >>
rect 13 23 22 29
rect 24 28 31 29
rect 24 24 26 28
rect 30 24 31 28
rect 24 23 31 24
rect 35 24 43 30
rect 45 29 53 30
rect 45 25 47 29
rect 51 25 53 29
rect 45 24 53 25
rect 13 22 20 23
rect 2 21 9 22
rect 2 17 3 21
rect 7 17 9 21
rect 2 16 9 17
rect 11 16 20 22
rect 13 12 20 16
rect 13 8 14 12
rect 18 8 20 12
rect 13 7 20 8
rect 35 12 41 24
rect 48 23 53 24
rect 55 23 60 30
rect 62 28 69 30
rect 62 24 64 28
rect 68 24 69 28
rect 62 23 69 24
rect 35 8 36 12
rect 40 8 41 12
rect 35 7 41 8
<< pdiffusion >>
rect 13 72 19 73
rect 13 68 14 72
rect 18 68 19 72
rect 13 63 19 68
rect 4 57 9 63
rect 2 56 9 57
rect 2 52 3 56
rect 7 52 9 56
rect 2 51 9 52
rect 11 51 21 63
rect 23 57 28 63
rect 23 56 30 57
rect 23 52 25 56
rect 29 52 30 56
rect 36 53 41 63
rect 23 51 30 52
rect 34 52 41 53
rect 34 48 35 52
rect 39 48 41 52
rect 34 47 41 48
rect 43 62 51 63
rect 43 58 45 62
rect 49 58 51 62
rect 43 55 51 58
rect 43 51 45 55
rect 49 51 51 55
rect 43 47 51 51
rect 53 62 61 63
rect 53 58 55 62
rect 59 58 61 62
rect 53 47 61 58
rect 63 62 70 63
rect 63 58 65 62
rect 69 58 70 62
rect 63 55 70 58
rect 63 51 65 55
rect 69 51 70 55
rect 63 50 70 51
rect 63 47 68 50
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect -2 72 74 78
rect -2 68 14 72
rect 18 68 74 72
rect 10 57 22 63
rect 54 62 60 68
rect 44 58 45 62
rect 49 58 50 62
rect 54 58 55 62
rect 59 58 60 62
rect 64 58 65 62
rect 69 58 70 62
rect 2 56 7 57
rect 2 52 3 56
rect 2 51 7 52
rect 2 21 6 51
rect 10 47 14 57
rect 25 56 29 57
rect 10 41 14 43
rect 18 37 22 47
rect 10 33 17 37
rect 21 33 22 37
rect 25 38 29 52
rect 34 52 39 56
rect 34 48 35 52
rect 44 55 50 58
rect 64 55 70 58
rect 44 51 45 55
rect 49 51 65 55
rect 69 51 70 55
rect 34 47 39 48
rect 34 43 46 47
rect 25 34 34 38
rect 38 34 39 38
rect 10 25 14 33
rect 25 28 31 34
rect 25 24 26 28
rect 30 24 31 28
rect 42 29 46 43
rect 57 43 70 47
rect 57 42 65 43
rect 69 39 70 43
rect 49 34 50 38
rect 54 34 60 38
rect 42 25 47 29
rect 51 25 52 29
rect 56 21 60 34
rect 65 33 70 39
rect 2 17 3 21
rect 7 17 60 21
rect 64 28 68 29
rect 64 12 68 24
rect -2 8 14 12
rect 18 8 36 12
rect 40 8 74 12
rect -2 2 74 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
<< ntransistor >>
rect 22 23 24 29
rect 43 24 45 30
rect 9 16 11 22
rect 53 23 55 30
rect 60 23 62 30
<< ptransistor >>
rect 9 51 11 63
rect 21 51 23 63
rect 41 47 43 63
rect 51 47 53 63
rect 61 47 63 63
<< polycontact >>
rect 10 43 14 47
rect 65 39 69 43
rect 17 33 21 37
rect 34 34 38 38
rect 50 34 54 38
<< ndcontact >>
rect 26 24 30 28
rect 47 25 51 29
rect 3 17 7 21
rect 14 8 18 12
rect 64 24 68 28
rect 36 8 40 12
<< pdcontact >>
rect 14 68 18 72
rect 3 52 7 56
rect 25 52 29 56
rect 35 48 39 52
rect 45 58 49 62
rect 45 51 49 55
rect 55 58 59 62
rect 65 58 69 62
rect 65 51 69 55
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
<< psubstratepdiff >>
rect 0 2 72 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 72 2
rect 0 -3 72 -2
<< nsubstratendiff >>
rect 0 82 72 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 72 82
rect 0 77 72 78
<< labels >>
rlabel polysilicon 38 36 38 36 6 bn
rlabel polycontact 52 36 52 36 6 a2n
rlabel pdcontact 4 54 4 54 6 a2n
rlabel metal1 12 28 12 28 6 b
rlabel metal1 20 40 20 40 6 b
rlabel metal1 12 52 12 52 6 a2
rlabel metal1 20 60 20 60 6 a2
rlabel metal1 36 6 36 6 6 vss
rlabel metal1 32 36 32 36 6 bn
rlabel metal1 36 52 36 52 6 z
rlabel metal1 27 40 27 40 6 bn
rlabel metal1 36 74 36 74 6 vdd
rlabel metal1 44 36 44 36 6 z
rlabel metal1 47 56 47 56 6 n1
rlabel metal1 31 19 31 19 6 a2n
rlabel metal1 60 44 60 44 6 a1
rlabel metal1 54 36 54 36 6 a2n
rlabel polycontact 68 40 68 40 6 a1
rlabel metal1 57 53 57 53 6 n1
rlabel metal1 67 56 67 56 6 n1
<< end >>
