magic
tech scmos
timestamp 1179387811
<< checkpaint >>
rect -22 -25 150 105
<< ab >>
rect 0 0 128 80
<< pwell >>
rect -4 -7 132 36
<< nwell >>
rect -4 36 132 87
<< polysilicon >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 39 70 41 74
rect 49 70 51 74
rect 69 70 71 74
rect 79 70 81 74
rect 89 70 91 74
rect 39 53 41 56
rect 49 53 51 56
rect 39 52 51 53
rect 39 51 46 52
rect 45 48 46 51
rect 50 48 51 52
rect 45 47 51 48
rect 100 64 116 65
rect 100 63 111 64
rect 100 60 102 63
rect 110 60 111 63
rect 115 60 116 64
rect 110 59 116 60
rect 110 56 112 59
rect 100 42 102 46
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 69 39 71 42
rect 79 39 81 42
rect 9 38 15 39
rect 9 34 10 38
rect 14 34 15 38
rect 9 33 15 34
rect 19 38 25 39
rect 19 34 20 38
rect 24 34 25 38
rect 29 38 65 39
rect 29 37 60 38
rect 19 33 25 34
rect 10 24 12 33
rect 19 29 21 33
rect 37 29 39 37
rect 59 34 60 37
rect 64 34 65 38
rect 59 33 65 34
rect 69 38 75 39
rect 69 34 70 38
rect 74 34 75 38
rect 69 33 75 34
rect 79 38 85 39
rect 79 34 80 38
rect 84 34 85 38
rect 89 38 91 42
rect 89 37 103 38
rect 89 36 98 37
rect 79 33 85 34
rect 97 33 98 36
rect 102 33 103 37
rect 49 32 55 33
rect 17 27 21 29
rect 17 24 19 27
rect 27 24 29 29
rect 49 28 50 32
rect 54 28 55 32
rect 49 27 55 28
rect 49 24 51 27
rect 72 24 74 33
rect 79 24 81 33
rect 97 32 103 33
rect 99 29 101 32
rect 110 30 112 42
rect 89 24 91 29
rect 37 12 39 16
rect 10 6 12 11
rect 17 6 19 11
rect 27 8 29 11
rect 49 8 51 13
rect 27 6 51 8
rect 99 12 101 16
rect 72 6 74 11
rect 79 6 81 11
rect 89 8 91 11
rect 110 8 112 19
rect 89 6 112 8
<< ndiffusion >>
rect 32 24 37 29
rect 2 12 10 24
rect 2 8 3 12
rect 7 11 10 12
rect 12 11 17 24
rect 19 22 27 24
rect 19 18 21 22
rect 25 18 27 22
rect 19 11 27 18
rect 29 23 37 24
rect 29 19 31 23
rect 35 19 37 23
rect 29 16 37 19
rect 39 24 47 29
rect 105 29 110 30
rect 94 24 99 29
rect 39 16 49 24
rect 29 11 34 16
rect 41 15 49 16
rect 41 11 42 15
rect 46 13 49 15
rect 51 23 58 24
rect 51 19 53 23
rect 57 19 58 23
rect 51 18 58 19
rect 51 13 56 18
rect 46 11 47 13
rect 7 8 8 11
rect 2 7 8 8
rect 41 10 47 11
rect 64 12 72 24
rect 64 8 65 12
rect 69 11 72 12
rect 74 11 79 24
rect 81 22 89 24
rect 81 18 83 22
rect 87 18 89 22
rect 81 11 89 18
rect 91 23 99 24
rect 91 19 93 23
rect 97 19 99 23
rect 91 16 99 19
rect 101 21 110 29
rect 101 17 103 21
rect 107 19 110 21
rect 112 29 119 30
rect 112 25 114 29
rect 118 25 119 29
rect 112 24 119 25
rect 112 19 117 24
rect 107 17 108 19
rect 101 16 108 17
rect 91 11 96 16
rect 69 8 70 11
rect 64 7 70 8
<< pdiffusion >>
rect 116 72 122 73
rect 4 63 9 70
rect 2 62 9 63
rect 2 58 3 62
rect 7 58 9 62
rect 2 57 9 58
rect 4 42 9 57
rect 11 54 19 70
rect 11 50 13 54
rect 17 50 19 54
rect 11 42 19 50
rect 21 54 29 70
rect 21 50 23 54
rect 27 50 29 54
rect 21 47 29 50
rect 21 43 23 47
rect 27 43 29 47
rect 21 42 29 43
rect 31 69 39 70
rect 31 65 33 69
rect 37 65 39 69
rect 31 56 39 65
rect 41 62 49 70
rect 41 58 43 62
rect 47 58 49 62
rect 41 56 49 58
rect 51 69 58 70
rect 51 65 53 69
rect 57 65 58 69
rect 51 62 58 65
rect 64 63 69 70
rect 51 58 53 62
rect 57 58 58 62
rect 51 56 58 58
rect 62 62 69 63
rect 62 58 63 62
rect 67 58 69 62
rect 62 57 69 58
rect 31 42 37 56
rect 64 42 69 57
rect 71 54 79 70
rect 71 50 73 54
rect 77 50 79 54
rect 71 42 79 50
rect 81 54 89 70
rect 81 50 83 54
rect 87 50 89 54
rect 81 47 89 50
rect 81 43 83 47
rect 87 43 89 47
rect 81 42 89 43
rect 91 69 98 70
rect 91 65 93 69
rect 97 65 98 69
rect 116 68 117 72
rect 121 68 122 72
rect 116 67 122 68
rect 91 60 98 65
rect 91 46 100 60
rect 102 56 107 60
rect 118 56 122 67
rect 102 51 110 56
rect 102 47 104 51
rect 108 47 110 51
rect 102 46 110 47
rect 91 42 98 46
rect 105 42 110 46
rect 112 42 122 56
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect 118 78 122 82
rect 126 78 130 82
rect -2 72 130 78
rect -2 69 117 72
rect -2 68 33 69
rect 32 65 33 68
rect 37 68 53 69
rect 37 65 38 68
rect 52 65 53 68
rect 57 68 93 69
rect 57 65 58 68
rect 92 65 93 68
rect 97 68 117 69
rect 121 68 130 72
rect 97 65 98 68
rect 52 62 58 65
rect 110 63 111 64
rect 2 58 3 62
rect 7 58 43 62
rect 47 58 48 62
rect 52 58 53 62
rect 57 58 58 62
rect 62 58 63 62
rect 67 58 94 62
rect 2 50 13 54
rect 17 50 18 54
rect 22 50 23 54
rect 27 50 28 54
rect 2 22 6 50
rect 22 47 28 50
rect 10 43 23 47
rect 27 43 28 47
rect 10 38 14 43
rect 32 38 36 58
rect 83 54 87 55
rect 41 52 54 54
rect 41 48 46 52
rect 19 34 20 38
rect 24 34 45 38
rect 10 30 14 34
rect 10 26 35 30
rect 31 23 35 26
rect 2 18 21 22
rect 25 18 26 22
rect 41 23 45 34
rect 50 32 54 52
rect 62 50 73 54
rect 77 50 78 54
rect 62 38 66 50
rect 83 47 87 50
rect 59 34 60 38
rect 64 34 66 38
rect 50 27 54 28
rect 41 19 53 23
rect 57 19 58 23
rect 62 22 66 34
rect 70 43 83 46
rect 70 42 87 43
rect 90 46 94 58
rect 106 60 111 63
rect 115 63 116 64
rect 115 60 118 63
rect 106 57 118 60
rect 104 51 108 52
rect 114 49 118 57
rect 104 46 108 47
rect 90 42 118 46
rect 70 38 74 42
rect 90 38 94 42
rect 79 34 80 38
rect 84 34 94 38
rect 98 37 111 39
rect 70 30 74 34
rect 102 33 111 37
rect 70 26 97 30
rect 105 26 111 33
rect 114 29 118 42
rect 93 23 97 26
rect 114 24 118 25
rect 31 18 35 19
rect 62 18 83 22
rect 87 18 88 22
rect 93 18 97 19
rect 103 21 107 22
rect 41 12 42 15
rect -2 8 3 12
rect 7 11 42 12
rect 46 12 47 15
rect 103 12 107 17
rect 46 11 65 12
rect 7 8 65 11
rect 69 8 130 12
rect -2 2 130 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 122 2
rect 126 -2 130 2
<< ntransistor >>
rect 10 11 12 24
rect 17 11 19 24
rect 27 11 29 24
rect 37 16 39 29
rect 49 13 51 24
rect 72 11 74 24
rect 79 11 81 24
rect 89 11 91 24
rect 99 16 101 29
rect 110 19 112 30
<< ptransistor >>
rect 9 42 11 70
rect 19 42 21 70
rect 29 42 31 70
rect 39 56 41 70
rect 49 56 51 70
rect 69 42 71 70
rect 79 42 81 70
rect 89 42 91 70
rect 100 46 102 60
rect 110 42 112 56
<< polycontact >>
rect 46 48 50 52
rect 111 60 115 64
rect 10 34 14 38
rect 20 34 24 38
rect 60 34 64 38
rect 70 34 74 38
rect 80 34 84 38
rect 98 33 102 37
rect 50 28 54 32
<< ndcontact >>
rect 3 8 7 12
rect 21 18 25 22
rect 31 19 35 23
rect 42 11 46 15
rect 53 19 57 23
rect 65 8 69 12
rect 83 18 87 22
rect 93 19 97 23
rect 103 17 107 21
rect 114 25 118 29
<< pdcontact >>
rect 3 58 7 62
rect 13 50 17 54
rect 23 50 27 54
rect 23 43 27 47
rect 33 65 37 69
rect 43 58 47 62
rect 53 65 57 69
rect 53 58 57 62
rect 63 58 67 62
rect 73 50 77 54
rect 83 50 87 54
rect 83 43 87 47
rect 93 65 97 69
rect 117 68 121 72
rect 104 47 108 51
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
rect 90 -2 94 2
rect 98 -2 102 2
rect 106 -2 110 2
rect 114 -2 118 2
rect 122 -2 126 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
rect 90 78 94 82
rect 98 78 102 82
rect 106 78 110 82
rect 114 78 118 82
rect 122 78 126 82
<< psubstratepdiff >>
rect 0 2 128 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 122 2
rect 126 -2 128 2
rect 0 -3 128 -2
<< nsubstratendiff >>
rect 0 82 128 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect 118 78 122 82
rect 126 78 128 82
rect 0 77 128 78
<< labels >>
rlabel polycontact 22 36 22 36 6 cn
rlabel ntransistor 73 22 73 22 6 an
rlabel polycontact 82 36 82 36 6 bn
rlabel metal1 20 20 20 20 6 z
rlabel metal1 12 20 12 20 6 z
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 52 12 52 6 z
rlabel metal1 44 52 44 52 6 c
rlabel metal1 34 48 34 48 6 cn
rlabel metal1 25 60 25 60 6 cn
rlabel metal1 64 6 64 6 6 vss
rlabel metal1 49 21 49 21 6 cn
rlabel polycontact 72 36 72 36 6 an
rlabel metal1 52 40 52 40 6 c
rlabel metal1 64 74 64 74 6 vdd
rlabel metal1 95 24 95 24 6 an
rlabel metal1 86 36 86 36 6 bn
rlabel polycontact 100 36 100 36 6 a
rlabel metal1 85 48 85 48 6 an
rlabel metal1 78 60 78 60 6 bn
rlabel metal1 108 32 108 32 6 a
rlabel metal1 116 35 116 35 6 bn
rlabel metal1 106 47 106 47 6 bn
rlabel metal1 116 56 116 56 6 b
rlabel metal1 108 60 108 60 6 b
<< end >>
