magic
tech scmos
timestamp 1179385105
<< checkpaint >>
rect -22 -22 78 94
<< ab >>
rect 0 0 56 72
<< pwell >>
rect -4 -4 60 32
<< nwell >>
rect -4 32 60 76
<< polysilicon >>
rect 9 66 11 70
rect 19 63 21 68
rect 29 63 31 68
rect 41 63 43 68
rect 19 43 21 54
rect 29 51 31 54
rect 29 50 37 51
rect 29 46 32 50
rect 36 46 37 50
rect 29 45 37 46
rect 19 42 25 43
rect 19 38 20 42
rect 24 38 25 42
rect 9 35 11 38
rect 19 37 25 38
rect 9 34 15 35
rect 9 30 10 34
rect 14 30 15 34
rect 9 29 15 30
rect 9 26 11 29
rect 22 22 24 37
rect 29 22 31 45
rect 41 31 43 54
rect 40 30 46 31
rect 40 27 41 30
rect 36 26 41 27
rect 45 26 46 30
rect 36 25 46 26
rect 36 22 38 25
rect 9 8 11 12
rect 22 8 24 13
rect 29 8 31 13
rect 36 8 38 13
<< ndiffusion >>
rect 4 19 9 26
rect 2 18 9 19
rect 2 14 3 18
rect 7 14 9 18
rect 2 12 9 14
rect 11 22 20 26
rect 11 13 22 22
rect 24 13 29 22
rect 31 13 36 22
rect 38 19 43 22
rect 38 18 45 19
rect 38 14 40 18
rect 44 14 45 18
rect 38 13 45 14
rect 11 12 20 13
rect 13 8 20 12
rect 13 4 14 8
rect 18 4 20 8
rect 13 3 20 4
<< pdiffusion >>
rect 33 68 39 69
rect 4 51 9 66
rect 2 50 9 51
rect 2 46 3 50
rect 7 46 9 50
rect 2 43 9 46
rect 2 39 3 43
rect 7 39 9 43
rect 2 38 9 39
rect 11 63 16 66
rect 33 64 34 68
rect 38 64 39 68
rect 33 63 39 64
rect 11 62 19 63
rect 11 58 13 62
rect 17 58 19 62
rect 11 54 19 58
rect 21 59 29 63
rect 21 55 23 59
rect 27 55 29 59
rect 21 54 29 55
rect 31 54 41 63
rect 43 60 48 63
rect 43 59 50 60
rect 43 55 45 59
rect 49 55 50 59
rect 43 54 50 55
rect 11 38 17 54
<< metal1 >>
rect -2 68 58 72
rect -2 64 34 68
rect 38 64 58 68
rect 13 62 17 64
rect 2 50 7 59
rect 13 57 17 58
rect 22 55 23 59
rect 27 55 45 59
rect 49 55 50 59
rect 22 50 26 55
rect 2 46 3 50
rect 2 43 7 46
rect 2 39 3 43
rect 2 38 7 39
rect 10 46 26 50
rect 31 46 32 50
rect 36 46 47 50
rect 2 18 6 38
rect 10 34 14 46
rect 17 38 20 42
rect 24 38 31 42
rect 41 38 47 46
rect 25 30 31 38
rect 41 30 47 34
rect 10 26 14 30
rect 45 26 47 30
rect 10 22 22 26
rect 25 22 47 26
rect 18 18 22 22
rect 2 14 3 18
rect 7 14 15 18
rect 18 14 40 18
rect 44 14 45 18
rect -2 4 14 8
rect 18 4 58 8
rect -2 0 58 4
<< ntransistor >>
rect 9 12 11 26
rect 22 13 24 22
rect 29 13 31 22
rect 36 13 38 22
<< ptransistor >>
rect 9 38 11 66
rect 19 54 21 63
rect 29 54 31 63
rect 41 54 43 63
<< polycontact >>
rect 32 46 36 50
rect 20 38 24 42
rect 10 30 14 34
rect 41 26 45 30
<< ndcontact >>
rect 3 14 7 18
rect 40 14 44 18
rect 14 4 18 8
<< pdcontact >>
rect 3 46 7 50
rect 3 39 7 43
rect 34 64 38 68
rect 13 58 17 62
rect 23 55 27 59
rect 45 55 49 59
<< labels >>
rlabel polycontact 12 32 12 32 6 zn
rlabel pdcontact 4 40 4 40 6 z
rlabel metal1 12 16 12 16 6 z
rlabel metal1 20 40 20 40 6 a
rlabel metal1 12 36 12 36 6 zn
rlabel metal1 28 4 28 4 6 vss
rlabel metal1 28 24 28 24 6 c
rlabel metal1 36 24 36 24 6 c
rlabel metal1 28 36 28 36 6 a
rlabel metal1 36 48 36 48 6 b
rlabel metal1 28 68 28 68 6 vdd
rlabel metal1 31 16 31 16 6 zn
rlabel polycontact 44 28 44 28 6 c
rlabel metal1 44 44 44 44 6 b
rlabel metal1 36 57 36 57 6 zn
<< end >>
