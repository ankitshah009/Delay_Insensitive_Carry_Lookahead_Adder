magic
tech scmos
timestamp 1179385621
<< checkpaint >>
rect -22 -25 134 105
<< ab >>
rect 0 0 112 80
<< pwell >>
rect -4 -7 116 36
<< nwell >>
rect -4 36 116 87
<< polysilicon >>
rect 25 72 110 74
rect 15 63 17 68
rect 25 64 27 72
rect 56 69 58 72
rect 35 64 37 68
rect 77 64 79 68
rect 87 64 89 72
rect 97 64 99 68
rect 56 44 58 47
rect 56 42 61 44
rect 15 39 17 42
rect 2 38 17 39
rect 2 34 3 38
rect 7 34 17 38
rect 25 39 27 42
rect 25 37 30 39
rect 2 33 17 34
rect 12 26 14 33
rect 28 31 30 37
rect 35 38 37 42
rect 59 40 61 42
rect 59 39 65 40
rect 77 39 79 42
rect 35 37 55 38
rect 35 36 50 37
rect 43 33 50 36
rect 54 33 55 37
rect 43 32 55 33
rect 59 35 60 39
rect 64 35 65 39
rect 59 34 65 35
rect 73 38 79 39
rect 73 34 74 38
rect 78 34 79 38
rect 87 37 89 42
rect 97 39 99 42
rect 94 37 99 39
rect 22 26 24 31
rect 28 29 34 31
rect 32 26 34 29
rect 12 11 14 16
rect 22 8 24 16
rect 32 12 34 16
rect 43 8 45 32
rect 59 30 61 34
rect 73 33 79 34
rect 94 33 96 37
rect 108 33 110 72
rect 73 31 83 33
rect 81 28 83 31
rect 91 31 96 33
rect 101 31 110 33
rect 91 28 93 31
rect 101 28 103 31
rect 59 15 61 20
rect 81 13 83 18
rect 91 8 93 18
rect 101 13 103 18
rect 22 6 93 8
<< ndiffusion >>
rect 3 21 12 26
rect 3 17 5 21
rect 9 17 12 21
rect 3 16 12 17
rect 14 25 22 26
rect 14 21 16 25
rect 20 21 22 25
rect 14 16 22 21
rect 24 25 32 26
rect 24 21 26 25
rect 30 21 32 25
rect 24 16 32 21
rect 34 23 39 26
rect 34 22 41 23
rect 34 18 36 22
rect 40 18 41 22
rect 34 16 41 18
rect 52 29 59 30
rect 52 25 53 29
rect 57 25 59 29
rect 52 24 59 25
rect 54 20 59 24
rect 61 28 66 30
rect 61 23 81 28
rect 61 20 71 23
rect 63 19 71 20
rect 75 19 81 23
rect 63 18 81 19
rect 83 27 91 28
rect 83 23 85 27
rect 89 23 91 27
rect 83 18 91 23
rect 93 23 101 28
rect 93 19 95 23
rect 99 19 101 23
rect 93 18 101 19
rect 103 27 110 28
rect 103 23 105 27
rect 109 23 110 27
rect 103 22 110 23
rect 103 18 108 22
<< pdiffusion >>
rect 20 63 25 64
rect 7 62 15 63
rect 7 58 9 62
rect 13 58 15 62
rect 7 55 15 58
rect 7 51 9 55
rect 13 51 15 55
rect 7 42 15 51
rect 17 54 25 63
rect 17 50 19 54
rect 23 50 25 54
rect 17 47 25 50
rect 17 43 19 47
rect 23 43 25 47
rect 17 42 25 43
rect 27 54 35 64
rect 27 50 29 54
rect 33 50 35 54
rect 27 47 35 50
rect 27 43 29 47
rect 33 43 35 47
rect 27 42 35 43
rect 37 55 42 64
rect 37 54 44 55
rect 37 50 39 54
rect 43 50 44 54
rect 51 53 56 69
rect 37 47 44 50
rect 49 52 56 53
rect 49 48 50 52
rect 54 48 56 52
rect 49 47 56 48
rect 58 68 75 69
rect 58 64 63 68
rect 67 64 75 68
rect 58 47 77 64
rect 37 43 39 47
rect 43 43 44 47
rect 37 42 44 43
rect 67 42 77 47
rect 79 54 87 64
rect 79 50 81 54
rect 85 50 87 54
rect 79 47 87 50
rect 79 43 81 47
rect 85 43 87 47
rect 79 42 87 43
rect 89 54 97 64
rect 89 50 91 54
rect 95 50 97 54
rect 89 47 97 50
rect 89 43 91 47
rect 95 43 97 47
rect 89 42 97 43
rect 99 63 106 64
rect 99 59 101 63
rect 105 59 106 63
rect 99 56 106 59
rect 99 52 101 56
rect 105 52 106 56
rect 99 51 106 52
rect 99 42 104 51
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect -2 68 114 78
rect 9 62 13 68
rect 62 64 63 68
rect 67 64 68 68
rect 9 55 13 58
rect 9 50 13 51
rect 19 61 52 63
rect 72 61 101 63
rect 19 59 101 61
rect 105 59 106 63
rect 19 54 23 59
rect 48 57 76 59
rect 100 56 106 59
rect 19 47 23 50
rect 2 41 14 47
rect 2 38 7 41
rect 19 38 23 43
rect 2 34 3 38
rect 2 25 7 34
rect 16 34 23 38
rect 26 54 33 55
rect 26 50 29 54
rect 26 47 33 50
rect 26 43 29 47
rect 26 42 33 43
rect 39 54 43 55
rect 81 54 85 55
rect 39 47 43 50
rect 16 25 20 34
rect 4 17 5 21
rect 9 17 10 21
rect 16 20 20 21
rect 26 31 30 42
rect 39 39 43 43
rect 50 52 54 53
rect 65 50 78 54
rect 39 35 46 39
rect 26 25 38 31
rect 42 22 46 35
rect 50 37 54 48
rect 57 39 63 46
rect 57 35 60 39
rect 64 35 70 39
rect 57 33 70 35
rect 74 38 78 50
rect 74 33 78 34
rect 81 47 85 50
rect 50 29 54 33
rect 81 30 85 43
rect 90 54 95 55
rect 90 50 91 54
rect 100 52 101 56
rect 90 47 95 50
rect 90 43 91 47
rect 90 39 95 43
rect 90 33 102 39
rect 50 25 53 29
rect 57 25 58 29
rect 62 27 89 30
rect 62 26 85 27
rect 62 22 66 26
rect 98 23 102 33
rect 26 17 30 21
rect 35 18 36 22
rect 40 18 66 22
rect 70 19 71 23
rect 75 19 76 23
rect 85 22 89 23
rect 4 12 10 17
rect 47 12 53 15
rect 70 12 76 19
rect 94 19 95 23
rect 99 19 102 23
rect 105 27 109 56
rect 105 22 109 23
rect 94 17 102 19
rect -2 2 114 12
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
<< ntransistor >>
rect 12 16 14 26
rect 22 16 24 26
rect 32 16 34 26
rect 59 20 61 30
rect 81 18 83 28
rect 91 18 93 28
rect 101 18 103 28
<< ptransistor >>
rect 15 42 17 63
rect 25 42 27 64
rect 35 42 37 64
rect 56 47 58 69
rect 77 42 79 64
rect 87 42 89 64
rect 97 42 99 64
<< polycontact >>
rect 3 34 7 38
rect 50 33 54 37
rect 60 35 64 39
rect 74 34 78 38
<< ndcontact >>
rect 5 17 9 21
rect 16 21 20 25
rect 26 21 30 25
rect 36 18 40 22
rect 53 25 57 29
rect 71 19 75 23
rect 85 23 89 27
rect 95 19 99 23
rect 105 23 109 27
<< pdcontact >>
rect 9 58 13 62
rect 9 51 13 55
rect 19 50 23 54
rect 19 43 23 47
rect 29 50 33 54
rect 29 43 33 47
rect 39 50 43 54
rect 50 48 54 52
rect 63 64 67 68
rect 39 43 43 47
rect 81 50 85 54
rect 81 43 85 47
rect 91 50 95 54
rect 91 43 95 47
rect 101 59 105 63
rect 101 52 105 56
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
rect 90 -2 94 2
rect 98 -2 102 2
rect 106 -2 110 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
rect 90 78 94 82
rect 98 78 102 82
rect 106 78 110 82
<< psubstratepdiff >>
rect 0 2 112 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 112 2
rect 0 -3 112 -2
<< nsubstratendiff >>
rect 0 82 112 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 112 82
rect 0 77 112 78
<< labels >>
rlabel polysilicon 49 35 49 35 6 sn
rlabel metal1 18 29 18 29 6 a0n
rlabel polycontact 4 36 4 36 6 a0
rlabel metal1 12 44 12 44 6 a0
rlabel metal1 36 28 36 28 6 z0
rlabel metal1 28 36 28 36 6 z0
rlabel pdcontact 41 45 41 45 6 a1n
rlabel metal1 21 48 21 48 6 a0n
rlabel metal1 56 6 56 6 6 vss
rlabel metal1 50 20 50 20 6 a1n
rlabel metal1 60 40 60 40 6 s
rlabel metal1 52 39 52 39 6 sn
rlabel metal1 56 74 56 74 6 vdd
rlabel metal1 75 28 75 28 6 a1n
rlabel metal1 68 36 68 36 6 s
rlabel metal1 76 40 76 40 6 a1
rlabel metal1 68 52 68 52 6 a1
rlabel metal1 83 40 83 40 6 a1n
rlabel metal1 100 28 100 28 6 z1
rlabel pdcontact 92 44 92 44 6 z1
rlabel metal1 107 39 107 39 6 a0n
rlabel metal1 89 61 89 61 6 a0n
<< end >>
