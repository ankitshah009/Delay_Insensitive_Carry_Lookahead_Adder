magic
tech scmos
timestamp 1170759807
<< checkpaint >>
rect -22 -26 86 114
<< pwell >>
rect -4 -8 68 40
<< nwell >>
rect -4 40 68 96
<< polysilicon >>
rect 2 77 11 83
rect 9 74 11 77
rect 21 82 30 83
rect 21 78 25 82
rect 29 78 30 82
rect 21 77 30 78
rect 34 77 43 83
rect 21 74 23 77
rect 41 74 43 77
rect 53 82 62 83
rect 53 78 54 82
rect 58 78 62 82
rect 53 77 62 78
rect 53 74 55 77
rect 9 43 11 46
rect 21 43 23 46
rect 41 43 43 46
rect 53 43 55 46
rect 2 42 14 43
rect 2 38 6 42
rect 10 38 14 42
rect 2 37 14 38
rect 18 37 30 43
rect 34 42 46 43
rect 34 38 38 42
rect 42 38 46 42
rect 34 37 46 38
rect 50 42 62 43
rect 50 38 54 42
rect 58 38 62 42
rect 50 37 62 38
rect 9 34 11 37
rect 21 34 23 37
rect 41 34 43 37
rect 53 34 55 37
rect 9 11 11 14
rect 2 5 11 11
rect 21 11 23 14
rect 41 11 43 14
rect 21 5 30 11
rect 34 5 43 11
rect 53 11 55 14
rect 53 5 62 11
<< ndiffusion >>
rect 2 30 9 34
rect 2 26 3 30
rect 7 26 9 30
rect 2 22 9 26
rect 2 18 3 22
rect 7 18 9 22
rect 2 14 9 18
rect 11 14 21 34
rect 23 19 30 34
rect 23 15 25 19
rect 29 15 30 19
rect 23 14 30 15
rect 34 30 41 34
rect 34 26 35 30
rect 39 26 41 30
rect 34 22 41 26
rect 34 18 35 22
rect 39 18 41 22
rect 34 14 41 18
rect 43 14 53 34
rect 55 26 62 34
rect 55 22 57 26
rect 61 22 62 26
rect 55 19 62 22
rect 55 15 57 19
rect 61 15 62 19
rect 55 14 62 15
rect 13 2 19 14
rect 45 2 51 14
<< pdiffusion >>
rect 13 74 19 86
rect 45 74 51 86
rect 2 73 9 74
rect 2 69 3 73
rect 7 69 9 73
rect 2 66 9 69
rect 2 62 3 66
rect 7 62 9 66
rect 2 46 9 62
rect 11 62 21 74
rect 11 58 14 62
rect 18 58 21 62
rect 11 54 21 58
rect 11 50 14 54
rect 18 50 21 54
rect 11 46 21 50
rect 23 73 30 74
rect 23 69 25 73
rect 29 69 30 73
rect 23 66 30 69
rect 23 62 25 66
rect 29 62 30 66
rect 23 46 30 62
rect 34 73 41 74
rect 34 69 35 73
rect 39 69 41 73
rect 34 66 41 69
rect 34 62 35 66
rect 39 62 41 66
rect 34 46 41 62
rect 43 58 53 74
rect 43 54 46 58
rect 50 54 53 58
rect 43 51 53 54
rect 43 47 46 51
rect 50 47 53 51
rect 43 46 53 47
rect 55 73 62 74
rect 55 69 57 73
rect 61 69 62 73
rect 55 66 62 69
rect 55 62 57 66
rect 61 62 62 66
rect 55 46 62 62
<< metal1 >>
rect -2 86 2 90
rect 10 86 22 90
rect 30 86 34 90
rect 42 86 54 90
rect 62 86 66 90
rect 6 82 10 86
rect 24 78 25 82
rect 29 78 54 82
rect 58 78 59 82
rect 6 74 10 78
rect 3 73 61 74
rect 7 70 25 73
rect 3 66 7 69
rect 29 70 35 73
rect 25 66 29 69
rect 3 61 7 62
rect 14 62 18 63
rect 25 61 29 62
rect 39 70 57 73
rect 35 66 39 69
rect 57 66 61 69
rect 35 61 39 62
rect 14 56 18 58
rect 46 58 50 63
rect 57 61 61 62
rect 6 42 10 55
rect 14 54 46 56
rect 18 52 50 54
rect 14 49 18 50
rect 46 51 50 52
rect 38 42 42 47
rect 6 34 42 38
rect 46 30 50 47
rect 54 42 58 55
rect 54 33 58 38
rect 2 26 3 30
rect 7 26 35 30
rect 39 26 50 30
rect 6 22 11 26
rect 2 18 3 22
rect 7 18 11 22
rect 35 25 50 26
rect 57 26 61 27
rect 35 22 39 25
rect 25 19 29 20
rect 35 17 39 18
rect 57 19 61 22
rect 25 10 29 15
rect 25 2 29 6
rect 57 10 61 15
rect 57 2 61 6
rect -2 -2 2 2
rect 10 -2 22 2
rect 30 -2 34 2
rect 42 -2 54 2
rect 62 -2 66 2
<< metal2 >>
rect -2 86 6 90
rect 10 86 22 90
rect 26 86 38 90
rect 42 86 54 90
rect 58 86 66 90
rect -2 82 66 86
rect -2 78 6 82
rect 10 78 66 82
rect -2 76 66 78
rect -2 10 66 12
rect -2 6 25 10
rect 29 6 57 10
rect 61 6 66 10
rect -2 2 66 6
rect -2 -2 6 2
rect 10 -2 22 2
rect 26 -2 38 2
rect 42 -2 54 2
rect 58 -2 66 2
<< ntransistor >>
rect 9 14 11 34
rect 21 14 23 34
rect 41 14 43 34
rect 53 14 55 34
<< ptransistor >>
rect 9 46 11 74
rect 21 46 23 74
rect 41 46 43 74
rect 53 46 55 74
<< polycontact >>
rect 25 78 29 82
rect 54 78 58 82
rect 6 38 10 42
rect 38 38 42 42
rect 54 38 58 42
<< ndcontact >>
rect 3 26 7 30
rect 3 18 7 22
rect 25 15 29 19
rect 35 26 39 30
rect 35 18 39 22
rect 57 22 61 26
rect 57 15 61 19
<< pdcontact >>
rect 3 69 7 73
rect 3 62 7 66
rect 14 58 18 62
rect 14 50 18 54
rect 25 69 29 73
rect 25 62 29 66
rect 35 69 39 73
rect 35 62 39 66
rect 46 54 50 58
rect 46 47 50 51
rect 57 69 61 73
rect 57 62 61 66
<< m2contact >>
rect 6 86 10 90
rect 22 86 26 90
rect 38 86 42 90
rect 54 86 58 90
rect 6 78 10 82
rect 25 6 29 10
rect 57 6 61 10
rect 6 -2 10 2
rect 22 -2 26 2
rect 38 -2 42 2
rect 54 -2 58 2
<< psubstratepcontact >>
rect 2 -2 6 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 58 -2 62 2
<< nsubstratencontact >>
rect 2 86 6 90
rect 26 86 30 90
rect 34 86 38 90
rect 58 86 62 90
<< psubstratepdiff >>
rect 0 2 7 3
rect 25 2 39 3
rect 57 2 64 3
rect 0 -2 2 2
rect 6 -2 7 2
rect 0 -3 7 -2
rect 25 -2 26 2
rect 30 -2 34 2
rect 38 -2 39 2
rect 25 -3 39 -2
rect 57 -2 58 2
rect 62 -2 64 2
rect 57 -3 64 -2
<< nsubstratendiff >>
rect 0 90 7 91
rect 0 86 2 90
rect 6 86 7 90
rect 25 90 39 91
rect 25 86 26 90
rect 30 86 34 90
rect 38 86 39 90
rect 57 90 64 91
rect 57 86 58 90
rect 62 86 64 90
rect 0 85 7 86
rect 25 85 39 86
rect 57 85 64 86
<< labels >>
rlabel metal1 8 24 8 24 6 z
rlabel metal1 8 48 8 48 6 b
rlabel metal1 16 28 16 28 6 z
rlabel metal1 16 36 16 36 6 b
rlabel metal1 24 28 24 28 6 z
rlabel metal1 32 28 32 28 6 z
rlabel metal1 32 36 32 36 6 b
rlabel metal1 24 36 24 36 6 b
rlabel metal1 40 28 40 28 6 z
rlabel metal1 40 44 40 44 6 b
rlabel metal1 48 44 48 44 6 z
rlabel metal1 56 44 56 44 6 a
rlabel metal2 32 6 32 6 6 vss
rlabel metal2 32 82 32 82 6 vdd
<< end >>
