magic
tech scmos
timestamp 1179386485
<< checkpaint >>
rect -22 -25 94 105
<< ab >>
rect 0 0 72 80
<< pwell >>
rect -4 -7 76 36
<< nwell >>
rect -4 36 76 87
<< polysilicon >>
rect 9 69 11 74
rect 19 69 21 74
rect 29 69 31 74
rect 39 69 41 74
rect 49 69 51 74
rect 59 69 61 74
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 39 39 41 42
rect 49 39 51 42
rect 59 39 61 42
rect 9 38 15 39
rect 9 34 10 38
rect 14 34 15 38
rect 9 33 15 34
rect 19 38 33 39
rect 19 34 26 38
rect 30 34 33 38
rect 19 33 33 34
rect 12 30 14 33
rect 19 30 21 33
rect 31 30 33 33
rect 38 38 51 39
rect 38 34 42 38
rect 46 34 51 38
rect 38 33 51 34
rect 55 38 61 39
rect 55 34 56 38
rect 60 34 61 38
rect 55 33 61 34
rect 38 30 40 33
rect 48 30 50 33
rect 55 30 57 33
rect 12 15 14 19
rect 19 14 21 19
rect 31 6 33 10
rect 38 6 40 10
rect 48 6 50 10
rect 55 6 57 10
<< ndiffusion >>
rect 5 29 12 30
rect 5 25 6 29
rect 10 25 12 29
rect 5 24 12 25
rect 7 19 12 24
rect 14 19 19 30
rect 21 19 31 30
rect 23 15 31 19
rect 23 11 24 15
rect 28 11 31 15
rect 23 10 31 11
rect 33 10 38 30
rect 40 22 48 30
rect 40 18 42 22
rect 46 18 48 22
rect 40 10 48 18
rect 50 10 55 30
rect 57 12 66 30
rect 57 10 60 12
rect 59 8 60 10
rect 64 8 66 12
rect 59 7 66 8
<< pdiffusion >>
rect 2 68 9 69
rect 2 64 3 68
rect 7 64 9 68
rect 2 61 9 64
rect 2 57 3 61
rect 7 57 9 61
rect 2 42 9 57
rect 11 62 19 69
rect 11 58 13 62
rect 17 58 19 62
rect 11 54 19 58
rect 11 50 13 54
rect 17 50 19 54
rect 11 42 19 50
rect 21 68 29 69
rect 21 64 23 68
rect 27 64 29 68
rect 21 61 29 64
rect 21 57 23 61
rect 27 57 29 61
rect 21 42 29 57
rect 31 62 39 69
rect 31 58 33 62
rect 37 58 39 62
rect 31 54 39 58
rect 31 50 33 54
rect 37 50 39 54
rect 31 42 39 50
rect 41 68 49 69
rect 41 64 43 68
rect 47 64 49 68
rect 41 61 49 64
rect 41 57 43 61
rect 47 57 49 61
rect 41 42 49 57
rect 51 62 59 69
rect 51 58 53 62
rect 57 58 59 62
rect 51 55 59 58
rect 51 51 53 55
rect 57 51 59 55
rect 51 42 59 51
rect 61 68 68 69
rect 61 64 63 68
rect 67 64 68 68
rect 61 61 68 64
rect 61 57 63 61
rect 67 57 68 61
rect 61 42 68 57
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect -2 68 74 78
rect 2 64 3 68
rect 7 64 8 68
rect 2 61 8 64
rect 22 64 23 68
rect 27 64 28 68
rect 2 57 3 61
rect 7 57 8 61
rect 13 62 17 63
rect 13 54 17 58
rect 22 61 28 64
rect 42 64 43 68
rect 47 64 48 68
rect 22 57 23 61
rect 27 57 28 61
rect 33 62 38 63
rect 37 58 38 62
rect 33 54 38 58
rect 42 61 48 64
rect 62 64 63 68
rect 67 64 68 68
rect 42 57 43 61
rect 47 57 48 61
rect 53 62 57 63
rect 53 55 57 58
rect 62 61 68 64
rect 62 57 63 61
rect 67 57 68 61
rect 2 50 13 54
rect 17 50 33 54
rect 37 51 53 54
rect 57 51 63 54
rect 37 50 63 51
rect 2 25 6 50
rect 25 42 63 46
rect 10 38 21 39
rect 14 34 21 38
rect 25 38 31 42
rect 55 38 61 42
rect 25 34 26 38
rect 30 34 31 38
rect 41 34 42 38
rect 46 34 47 38
rect 55 34 56 38
rect 60 34 61 38
rect 10 33 21 34
rect 17 30 21 33
rect 41 30 47 34
rect 10 25 11 29
rect 17 26 55 30
rect 7 22 11 25
rect 7 18 42 22
rect 46 18 47 22
rect 23 12 24 15
rect -2 11 24 12
rect 28 12 29 15
rect 28 11 60 12
rect -2 8 60 11
rect 64 8 74 12
rect -2 2 74 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
<< ntransistor >>
rect 12 19 14 30
rect 19 19 21 30
rect 31 10 33 30
rect 38 10 40 30
rect 48 10 50 30
rect 55 10 57 30
<< ptransistor >>
rect 9 42 11 69
rect 19 42 21 69
rect 29 42 31 69
rect 39 42 41 69
rect 49 42 51 69
rect 59 42 61 69
<< polycontact >>
rect 10 34 14 38
rect 26 34 30 38
rect 42 34 46 38
rect 56 34 60 38
<< ndcontact >>
rect 6 25 10 29
rect 24 11 28 15
rect 42 18 46 22
rect 60 8 64 12
<< pdcontact >>
rect 3 64 7 68
rect 3 57 7 61
rect 13 58 17 62
rect 13 50 17 54
rect 23 64 27 68
rect 23 57 27 61
rect 33 58 37 62
rect 33 50 37 54
rect 43 64 47 68
rect 43 57 47 61
rect 53 58 57 62
rect 53 51 57 55
rect 63 64 67 68
rect 63 57 67 61
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
<< psubstratepdiff >>
rect 0 2 72 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 72 2
rect 0 -3 72 -2
<< nsubstratendiff >>
rect 0 82 72 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 72 82
rect 0 77 72 78
<< labels >>
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 20 12 20 6 z
rlabel metal1 20 20 20 20 6 z
rlabel metal1 20 28 20 28 6 b
rlabel polycontact 12 36 12 36 6 b
rlabel metal1 20 52 20 52 6 z
rlabel metal1 12 52 12 52 6 z
rlabel metal1 36 6 36 6 6 vss
rlabel metal1 28 20 28 20 6 z
rlabel metal1 28 28 28 28 6 b
rlabel metal1 36 20 36 20 6 z
rlabel metal1 36 28 36 28 6 b
rlabel metal1 28 40 28 40 6 a
rlabel metal1 36 44 36 44 6 a
rlabel metal1 28 52 28 52 6 z
rlabel metal1 36 56 36 56 6 z
rlabel metal1 36 74 36 74 6 vdd
rlabel ndcontact 44 20 44 20 6 z
rlabel metal1 52 28 52 28 6 b
rlabel metal1 44 32 44 32 6 b
rlabel metal1 44 44 44 44 6 a
rlabel metal1 52 44 52 44 6 a
rlabel metal1 52 52 52 52 6 z
rlabel metal1 44 52 44 52 6 z
rlabel metal1 60 44 60 44 6 a
rlabel metal1 60 52 60 52 6 z
<< end >>
