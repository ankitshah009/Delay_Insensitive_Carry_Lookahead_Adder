magic
tech scmos
timestamp 1179386940
<< checkpaint >>
rect -22 -22 134 94
<< ab >>
rect 0 0 112 72
<< pwell >>
rect -4 -4 116 32
<< nwell >>
rect -4 32 116 76
<< polysilicon >>
rect 14 65 16 70
rect 21 65 23 70
rect 28 65 30 70
rect 35 65 37 70
rect 47 65 49 70
rect 54 65 56 70
rect 61 65 63 70
rect 68 65 70 70
rect 78 65 80 70
rect 85 65 87 70
rect 92 65 94 70
rect 99 65 101 70
rect 14 37 16 40
rect 9 36 16 37
rect 9 32 10 36
rect 14 32 16 36
rect 9 31 16 32
rect 10 18 12 31
rect 21 27 23 40
rect 17 26 23 27
rect 17 22 18 26
rect 22 22 23 26
rect 17 21 23 22
rect 28 27 30 40
rect 35 35 37 40
rect 47 35 49 38
rect 35 34 49 35
rect 35 33 39 34
rect 38 30 39 33
rect 43 33 49 34
rect 43 30 44 33
rect 38 29 44 30
rect 28 26 34 27
rect 28 22 29 26
rect 33 22 34 26
rect 28 21 34 22
rect 20 18 22 21
rect 32 18 34 21
rect 42 18 44 29
rect 54 27 56 38
rect 61 29 63 38
rect 68 35 70 38
rect 78 35 80 38
rect 68 34 81 35
rect 68 33 76 34
rect 75 30 76 33
rect 80 30 81 34
rect 75 29 81 30
rect 61 28 71 29
rect 61 27 66 28
rect 48 26 56 27
rect 48 22 49 26
rect 53 22 56 26
rect 65 24 66 27
rect 70 25 71 28
rect 85 25 87 38
rect 70 24 87 25
rect 65 23 87 24
rect 48 21 56 22
rect 54 19 56 21
rect 92 19 94 38
rect 10 2 12 7
rect 20 2 22 7
rect 54 17 94 19
rect 99 19 101 38
rect 99 18 105 19
rect 99 14 100 18
rect 104 14 105 18
rect 99 13 105 14
rect 32 2 34 7
rect 42 2 44 7
<< ndiffusion >>
rect 2 8 10 18
rect 2 4 3 8
rect 7 7 10 8
rect 12 17 20 18
rect 12 13 14 17
rect 18 13 20 17
rect 12 7 20 13
rect 22 8 32 18
rect 22 7 25 8
rect 7 4 8 7
rect 2 3 8 4
rect 24 4 25 7
rect 29 7 32 8
rect 34 17 42 18
rect 34 13 36 17
rect 40 13 42 17
rect 34 7 42 13
rect 44 8 52 18
rect 44 7 47 8
rect 29 4 30 7
rect 24 3 30 4
rect 46 4 47 7
rect 51 4 52 8
rect 46 3 52 4
<< pdiffusion >>
rect 39 68 45 69
rect 39 65 40 68
rect 9 59 14 65
rect 7 58 14 59
rect 7 54 8 58
rect 12 54 14 58
rect 7 53 14 54
rect 9 40 14 53
rect 16 40 21 65
rect 23 40 28 65
rect 30 40 35 65
rect 37 64 40 65
rect 44 65 45 68
rect 44 64 47 65
rect 37 40 47 64
rect 39 38 47 40
rect 49 38 54 65
rect 56 38 61 65
rect 63 38 68 65
rect 70 58 78 65
rect 70 54 72 58
rect 76 54 78 58
rect 70 38 78 54
rect 80 38 85 65
rect 87 38 92 65
rect 94 38 99 65
rect 101 64 108 65
rect 101 60 103 64
rect 107 60 108 64
rect 101 57 108 60
rect 101 53 103 57
rect 107 53 108 57
rect 101 38 108 53
<< metal1 >>
rect -2 68 114 72
rect -2 64 40 68
rect 44 64 114 68
rect 102 60 103 64
rect 107 60 108 64
rect 2 54 8 58
rect 12 54 72 58
rect 76 54 79 58
rect 102 57 108 60
rect 2 19 6 54
rect 102 53 103 57
rect 107 53 108 57
rect 10 46 80 50
rect 10 36 14 46
rect 10 29 14 32
rect 18 38 70 42
rect 18 26 22 38
rect 38 30 39 34
rect 43 30 62 34
rect 28 22 29 26
rect 33 22 49 26
rect 53 22 54 26
rect 18 21 22 22
rect 2 13 14 19
rect 33 17 41 18
rect 18 13 36 17
rect 40 13 41 17
rect 50 13 54 22
rect 58 18 62 30
rect 66 28 70 38
rect 74 34 80 46
rect 74 30 76 34
rect 74 29 80 30
rect 66 23 70 24
rect 58 14 100 18
rect 104 14 105 18
rect -2 4 3 8
rect 7 4 25 8
rect 29 4 47 8
rect 51 4 64 8
rect 68 4 72 8
rect 76 4 80 8
rect 84 4 88 8
rect 92 4 96 8
rect 100 4 104 8
rect 108 4 114 8
rect -2 0 114 4
<< ntransistor >>
rect 10 7 12 18
rect 20 7 22 18
rect 32 7 34 18
rect 42 7 44 18
<< ptransistor >>
rect 14 40 16 65
rect 21 40 23 65
rect 28 40 30 65
rect 35 40 37 65
rect 47 38 49 65
rect 54 38 56 65
rect 61 38 63 65
rect 68 38 70 65
rect 78 38 80 65
rect 85 38 87 65
rect 92 38 94 65
rect 99 38 101 65
<< polycontact >>
rect 10 32 14 36
rect 18 22 22 26
rect 39 30 43 34
rect 29 22 33 26
rect 76 30 80 34
rect 49 22 53 26
rect 66 24 70 28
rect 100 14 104 18
<< ndcontact >>
rect 3 4 7 8
rect 14 13 18 17
rect 25 4 29 8
rect 36 13 40 17
rect 47 4 51 8
<< pdcontact >>
rect 8 54 12 58
rect 40 64 44 68
rect 72 54 76 58
rect 103 60 107 64
rect 103 53 107 57
<< psubstratepcontact >>
rect 64 4 68 8
rect 72 4 76 8
rect 80 4 84 8
rect 88 4 92 8
rect 96 4 100 8
rect 104 4 108 8
<< psubstratepdiff >>
rect 63 8 109 9
rect 63 4 64 8
rect 68 4 72 8
rect 76 4 80 8
rect 84 4 88 8
rect 92 4 96 8
rect 100 4 104 8
rect 108 4 109 8
rect 63 3 109 4
<< labels >>
rlabel metal1 12 16 12 16 6 z
rlabel metal1 4 32 4 32 6 z
rlabel metal1 12 36 12 36 6 d
rlabel metal1 12 56 12 56 6 z
rlabel metal1 36 16 36 16 6 z
rlabel metal1 36 24 36 24 6 b
rlabel metal1 20 28 20 28 6 c
rlabel metal1 28 40 28 40 6 c
rlabel metal1 36 40 36 40 6 c
rlabel metal1 20 48 20 48 6 d
rlabel metal1 28 48 28 48 6 d
rlabel metal1 36 48 36 48 6 d
rlabel metal1 28 56 28 56 6 z
rlabel metal1 36 56 36 56 6 z
rlabel metal1 20 56 20 56 6 z
rlabel metal1 56 4 56 4 6 vss
rlabel metal1 52 16 52 16 6 b
rlabel metal1 44 24 44 24 6 b
rlabel metal1 60 24 60 24 6 a
rlabel metal1 52 32 52 32 6 a
rlabel metal1 44 32 44 32 6 a
rlabel metal1 44 40 44 40 6 c
rlabel metal1 52 40 52 40 6 c
rlabel metal1 60 40 60 40 6 c
rlabel metal1 44 48 44 48 6 d
rlabel metal1 52 48 52 48 6 d
rlabel metal1 60 48 60 48 6 d
rlabel metal1 52 56 52 56 6 z
rlabel metal1 60 56 60 56 6 z
rlabel metal1 44 56 44 56 6 z
rlabel metal1 56 68 56 68 6 vdd
rlabel metal1 76 16 76 16 6 a
rlabel metal1 84 16 84 16 6 a
rlabel metal1 68 16 68 16 6 a
rlabel metal1 68 32 68 32 6 c
rlabel metal1 76 40 76 40 6 d
rlabel metal1 68 48 68 48 6 d
rlabel metal1 76 56 76 56 6 z
rlabel metal1 68 56 68 56 6 z
rlabel metal1 100 16 100 16 6 a
rlabel metal1 92 16 92 16 6 a
<< end >>
