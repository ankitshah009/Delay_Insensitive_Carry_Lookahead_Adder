magic
tech scmos
timestamp 1179387612
<< checkpaint >>
rect -22 -25 158 105
<< ab >>
rect 0 0 136 80
<< pwell >>
rect -4 -7 140 36
<< nwell >>
rect -4 36 140 87
<< polysilicon >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 39 70 41 74
rect 49 70 51 74
rect 59 70 61 74
rect 66 70 68 74
rect 78 72 104 74
rect 78 63 80 72
rect 85 66 97 68
rect 85 63 87 66
rect 95 63 97 66
rect 102 63 104 72
rect 115 70 117 74
rect 125 61 127 65
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 39 39 41 42
rect 49 39 51 42
rect 59 39 61 42
rect 9 37 21 39
rect 25 38 51 39
rect 9 36 15 37
rect 9 32 10 36
rect 14 32 15 36
rect 25 34 26 38
rect 30 37 51 38
rect 55 38 61 39
rect 30 34 31 37
rect 25 33 31 34
rect 55 34 56 38
rect 60 34 61 38
rect 66 39 68 42
rect 78 39 80 42
rect 66 37 80 39
rect 85 39 87 42
rect 85 38 91 39
rect 95 38 97 42
rect 102 39 104 42
rect 115 39 117 42
rect 125 39 127 42
rect 101 38 107 39
rect 55 33 61 34
rect 85 34 86 38
rect 90 34 91 38
rect 101 34 102 38
rect 106 34 107 38
rect 85 33 91 34
rect 9 31 15 32
rect 19 31 31 33
rect 12 28 14 31
rect 19 28 21 31
rect 29 28 31 31
rect 36 28 38 33
rect 55 30 57 33
rect 12 8 14 16
rect 19 12 21 16
rect 29 12 31 16
rect 36 8 38 16
rect 12 6 38 8
rect 75 29 77 33
rect 85 29 87 33
rect 95 32 107 34
rect 95 29 97 32
rect 105 29 107 32
rect 115 38 127 39
rect 115 34 122 38
rect 126 34 127 38
rect 115 33 127 34
rect 115 30 117 33
rect 125 30 127 33
rect 55 10 57 15
rect 125 16 127 20
rect 85 12 87 16
rect 95 12 97 16
rect 105 12 107 16
rect 75 8 77 11
rect 115 8 117 16
rect 75 6 117 8
<< ndiffusion >>
rect 40 28 55 30
rect 3 16 12 28
rect 14 16 19 28
rect 21 22 29 28
rect 21 18 23 22
rect 27 18 29 22
rect 21 16 29 18
rect 31 16 36 28
rect 38 16 55 28
rect 3 12 10 16
rect 3 8 5 12
rect 9 8 10 12
rect 3 7 10 8
rect 40 15 55 16
rect 57 29 64 30
rect 109 29 115 30
rect 57 25 59 29
rect 63 25 64 29
rect 57 24 64 25
rect 57 15 62 24
rect 70 23 75 29
rect 68 22 75 23
rect 68 18 69 22
rect 73 18 75 22
rect 68 17 75 18
rect 40 12 53 15
rect 40 8 41 12
rect 45 8 48 12
rect 52 8 53 12
rect 70 11 75 17
rect 77 28 85 29
rect 77 24 79 28
rect 83 24 85 28
rect 77 21 85 24
rect 77 17 79 21
rect 83 17 85 21
rect 77 16 85 17
rect 87 21 95 29
rect 87 17 89 21
rect 93 17 95 21
rect 87 16 95 17
rect 97 28 105 29
rect 97 24 99 28
rect 103 24 105 28
rect 97 21 105 24
rect 97 17 99 21
rect 103 17 105 21
rect 97 16 105 17
rect 107 21 115 29
rect 107 17 109 21
rect 113 17 115 21
rect 107 16 115 17
rect 117 29 125 30
rect 117 25 119 29
rect 123 25 125 29
rect 117 20 125 25
rect 127 25 134 30
rect 127 21 129 25
rect 133 21 134 25
rect 127 20 134 21
rect 117 16 122 20
rect 77 11 82 16
rect 40 7 53 8
<< pdiffusion >>
rect 70 72 76 73
rect 70 70 71 72
rect 4 63 9 70
rect 2 62 9 63
rect 2 58 3 62
rect 7 58 9 62
rect 2 55 9 58
rect 2 51 3 55
rect 7 51 9 55
rect 2 50 9 51
rect 4 42 9 50
rect 11 55 19 70
rect 11 51 13 55
rect 17 51 19 55
rect 11 47 19 51
rect 11 43 13 47
rect 17 43 19 47
rect 11 42 19 43
rect 21 62 29 70
rect 21 58 23 62
rect 27 58 29 62
rect 21 42 29 58
rect 31 47 39 70
rect 31 43 33 47
rect 37 43 39 47
rect 31 42 39 43
rect 41 62 49 70
rect 41 58 43 62
rect 47 58 49 62
rect 41 42 49 58
rect 51 47 59 70
rect 51 43 53 47
rect 57 43 59 47
rect 51 42 59 43
rect 61 42 66 70
rect 68 68 71 70
rect 75 68 76 72
rect 68 63 76 68
rect 106 72 113 73
rect 106 68 108 72
rect 112 70 113 72
rect 112 68 115 70
rect 106 63 115 68
rect 68 42 78 63
rect 80 42 85 63
rect 87 54 95 63
rect 87 50 89 54
rect 93 50 95 54
rect 87 47 95 50
rect 87 43 89 47
rect 93 43 95 47
rect 87 42 95 43
rect 97 42 102 63
rect 104 42 115 63
rect 117 61 122 70
rect 117 55 125 61
rect 117 51 119 55
rect 123 51 125 55
rect 117 48 125 51
rect 117 44 119 48
rect 123 44 125 48
rect 117 42 125 44
rect 127 60 134 61
rect 127 56 129 60
rect 133 56 134 60
rect 127 42 134 56
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect 118 78 122 82
rect 126 78 130 82
rect 134 78 138 82
rect -2 72 138 78
rect -2 68 71 72
rect 75 68 108 72
rect 112 68 138 72
rect 2 58 3 62
rect 7 58 23 62
rect 27 58 43 62
rect 47 58 48 62
rect 54 59 123 63
rect 2 55 7 58
rect 54 55 58 59
rect 119 55 123 59
rect 129 60 133 68
rect 129 55 133 56
rect 2 51 3 55
rect 12 51 13 55
rect 17 51 58 55
rect 64 54 93 55
rect 64 51 89 54
rect 2 50 7 51
rect 2 22 6 50
rect 24 47 28 51
rect 64 47 68 51
rect 89 47 93 50
rect 119 48 123 51
rect 12 43 13 47
rect 17 43 28 47
rect 32 43 33 47
rect 37 43 53 47
rect 57 43 68 47
rect 24 38 28 43
rect 10 36 14 37
rect 24 34 26 38
rect 30 34 31 38
rect 10 30 14 32
rect 34 30 38 43
rect 74 38 78 47
rect 89 42 93 43
rect 106 39 110 47
rect 98 38 110 39
rect 49 34 56 38
rect 60 34 86 38
rect 90 34 91 38
rect 98 34 102 38
rect 106 34 110 38
rect 98 33 110 34
rect 10 29 103 30
rect 10 26 59 29
rect 58 25 59 26
rect 63 28 103 29
rect 63 26 79 28
rect 63 25 64 26
rect 83 26 99 28
rect 2 18 23 22
rect 27 18 69 22
rect 73 18 74 22
rect 79 21 83 24
rect 106 25 110 33
rect 114 44 119 47
rect 114 43 123 44
rect 114 29 118 43
rect 130 39 134 47
rect 122 38 134 39
rect 126 34 134 38
rect 122 33 134 34
rect 114 25 119 29
rect 123 25 124 29
rect 129 25 133 26
rect 99 21 103 24
rect 79 16 83 17
rect 88 17 89 21
rect 93 17 94 21
rect 88 12 94 17
rect 99 16 103 17
rect 108 17 109 21
rect 113 17 114 21
rect 108 12 114 17
rect 129 12 133 21
rect -2 8 5 12
rect 9 8 41 12
rect 45 8 48 12
rect 52 8 138 12
rect -2 2 138 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 122 2
rect 126 -2 130 2
rect 134 -2 138 2
<< ntransistor >>
rect 12 16 14 28
rect 19 16 21 28
rect 29 16 31 28
rect 36 16 38 28
rect 55 15 57 30
rect 75 11 77 29
rect 85 16 87 29
rect 95 16 97 29
rect 105 16 107 29
rect 115 16 117 30
rect 125 20 127 30
<< ptransistor >>
rect 9 42 11 70
rect 19 42 21 70
rect 29 42 31 70
rect 39 42 41 70
rect 49 42 51 70
rect 59 42 61 70
rect 66 42 68 70
rect 78 42 80 63
rect 85 42 87 63
rect 95 42 97 63
rect 102 42 104 63
rect 115 42 117 70
rect 125 42 127 61
<< polycontact >>
rect 10 32 14 36
rect 26 34 30 38
rect 56 34 60 38
rect 86 34 90 38
rect 102 34 106 38
rect 122 34 126 38
<< ndcontact >>
rect 23 18 27 22
rect 5 8 9 12
rect 59 25 63 29
rect 69 18 73 22
rect 41 8 45 12
rect 48 8 52 12
rect 79 24 83 28
rect 79 17 83 21
rect 89 17 93 21
rect 99 24 103 28
rect 99 17 103 21
rect 109 17 113 21
rect 119 25 123 29
rect 129 21 133 25
<< pdcontact >>
rect 3 58 7 62
rect 3 51 7 55
rect 13 51 17 55
rect 13 43 17 47
rect 23 58 27 62
rect 33 43 37 47
rect 43 58 47 62
rect 53 43 57 47
rect 71 68 75 72
rect 108 68 112 72
rect 89 50 93 54
rect 89 43 93 47
rect 119 51 123 55
rect 119 44 123 48
rect 129 56 133 60
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
rect 90 -2 94 2
rect 98 -2 102 2
rect 106 -2 110 2
rect 114 -2 118 2
rect 122 -2 126 2
rect 130 -2 134 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
rect 90 78 94 82
rect 98 78 102 82
rect 106 78 110 82
rect 114 78 118 82
rect 122 78 126 82
rect 130 78 134 82
<< psubstratepdiff >>
rect 0 2 136 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 122 2
rect 126 -2 130 2
rect 134 -2 136 2
rect 0 -3 136 -2
<< nsubstratendiff >>
rect 0 82 136 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect 118 78 122 82
rect 126 78 130 82
rect 134 78 136 82
rect 0 77 136 78
<< labels >>
rlabel ntransistor 13 22 13 22 6 an
rlabel polycontact 28 35 28 35 6 bn
rlabel metal1 12 20 12 20 6 z
rlabel metal1 20 20 20 20 6 z
rlabel metal1 12 31 12 31 6 an
rlabel metal1 4 40 4 40 6 z
rlabel metal1 12 60 12 60 6 z
rlabel metal1 20 60 20 60 6 z
rlabel metal1 28 20 28 20 6 z
rlabel metal1 36 20 36 20 6 z
rlabel metal1 44 20 44 20 6 z
rlabel metal1 20 45 20 45 6 bn
rlabel metal1 26 44 26 44 6 bn
rlabel metal1 28 60 28 60 6 z
rlabel metal1 36 60 36 60 6 z
rlabel pdcontact 44 60 44 60 6 z
rlabel metal1 68 6 68 6 6 vss
rlabel metal1 52 20 52 20 6 z
rlabel metal1 60 20 60 20 6 z
rlabel metal1 68 20 68 20 6 z
rlabel metal1 52 36 52 36 6 a2
rlabel metal1 50 45 50 45 6 an
rlabel metal1 60 36 60 36 6 a2
rlabel metal1 68 36 68 36 6 a2
rlabel metal1 76 40 76 40 6 a2
rlabel metal1 35 53 35 53 6 bn
rlabel metal1 68 74 68 74 6 vdd
rlabel metal1 101 23 101 23 6 an
rlabel metal1 81 23 81 23 6 an
rlabel metal1 56 28 56 28 6 an
rlabel metal1 84 36 84 36 6 a2
rlabel metal1 100 36 100 36 6 a1
rlabel metal1 108 36 108 36 6 a1
rlabel metal1 91 48 91 48 6 an
rlabel metal1 119 27 119 27 6 bn
rlabel polycontact 124 36 124 36 6 b
rlabel metal1 132 40 132 40 6 b
rlabel pdcontact 121 53 121 53 6 bn
<< end >>
