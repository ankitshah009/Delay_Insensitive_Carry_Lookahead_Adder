magic
tech scmos
timestamp 1179385780
<< checkpaint >>
rect -22 -22 86 94
<< ab >>
rect 0 0 64 72
<< pwell >>
rect -4 -4 68 32
<< nwell >>
rect -4 32 68 76
<< polysilicon >>
rect 9 64 11 70
rect 20 68 26 69
rect 20 64 21 68
rect 25 64 26 68
rect 20 63 26 64
rect 9 43 11 46
rect 9 42 18 43
rect 9 41 13 42
rect 12 38 13 41
rect 17 38 18 42
rect 12 26 18 38
rect 22 36 26 63
rect 36 57 38 62
rect 43 57 45 62
rect 36 46 38 49
rect 43 46 45 49
rect 32 45 38 46
rect 32 41 33 45
rect 37 41 38 45
rect 32 40 38 41
rect 42 45 48 46
rect 42 41 43 45
rect 47 41 48 45
rect 42 40 48 41
rect 22 34 37 36
rect 9 24 18 26
rect 23 29 29 30
rect 23 25 24 29
rect 28 25 29 29
rect 23 24 29 25
rect 33 28 37 34
rect 33 24 49 28
rect 9 21 11 24
rect 16 21 18 24
rect 26 21 28 24
rect 33 21 35 24
rect 40 21 42 24
rect 47 21 49 24
rect 26 10 28 15
rect 33 10 35 15
rect 40 10 42 15
rect 47 11 49 15
rect 9 2 11 6
rect 16 2 18 6
<< ndiffusion >>
rect 2 20 9 21
rect 2 16 3 20
rect 7 16 9 20
rect 2 6 9 16
rect 11 6 16 21
rect 18 20 26 21
rect 18 16 20 20
rect 24 16 26 20
rect 18 15 26 16
rect 28 15 33 21
rect 35 15 40 21
rect 42 15 47 21
rect 49 20 56 21
rect 49 16 51 20
rect 55 16 56 20
rect 49 15 56 16
rect 18 6 24 15
<< pdiffusion >>
rect 2 59 9 64
rect 2 55 3 59
rect 7 55 9 59
rect 2 51 9 55
rect 2 47 3 51
rect 7 47 9 51
rect 2 46 9 47
rect 11 63 18 64
rect 11 59 13 63
rect 17 59 18 63
rect 11 46 18 59
rect 28 68 34 69
rect 28 64 29 68
rect 33 64 34 68
rect 28 57 34 64
rect 28 49 36 57
rect 38 49 43 57
rect 45 54 56 57
rect 45 50 51 54
rect 55 50 56 54
rect 45 49 56 50
<< metal1 >>
rect -2 68 66 72
rect -2 64 21 68
rect 25 64 29 68
rect 33 64 52 68
rect 56 64 66 68
rect 12 63 18 64
rect 12 59 13 63
rect 17 59 18 63
rect 2 55 3 59
rect 7 55 8 59
rect 12 56 18 59
rect 2 52 8 55
rect 22 54 56 59
rect 22 53 51 54
rect 2 51 18 52
rect 2 47 3 51
rect 7 47 18 51
rect 2 46 18 47
rect 2 34 8 46
rect 22 42 28 53
rect 50 50 51 53
rect 55 50 56 54
rect 12 38 13 42
rect 17 38 28 42
rect 33 45 39 46
rect 37 41 39 45
rect 33 34 39 41
rect 2 28 19 34
rect 23 30 39 34
rect 43 45 47 49
rect 23 29 29 30
rect 2 20 8 28
rect 23 25 24 29
rect 28 25 29 29
rect 23 24 29 25
rect 2 16 3 20
rect 7 16 8 20
rect 2 13 8 16
rect 19 16 20 20
rect 24 16 25 20
rect 19 8 25 16
rect 43 8 47 41
rect 50 20 56 50
rect 50 16 51 20
rect 55 16 56 20
rect 50 13 56 16
rect -2 4 52 8
rect 56 4 66 8
rect -2 0 66 4
<< ntransistor >>
rect 9 6 11 21
rect 16 6 18 21
rect 26 15 28 21
rect 33 15 35 21
rect 40 15 42 21
rect 47 15 49 21
<< ptransistor >>
rect 9 46 11 64
rect 36 49 38 57
rect 43 49 45 57
<< polycontact >>
rect 21 64 25 68
rect 13 38 17 42
rect 33 41 37 45
rect 43 41 47 45
rect 24 25 28 29
<< ndcontact >>
rect 3 16 7 20
rect 20 16 24 20
rect 51 16 55 20
<< pdcontact >>
rect 3 55 7 59
rect 3 47 7 51
rect 13 59 17 63
rect 29 64 33 68
rect 51 50 55 54
<< psubstratepcontact >>
rect 52 4 56 8
<< nsubstratencontact >>
rect 52 64 56 68
<< psubstratepdiff >>
rect 51 8 57 9
rect 51 4 52 8
rect 56 4 57 8
rect 51 3 57 4
<< nsubstratendiff >>
rect 51 68 57 69
rect 51 64 52 68
rect 56 64 57 68
rect 51 63 57 64
<< labels >>
rlabel polysilicon 15 33 15 33 6 an
rlabel metal1 12 32 12 32 6 z
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 48 12 48 6 z
rlabel metal1 28 32 28 32 6 a
rlabel metal1 20 40 20 40 6 an
rlabel metal1 32 4 32 4 6 vss
rlabel metal1 36 36 36 36 6 a
rlabel metal1 32 68 32 68 6 vdd
rlabel metal1 53 36 53 36 6 an
<< end >>
