magic
tech scmos
timestamp 1179384962
<< checkpaint >>
rect -22 -25 62 105
<< ab >>
rect 0 0 40 80
<< pwell >>
rect -4 -7 44 36
<< nwell >>
rect -4 36 44 87
<< polysilicon >>
rect 9 61 11 65
rect 19 63 21 68
rect 29 63 31 68
rect 9 39 11 43
rect 19 39 21 50
rect 29 47 31 50
rect 29 46 35 47
rect 29 42 30 46
rect 34 42 35 46
rect 29 41 35 42
rect 9 38 15 39
rect 9 34 10 38
rect 14 34 15 38
rect 9 33 15 34
rect 19 38 25 39
rect 19 34 20 38
rect 24 34 25 38
rect 19 33 25 34
rect 9 28 11 33
rect 22 28 24 33
rect 29 28 31 41
rect 9 15 11 19
rect 22 12 24 17
rect 29 12 31 17
<< ndiffusion >>
rect 4 25 9 28
rect 2 24 9 25
rect 2 20 3 24
rect 7 20 9 24
rect 2 19 9 20
rect 11 19 22 28
rect 13 17 22 19
rect 24 17 29 28
rect 31 23 36 28
rect 31 22 38 23
rect 31 18 33 22
rect 37 18 38 22
rect 31 17 38 18
rect 13 12 20 17
rect 13 8 14 12
rect 18 8 20 12
rect 13 7 20 8
<< pdiffusion >>
rect 13 61 19 63
rect 4 56 9 61
rect 2 55 9 56
rect 2 51 3 55
rect 7 51 9 55
rect 2 48 9 51
rect 2 44 3 48
rect 7 44 9 48
rect 2 43 9 44
rect 11 60 19 61
rect 11 56 13 60
rect 17 56 19 60
rect 11 50 19 56
rect 21 62 29 63
rect 21 58 23 62
rect 27 58 29 62
rect 21 55 29 58
rect 21 51 23 55
rect 27 51 29 55
rect 21 50 29 51
rect 31 62 38 63
rect 31 58 33 62
rect 37 58 38 62
rect 31 50 38 58
rect 11 43 17 50
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect -2 68 42 78
rect 12 60 18 68
rect 12 56 13 60
rect 17 56 18 60
rect 23 62 27 63
rect 32 62 38 68
rect 32 58 33 62
rect 37 58 38 62
rect 2 55 7 56
rect 2 51 3 55
rect 23 55 27 58
rect 2 48 7 51
rect 2 44 3 48
rect 2 43 7 44
rect 10 51 23 53
rect 10 49 27 51
rect 2 25 6 43
rect 10 38 14 49
rect 25 42 30 46
rect 34 42 38 55
rect 17 34 20 38
rect 24 34 31 38
rect 10 30 14 34
rect 10 26 22 30
rect 2 24 7 25
rect 2 20 3 24
rect 7 20 14 23
rect 2 17 14 20
rect 18 22 22 26
rect 26 25 31 34
rect 18 18 33 22
rect 37 18 38 22
rect -2 8 14 12
rect 18 8 42 12
rect -2 2 42 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
<< ntransistor >>
rect 9 19 11 28
rect 22 17 24 28
rect 29 17 31 28
<< ptransistor >>
rect 9 43 11 61
rect 19 50 21 63
rect 29 50 31 63
<< polycontact >>
rect 30 42 34 46
rect 10 34 14 38
rect 20 34 24 38
<< ndcontact >>
rect 3 20 7 24
rect 33 18 37 22
rect 14 8 18 12
<< pdcontact >>
rect 3 51 7 55
rect 3 44 7 48
rect 13 56 17 60
rect 23 58 27 62
rect 23 51 27 55
rect 33 58 37 62
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
<< psubstratepdiff >>
rect 0 2 40 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 40 2
rect 0 -3 40 -2
<< nsubstratendiff >>
rect 0 82 40 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 40 82
rect 0 77 40 78
<< labels >>
rlabel polycontact 12 36 12 36 6 zn
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 20 12 20 6 z
rlabel metal1 12 39 12 39 6 zn
rlabel metal1 20 6 20 6 6 vss
rlabel metal1 20 36 20 36 6 a
rlabel metal1 28 32 28 32 6 a
rlabel metal1 28 44 28 44 6 b
rlabel metal1 25 56 25 56 6 zn
rlabel metal1 20 74 20 74 6 vdd
rlabel metal1 28 20 28 20 6 zn
rlabel metal1 36 52 36 52 6 b
<< end >>
