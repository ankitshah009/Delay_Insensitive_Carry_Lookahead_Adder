magic
tech scmos
timestamp 1185094666
<< checkpaint >>
rect -22 -22 72 122
<< ab >>
rect 0 0 50 100
<< pwell >>
rect -4 -4 54 48
<< nwell >>
rect -4 48 54 104
<< polysilicon >>
rect 13 94 15 98
rect 25 94 27 98
rect 37 94 39 98
rect 13 43 15 56
rect 25 43 27 56
rect 37 53 39 56
rect 32 52 39 53
rect 32 48 33 52
rect 37 48 39 52
rect 32 47 39 48
rect 13 42 27 43
rect 13 38 22 42
rect 26 38 27 42
rect 13 37 27 38
rect 13 34 15 37
rect 25 34 27 37
rect 37 34 39 47
rect 13 11 15 15
rect 25 10 27 15
rect 37 10 39 15
<< ndiffusion >>
rect 4 22 13 34
rect 4 18 6 22
rect 10 18 13 22
rect 4 15 13 18
rect 15 32 25 34
rect 15 28 18 32
rect 22 28 25 32
rect 15 22 25 28
rect 15 18 18 22
rect 22 18 25 22
rect 15 15 25 18
rect 27 32 37 34
rect 27 28 30 32
rect 34 28 37 32
rect 27 22 37 28
rect 27 18 30 22
rect 34 18 37 22
rect 27 15 37 18
rect 39 33 47 34
rect 39 29 42 33
rect 46 29 47 33
rect 39 25 47 29
rect 39 21 42 25
rect 46 21 47 25
rect 39 20 47 21
rect 39 15 44 20
<< pdiffusion >>
rect 4 92 13 94
rect 4 88 6 92
rect 10 88 13 92
rect 4 82 13 88
rect 4 78 6 82
rect 10 78 13 82
rect 4 72 13 78
rect 4 68 6 72
rect 10 68 13 72
rect 4 56 13 68
rect 15 72 25 94
rect 15 68 18 72
rect 22 68 25 72
rect 15 62 25 68
rect 15 58 18 62
rect 22 58 25 62
rect 15 56 25 58
rect 27 92 37 94
rect 27 88 30 92
rect 34 88 37 92
rect 27 82 37 88
rect 27 78 30 82
rect 34 78 37 82
rect 27 56 37 78
rect 39 70 44 94
rect 39 69 47 70
rect 39 65 42 69
rect 46 65 47 69
rect 39 61 47 65
rect 39 57 42 61
rect 46 57 47 61
rect 39 56 47 57
<< metal1 >>
rect -2 92 52 100
rect -2 88 6 92
rect 10 88 30 92
rect 34 88 52 92
rect 6 82 10 88
rect 6 72 10 78
rect 30 82 34 88
rect 30 77 34 78
rect 6 67 10 68
rect 18 72 22 73
rect 18 63 22 68
rect 8 62 22 63
rect 8 58 18 62
rect 8 57 22 58
rect 8 33 12 57
rect 28 52 32 73
rect 42 69 46 70
rect 42 61 46 65
rect 17 48 33 52
rect 37 48 38 52
rect 42 42 46 57
rect 21 38 22 42
rect 26 38 46 42
rect 42 33 46 38
rect 8 32 22 33
rect 8 28 18 32
rect 8 27 22 28
rect 6 22 10 23
rect 6 12 10 18
rect 18 22 22 27
rect 18 17 22 18
rect 30 32 34 33
rect 30 22 34 28
rect 42 25 46 29
rect 42 20 46 21
rect 30 12 34 18
rect -2 8 52 12
rect -2 4 8 8
rect 12 4 18 8
rect 22 4 52 8
rect -2 0 52 4
<< ntransistor >>
rect 13 15 15 34
rect 25 15 27 34
rect 37 15 39 34
<< ptransistor >>
rect 13 56 15 94
rect 25 56 27 94
rect 37 56 39 94
<< polycontact >>
rect 33 48 37 52
rect 22 38 26 42
<< ndcontact >>
rect 6 18 10 22
rect 18 28 22 32
rect 18 18 22 22
rect 30 28 34 32
rect 30 18 34 22
rect 42 29 46 33
rect 42 21 46 25
<< pdcontact >>
rect 6 88 10 92
rect 6 78 10 82
rect 6 68 10 72
rect 18 68 22 72
rect 18 58 22 62
rect 30 88 34 92
rect 30 78 34 82
rect 42 65 46 69
rect 42 57 46 61
<< psubstratepcontact >>
rect 8 4 12 8
rect 18 4 22 8
<< psubstratepdiff >>
rect 7 8 23 9
rect 7 4 8 8
rect 12 4 18 8
rect 22 4 23 8
rect 7 3 23 4
<< labels >>
rlabel polysilicon 20 40 20 40 6 an
rlabel metal1 20 25 20 25 6 z
rlabel metal1 10 45 10 45 6 z
rlabel metal1 20 50 20 50 6 a
rlabel metal1 20 65 20 65 6 z
rlabel metal1 25 6 25 6 6 vss
rlabel metal1 30 60 30 60 6 a
rlabel metal1 25 94 25 94 6 vdd
rlabel metal1 33 40 33 40 6 an
rlabel metal1 44 45 44 45 6 an
<< end >>
