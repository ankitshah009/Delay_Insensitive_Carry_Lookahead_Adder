magic
tech scmos
timestamp 1179385404
<< checkpaint >>
rect -22 -25 78 105
<< ab >>
rect 0 0 56 80
<< pwell >>
rect -4 -7 60 36
<< nwell >>
rect -4 36 60 87
<< polysilicon >>
rect 31 66 33 71
rect 41 66 43 71
rect 9 57 11 62
rect 19 57 21 62
rect 31 48 33 51
rect 31 47 37 48
rect 31 43 32 47
rect 36 43 37 47
rect 9 38 11 43
rect 19 40 21 43
rect 31 42 37 43
rect 19 39 27 40
rect 19 38 22 39
rect 9 37 15 38
rect 9 33 10 37
rect 14 34 15 37
rect 21 35 22 38
rect 26 35 27 39
rect 21 34 27 35
rect 14 33 17 34
rect 9 32 17 33
rect 15 29 17 32
rect 22 29 24 34
rect 34 30 36 42
rect 41 39 43 51
rect 41 38 47 39
rect 41 34 42 38
rect 46 34 47 38
rect 41 33 47 34
rect 41 30 43 33
rect 15 12 17 17
rect 22 12 24 17
rect 34 12 36 17
rect 41 12 43 17
<< ndiffusion >>
rect 26 29 34 30
rect 10 23 15 29
rect 8 22 15 23
rect 8 18 9 22
rect 13 18 15 22
rect 8 17 15 18
rect 17 17 22 29
rect 24 17 34 29
rect 36 17 41 30
rect 43 23 48 30
rect 43 22 50 23
rect 43 18 45 22
rect 49 18 50 22
rect 43 17 50 18
rect 26 12 32 17
rect 26 8 27 12
rect 31 8 32 12
rect 26 7 32 8
<< pdiffusion >>
rect 23 72 29 73
rect 23 68 24 72
rect 28 68 29 72
rect 23 66 29 68
rect 23 57 31 66
rect 2 56 9 57
rect 2 52 3 56
rect 7 52 9 56
rect 2 43 9 52
rect 11 55 19 57
rect 11 51 13 55
rect 17 51 19 55
rect 11 48 19 51
rect 11 44 13 48
rect 17 44 19 48
rect 11 43 19 44
rect 21 51 31 57
rect 33 62 41 66
rect 33 58 35 62
rect 39 58 41 62
rect 33 51 41 58
rect 43 65 50 66
rect 43 61 45 65
rect 49 61 50 65
rect 43 57 50 61
rect 43 53 45 57
rect 49 53 50 57
rect 43 51 50 53
rect 21 43 29 51
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect -2 72 58 78
rect -2 68 24 72
rect 28 68 58 72
rect 3 56 7 68
rect 45 65 49 68
rect 23 58 35 62
rect 39 58 40 62
rect 3 51 7 52
rect 13 55 17 56
rect 13 48 17 51
rect 2 44 13 47
rect 2 43 17 44
rect 2 23 6 43
rect 23 39 27 58
rect 45 57 49 61
rect 33 48 39 54
rect 45 52 49 53
rect 32 47 39 48
rect 36 46 39 47
rect 36 43 47 46
rect 32 42 47 43
rect 10 37 14 39
rect 19 35 22 39
rect 10 31 14 33
rect 10 27 22 31
rect 2 22 14 23
rect 2 18 9 22
rect 13 18 14 22
rect 2 17 14 18
rect 18 17 22 27
rect 26 22 30 39
rect 34 34 42 38
rect 46 34 47 38
rect 34 25 38 34
rect 26 18 45 22
rect 49 18 50 22
rect -2 8 27 12
rect 31 8 58 12
rect -2 2 58 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
<< ntransistor >>
rect 15 17 17 29
rect 22 17 24 29
rect 34 17 36 30
rect 41 17 43 30
<< ptransistor >>
rect 9 43 11 57
rect 19 43 21 57
rect 31 51 33 66
rect 41 51 43 66
<< polycontact >>
rect 32 43 36 47
rect 10 33 14 37
rect 22 35 26 39
rect 42 34 46 38
<< ndcontact >>
rect 9 18 13 22
rect 45 18 49 22
rect 27 8 31 12
<< pdcontact >>
rect 24 68 28 72
rect 3 52 7 56
rect 13 51 17 55
rect 13 44 17 48
rect 35 58 39 62
rect 45 61 49 65
rect 45 53 49 57
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
<< psubstratepdiff >>
rect 0 2 56 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 56 2
rect 0 -3 56 -2
<< nsubstratendiff >>
rect 0 82 56 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 56 82
rect 0 77 56 78
<< labels >>
rlabel polycontact 24 37 24 37 6 an
rlabel metal1 4 32 4 32 6 z
rlabel ndcontact 12 20 12 20 6 z
rlabel polycontact 12 36 12 36 6 b
rlabel metal1 20 24 20 24 6 b
rlabel metal1 28 6 28 6 6 vss
rlabel polycontact 24 37 24 37 6 an
rlabel metal1 36 28 36 28 6 a1
rlabel metal1 36 48 36 48 6 a2
rlabel metal1 31 60 31 60 6 an
rlabel metal1 28 74 28 74 6 vdd
rlabel metal1 38 20 38 20 6 an
rlabel polycontact 44 36 44 36 6 a1
rlabel metal1 44 44 44 44 6 a2
<< end >>
