magic
tech scmos
timestamp 1179385095
<< checkpaint >>
rect -22 -22 78 94
<< ab >>
rect 0 0 56 72
<< pwell >>
rect -4 -4 60 32
<< nwell >>
rect -4 32 60 76
<< polysilicon >>
rect 9 60 11 65
rect 19 60 21 65
rect 29 60 31 65
rect 41 60 43 65
rect 19 43 21 54
rect 29 51 31 54
rect 29 50 37 51
rect 29 46 32 50
rect 36 46 37 50
rect 29 45 37 46
rect 19 42 25 43
rect 9 35 11 42
rect 19 38 20 42
rect 24 38 25 42
rect 19 37 25 38
rect 9 34 15 35
rect 9 30 10 34
rect 14 30 15 34
rect 9 29 15 30
rect 9 22 11 29
rect 22 19 24 37
rect 29 19 31 45
rect 41 28 43 54
rect 40 27 46 28
rect 40 24 41 27
rect 36 23 41 24
rect 45 23 46 27
rect 36 22 46 23
rect 36 19 38 22
rect 9 8 11 13
rect 22 8 24 13
rect 29 8 31 13
rect 36 8 38 13
<< ndiffusion >>
rect 4 19 9 22
rect 2 18 9 19
rect 2 14 3 18
rect 7 14 9 18
rect 2 13 9 14
rect 11 19 20 22
rect 11 13 22 19
rect 24 13 29 19
rect 31 13 36 19
rect 38 18 45 19
rect 38 14 40 18
rect 44 14 45 18
rect 38 13 45 14
rect 13 8 20 13
rect 13 4 14 8
rect 18 4 20 8
rect 13 3 20 4
<< pdiffusion >>
rect 33 68 39 69
rect 33 64 34 68
rect 38 64 39 68
rect 33 60 39 64
rect 4 55 9 60
rect 2 54 9 55
rect 2 50 3 54
rect 7 50 9 54
rect 2 47 9 50
rect 2 43 3 47
rect 7 43 9 47
rect 2 42 9 43
rect 11 59 19 60
rect 11 55 13 59
rect 17 55 19 59
rect 11 54 19 55
rect 21 59 29 60
rect 21 55 23 59
rect 27 55 29 59
rect 21 54 29 55
rect 31 54 41 60
rect 43 59 50 60
rect 43 55 45 59
rect 49 55 50 59
rect 43 54 50 55
rect 11 42 17 54
<< metal1 >>
rect -2 68 58 72
rect -2 64 34 68
rect 38 64 58 68
rect 13 59 17 64
rect 2 54 7 59
rect 13 54 17 55
rect 22 55 23 59
rect 27 55 45 59
rect 49 55 50 59
rect 2 50 3 54
rect 22 50 26 55
rect 2 47 7 50
rect 2 43 3 47
rect 2 42 7 43
rect 10 46 26 50
rect 31 46 32 50
rect 36 46 47 50
rect 2 18 6 42
rect 10 34 14 46
rect 17 38 20 42
rect 24 38 31 42
rect 41 38 47 46
rect 25 30 31 38
rect 10 26 14 30
rect 41 27 47 34
rect 10 22 22 26
rect 25 23 41 26
rect 45 23 47 27
rect 25 22 47 23
rect 18 18 22 22
rect 2 14 3 18
rect 7 14 15 18
rect 18 14 40 18
rect 44 14 45 18
rect -2 4 14 8
rect 18 4 58 8
rect -2 0 58 4
<< ntransistor >>
rect 9 13 11 22
rect 22 13 24 19
rect 29 13 31 19
rect 36 13 38 19
<< ptransistor >>
rect 9 42 11 60
rect 19 54 21 60
rect 29 54 31 60
rect 41 54 43 60
<< polycontact >>
rect 32 46 36 50
rect 20 38 24 42
rect 10 30 14 34
rect 41 23 45 27
<< ndcontact >>
rect 3 14 7 18
rect 40 14 44 18
rect 14 4 18 8
<< pdcontact >>
rect 34 64 38 68
rect 3 50 7 54
rect 3 43 7 47
rect 13 55 17 59
rect 23 55 27 59
rect 45 55 49 59
<< labels >>
rlabel polycontact 12 32 12 32 6 zn
rlabel metal1 4 40 4 40 6 z
rlabel metal1 12 16 12 16 6 z
rlabel metal1 20 40 20 40 6 a
rlabel metal1 12 36 12 36 6 zn
rlabel metal1 28 4 28 4 6 vss
rlabel metal1 28 24 28 24 6 c
rlabel metal1 36 24 36 24 6 c
rlabel metal1 28 36 28 36 6 a
rlabel metal1 36 48 36 48 6 b
rlabel metal1 28 68 28 68 6 vdd
rlabel metal1 31 16 31 16 6 zn
rlabel metal1 44 28 44 28 6 c
rlabel metal1 44 44 44 44 6 b
rlabel metal1 36 57 36 57 6 zn
<< end >>
