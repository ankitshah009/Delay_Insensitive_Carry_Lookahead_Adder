magic
tech scmos
timestamp 1180600647
<< checkpaint >>
rect -22 -22 232 122
<< ab >>
rect 0 0 210 100
<< pwell >>
rect -4 -4 214 48
<< nwell >>
rect -4 48 214 104
<< polysilicon >>
rect 81 94 83 98
rect 93 94 95 98
rect 105 94 107 98
rect 117 94 119 98
rect 11 83 13 87
rect 23 83 25 87
rect 35 83 37 87
rect 47 83 49 87
rect 57 83 59 87
rect 11 43 13 65
rect 23 43 25 65
rect 35 53 37 65
rect 7 42 13 43
rect 7 38 8 42
rect 12 38 13 42
rect 7 37 13 38
rect 17 42 25 43
rect 17 38 18 42
rect 22 38 25 42
rect 17 37 25 38
rect 33 52 43 53
rect 33 48 38 52
rect 42 48 43 52
rect 33 47 43 48
rect 11 27 13 37
rect 21 29 23 37
rect 33 25 35 47
rect 47 43 49 57
rect 57 53 59 57
rect 131 83 133 87
rect 143 83 145 87
rect 153 83 155 87
rect 165 84 167 88
rect 57 52 63 53
rect 57 48 58 52
rect 62 48 63 52
rect 57 47 63 48
rect 47 42 53 43
rect 47 39 48 42
rect 45 38 48 39
rect 52 38 53 42
rect 45 37 53 38
rect 45 25 47 37
rect 57 25 59 47
rect 81 43 83 55
rect 93 43 95 55
rect 75 42 95 43
rect 75 38 76 42
rect 80 38 95 42
rect 75 37 95 38
rect 81 25 83 37
rect 93 25 95 37
rect 105 43 107 55
rect 117 43 119 55
rect 131 43 133 69
rect 143 67 145 70
rect 153 67 155 70
rect 141 65 145 67
rect 151 65 155 67
rect 177 79 179 83
rect 187 79 189 83
rect 197 79 199 83
rect 141 43 143 65
rect 151 43 153 65
rect 165 63 167 66
rect 163 61 167 63
rect 163 43 165 61
rect 177 53 179 65
rect 187 53 189 65
rect 177 52 183 53
rect 177 49 178 52
rect 105 42 123 43
rect 105 38 118 42
rect 122 38 123 42
rect 105 37 123 38
rect 127 42 133 43
rect 127 38 128 42
rect 132 38 133 42
rect 127 37 133 38
rect 137 42 143 43
rect 137 38 138 42
rect 142 38 143 42
rect 137 37 143 38
rect 147 42 153 43
rect 147 38 148 42
rect 152 38 153 42
rect 147 37 153 38
rect 157 42 165 43
rect 157 38 158 42
rect 162 38 165 42
rect 157 37 165 38
rect 105 25 107 37
rect 117 25 119 37
rect 131 25 133 37
rect 141 25 143 37
rect 151 25 153 37
rect 163 27 165 37
rect 175 48 178 49
rect 182 48 183 52
rect 175 47 183 48
rect 187 52 193 53
rect 187 48 188 52
rect 192 48 193 52
rect 187 47 193 48
rect 11 13 13 17
rect 21 13 23 17
rect 33 13 35 17
rect 45 13 47 17
rect 57 13 59 17
rect 175 25 177 47
rect 187 29 189 47
rect 185 27 189 29
rect 197 43 199 65
rect 197 42 203 43
rect 197 38 198 42
rect 202 38 203 42
rect 197 37 203 38
rect 185 24 187 27
rect 197 25 199 37
rect 131 13 133 17
rect 141 13 143 17
rect 151 13 153 17
rect 163 13 165 17
rect 175 13 177 17
rect 185 13 187 17
rect 197 13 199 17
rect 81 2 83 6
rect 93 2 95 6
rect 105 2 107 6
rect 117 2 119 6
<< ndiffusion >>
rect 16 27 21 29
rect 3 17 11 27
rect 13 17 21 27
rect 23 25 31 29
rect 158 25 163 27
rect 23 22 33 25
rect 23 18 26 22
rect 30 18 33 22
rect 23 17 33 18
rect 35 22 45 25
rect 35 18 38 22
rect 42 18 45 22
rect 35 17 45 18
rect 47 17 57 25
rect 59 22 67 25
rect 59 18 62 22
rect 66 18 67 22
rect 59 17 67 18
rect 73 22 81 25
rect 73 18 74 22
rect 78 18 81 22
rect 3 12 9 17
rect 3 8 4 12
rect 8 8 9 12
rect 49 12 55 17
rect 3 7 9 8
rect 49 8 50 12
rect 54 8 55 12
rect 49 7 55 8
rect 73 12 81 18
rect 73 8 74 12
rect 78 8 81 12
rect 73 6 81 8
rect 83 22 93 25
rect 83 18 86 22
rect 90 18 93 22
rect 83 6 93 18
rect 95 12 105 25
rect 95 8 98 12
rect 102 8 105 12
rect 95 6 105 8
rect 107 22 117 25
rect 107 18 110 22
rect 114 18 117 22
rect 107 6 117 18
rect 119 17 131 25
rect 133 17 141 25
rect 143 17 151 25
rect 153 22 163 25
rect 153 18 156 22
rect 160 18 163 22
rect 153 17 163 18
rect 165 25 170 27
rect 165 22 175 25
rect 165 18 168 22
rect 172 18 175 22
rect 165 17 175 18
rect 177 24 182 25
rect 192 24 197 25
rect 177 17 185 24
rect 187 22 197 24
rect 187 18 190 22
rect 194 18 197 22
rect 187 17 197 18
rect 199 22 207 25
rect 199 18 202 22
rect 206 18 207 22
rect 199 17 207 18
rect 119 12 129 17
rect 119 8 122 12
rect 126 8 129 12
rect 179 11 183 17
rect 119 6 129 8
rect 178 10 184 11
rect 178 6 179 10
rect 183 6 184 10
rect 178 5 184 6
<< pdiffusion >>
rect 15 92 21 93
rect 15 88 16 92
rect 20 88 21 92
rect 146 94 152 95
rect 73 92 81 94
rect 15 83 21 88
rect 73 88 74 92
rect 78 88 81 92
rect 3 82 11 83
rect 3 78 4 82
rect 8 78 11 82
rect 3 65 11 78
rect 13 65 23 83
rect 25 82 35 83
rect 25 78 28 82
rect 32 78 35 82
rect 25 65 35 78
rect 37 72 47 83
rect 37 68 40 72
rect 44 68 47 72
rect 37 65 47 68
rect 40 57 47 65
rect 49 57 57 83
rect 59 82 67 83
rect 59 78 62 82
rect 66 78 67 82
rect 59 57 67 78
rect 73 55 81 88
rect 83 72 93 94
rect 83 68 86 72
rect 90 68 93 72
rect 83 62 93 68
rect 83 58 86 62
rect 90 58 93 62
rect 83 55 93 58
rect 95 92 105 94
rect 95 88 98 92
rect 102 88 105 92
rect 95 55 105 88
rect 107 72 117 94
rect 107 68 110 72
rect 114 68 117 72
rect 107 62 117 68
rect 107 58 110 62
rect 114 58 117 62
rect 107 55 117 58
rect 119 92 129 94
rect 119 88 122 92
rect 126 88 129 92
rect 146 90 147 94
rect 151 90 152 94
rect 146 89 152 90
rect 119 83 129 88
rect 147 83 151 89
rect 157 83 165 84
rect 119 69 131 83
rect 133 82 143 83
rect 133 78 136 82
rect 140 78 143 82
rect 133 70 143 78
rect 145 70 153 83
rect 155 82 165 83
rect 155 78 158 82
rect 162 78 165 82
rect 155 70 165 78
rect 133 69 138 70
rect 119 55 127 69
rect 157 66 165 70
rect 167 79 174 84
rect 201 82 207 83
rect 201 79 202 82
rect 167 72 177 79
rect 167 68 170 72
rect 174 68 177 72
rect 167 66 177 68
rect 172 65 177 66
rect 179 65 187 79
rect 189 65 197 79
rect 199 78 202 79
rect 206 78 207 82
rect 199 65 207 78
<< metal1 >>
rect -2 96 212 100
rect -2 92 30 96
rect 34 92 38 96
rect 42 92 46 96
rect 50 92 54 96
rect 58 92 62 96
rect 66 94 160 96
rect 66 92 147 94
rect -2 88 16 92
rect 20 88 74 92
rect 78 88 98 92
rect 102 88 122 92
rect 126 90 147 92
rect 151 92 160 94
rect 164 92 168 96
rect 172 92 176 96
rect 180 92 184 96
rect 188 92 192 96
rect 196 92 212 96
rect 151 90 212 92
rect 126 88 212 90
rect 3 78 4 82
rect 8 78 28 82
rect 32 78 62 82
rect 66 78 67 82
rect 74 78 124 82
rect 135 78 136 82
rect 140 78 158 82
rect 162 78 202 82
rect 206 78 207 82
rect 8 42 12 73
rect 8 17 12 38
rect 18 42 22 73
rect 74 72 78 78
rect 88 72 92 73
rect 18 27 22 38
rect 28 68 40 72
rect 44 68 78 72
rect 85 68 86 72
rect 90 68 92 72
rect 28 22 32 68
rect 38 52 42 63
rect 38 27 42 48
rect 48 42 52 63
rect 48 27 52 38
rect 58 52 62 63
rect 58 27 62 48
rect 74 42 78 68
rect 88 62 92 68
rect 85 58 86 62
rect 90 58 92 62
rect 74 38 76 42
rect 80 38 81 42
rect 74 22 78 23
rect 88 22 92 58
rect 25 18 26 22
rect 30 18 32 22
rect 37 18 38 22
rect 42 18 62 22
rect 66 18 67 22
rect 85 18 86 22
rect 90 18 92 22
rect 74 12 78 18
rect 88 17 92 18
rect 108 72 112 73
rect 120 72 124 78
rect 168 72 172 73
rect 108 68 110 72
rect 114 68 115 72
rect 120 68 162 72
rect 108 62 112 68
rect 108 58 110 62
rect 114 58 115 62
rect 108 22 112 58
rect 118 42 122 43
rect 118 32 122 38
rect 128 42 132 63
rect 128 37 132 38
rect 138 42 142 63
rect 118 28 132 32
rect 128 22 132 28
rect 138 27 142 38
rect 148 42 152 63
rect 148 27 152 38
rect 158 42 162 68
rect 158 37 162 38
rect 168 68 170 72
rect 174 68 175 72
rect 168 32 172 68
rect 158 28 172 32
rect 178 52 182 63
rect 158 22 162 28
rect 178 27 182 48
rect 188 52 192 73
rect 188 27 192 48
rect 198 42 202 73
rect 198 27 202 38
rect 202 22 206 23
rect 108 18 110 22
rect 114 18 115 22
rect 128 18 156 22
rect 160 18 162 22
rect 167 18 168 22
rect 172 18 190 22
rect 194 18 195 22
rect 108 17 112 18
rect 158 17 162 18
rect 202 12 206 18
rect -2 8 4 12
rect 8 10 50 12
rect 8 8 18 10
rect -2 6 18 8
rect 22 6 28 10
rect 32 6 38 10
rect 42 8 50 10
rect 54 8 74 12
rect 78 8 98 12
rect 102 8 122 12
rect 126 10 212 12
rect 126 8 136 10
rect 42 6 136 8
rect 140 6 146 10
rect 150 6 156 10
rect 160 6 167 10
rect 171 6 179 10
rect 183 6 192 10
rect 196 6 200 10
rect 204 6 212 10
rect -2 0 212 6
<< ntransistor >>
rect 11 17 13 27
rect 21 17 23 29
rect 33 17 35 25
rect 45 17 47 25
rect 57 17 59 25
rect 81 6 83 25
rect 93 6 95 25
rect 105 6 107 25
rect 117 6 119 25
rect 131 17 133 25
rect 141 17 143 25
rect 151 17 153 25
rect 163 17 165 27
rect 175 17 177 25
rect 185 17 187 24
rect 197 17 199 25
<< ptransistor >>
rect 11 65 13 83
rect 23 65 25 83
rect 35 65 37 83
rect 47 57 49 83
rect 57 57 59 83
rect 81 55 83 94
rect 93 55 95 94
rect 105 55 107 94
rect 117 55 119 94
rect 131 69 133 83
rect 143 70 145 83
rect 153 70 155 83
rect 165 66 167 84
rect 177 65 179 79
rect 187 65 189 79
rect 197 65 199 79
<< polycontact >>
rect 8 38 12 42
rect 18 38 22 42
rect 38 48 42 52
rect 58 48 62 52
rect 48 38 52 42
rect 76 38 80 42
rect 118 38 122 42
rect 128 38 132 42
rect 138 38 142 42
rect 148 38 152 42
rect 158 38 162 42
rect 178 48 182 52
rect 188 48 192 52
rect 198 38 202 42
<< ndcontact >>
rect 26 18 30 22
rect 38 18 42 22
rect 62 18 66 22
rect 74 18 78 22
rect 4 8 8 12
rect 50 8 54 12
rect 74 8 78 12
rect 86 18 90 22
rect 98 8 102 12
rect 110 18 114 22
rect 156 18 160 22
rect 168 18 172 22
rect 190 18 194 22
rect 202 18 206 22
rect 122 8 126 12
rect 179 6 183 10
<< pdcontact >>
rect 16 88 20 92
rect 74 88 78 92
rect 4 78 8 82
rect 28 78 32 82
rect 40 68 44 72
rect 62 78 66 82
rect 86 68 90 72
rect 86 58 90 62
rect 98 88 102 92
rect 110 68 114 72
rect 110 58 114 62
rect 122 88 126 92
rect 147 90 151 94
rect 136 78 140 82
rect 158 78 162 82
rect 170 68 174 72
rect 202 78 206 82
<< psubstratepcontact >>
rect 18 6 22 10
rect 28 6 32 10
rect 38 6 42 10
rect 136 6 140 10
rect 146 6 150 10
rect 156 6 160 10
rect 167 6 171 10
rect 192 6 196 10
rect 200 6 204 10
<< nsubstratencontact >>
rect 30 92 34 96
rect 38 92 42 96
rect 46 92 50 96
rect 54 92 58 96
rect 62 92 66 96
rect 160 92 164 96
rect 168 92 172 96
rect 176 92 180 96
rect 184 92 188 96
rect 192 92 196 96
<< psubstratepdiff >>
rect 17 10 43 11
rect 17 6 18 10
rect 22 6 28 10
rect 32 6 38 10
rect 42 6 43 10
rect 135 10 172 11
rect 135 6 136 10
rect 140 6 146 10
rect 150 6 156 10
rect 160 6 167 10
rect 171 6 172 10
rect 17 5 43 6
rect 135 5 172 6
rect 191 10 205 11
rect 191 6 192 10
rect 196 6 200 10
rect 204 6 205 10
rect 191 5 205 6
<< nsubstratendiff >>
rect 29 96 67 97
rect 29 92 30 96
rect 34 92 38 96
rect 42 92 46 96
rect 50 92 54 96
rect 58 92 62 96
rect 66 92 67 96
rect 159 96 197 97
rect 29 91 67 92
rect 159 92 160 96
rect 164 92 168 96
rect 172 92 176 96
rect 180 92 184 96
rect 188 92 192 96
rect 196 92 197 96
rect 159 91 197 92
<< labels >>
rlabel metal1 20 50 20 50 6 b1
rlabel metal1 10 45 10 45 6 a1
rlabel metal1 40 45 40 45 6 cin1
rlabel metal1 50 45 50 45 6 a2
rlabel metal1 60 45 60 45 6 b2
rlabel metal1 105 6 105 6 6 vss
rlabel metal1 90 45 90 45 6 cout
rlabel metal1 110 45 110 45 6 sout
rlabel metal1 105 94 105 94 6 vdd
rlabel metal1 130 50 130 50 6 a3
rlabel metal1 140 45 140 45 6 b3
rlabel metal1 150 45 150 45 6 cin2
rlabel metal1 200 50 200 50 6 b4
rlabel polycontact 190 50 190 50 6 a4
rlabel metal1 180 45 180 45 6 cin3
<< end >>
