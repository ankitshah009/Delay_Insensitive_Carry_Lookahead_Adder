.subckt iv1v0x6 a vdd vss z
*   SPICE3 file   created from iv1v0x6.ext -      technology: scmos
m00 vdd    vdd    w1     vdd p w=28u  l=2.3636u ad=186p     pd=60u      as=196p     ps=70u
m01 z      a      vdd    vdd p w=28u  l=2.3636u ad=182.667p pd=56.6667u as=186p     ps=60u
m02 z      a      vdd    vdd p w=28u  l=2.3636u ad=182.667p pd=56.6667u as=186p     ps=60u
m03 vdd    a      z      vdd p w=28u  l=2.3636u ad=186p     pd=60u      as=182.667p ps=56.6667u
m04 vss    vdd    w2     vss n w=20u  l=2.3636u ad=138p     pd=48u      as=140p     ps=54u
m05 z      a      vss    vss n w=20u  l=2.3636u ad=137.333p pd=46u      as=138p     ps=48u
m06 z      a      vss    vss n w=20u  l=2.3636u ad=137.333p pd=46u      as=138p     ps=48u
m07 vss    a      z      vss n w=20u  l=2.3636u ad=138p     pd=48u      as=137.333p ps=46u
C0  z      vdd    0.250f
C1  vss    z      0.237f
C2  vss    vdd    0.017f
C3  z      a      0.326f
C4  a      vdd    0.520f
C5  vss    a      0.099f
C7  z      vss    0.010f
C8  a      vss    0.144f
.ends
