.subckt inv_x8 i nq vdd vss
*   SPICE3 file   created from inv_x8.ext -      technology: scmos
m00 nq     i      vdd    vdd p w=39u  l=2.3636u ad=195p     pd=49u      as=237p     ps=71.5u
m01 vdd    i      nq     vdd p w=39u  l=2.3636u ad=237p     pd=71.5u    as=195p     ps=49u
m02 nq     i      vdd    vdd p w=39u  l=2.3636u ad=195p     pd=49u      as=237p     ps=71.5u
m03 vdd    i      nq     vdd p w=39u  l=2.3636u ad=237p     pd=71.5u    as=195p     ps=49u
m04 nq     i      vss    vss n w=18u  l=2.3636u ad=90p      pd=28u      as=117p     ps=40u
m05 vss    i      nq     vss n w=18u  l=2.3636u ad=117p     pd=40u      as=90p      ps=28u
m06 nq     i      vss    vss n w=18u  l=2.3636u ad=90p      pd=28u      as=117p     ps=40u
m07 vss    i      nq     vss n w=18u  l=2.3636u ad=117p     pd=40u      as=90p      ps=28u
C0  vss    nq     0.254f
C1  nq     vdd    0.399f
C2  vss    i      0.082f
C3  vdd    i      0.156f
C4  vss    vdd    0.024f
C5  nq     i      0.441f
C7  nq     vss    0.032f
C9  i      vss    0.123f
.ends
