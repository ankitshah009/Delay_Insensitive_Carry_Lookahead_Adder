magic
tech scmos
timestamp 1179385133
<< checkpaint >>
rect -22 -22 86 94
<< ab >>
rect 0 0 64 72
<< pwell >>
rect -4 -4 68 32
<< nwell >>
rect -4 32 68 76
<< polysilicon >>
rect 20 61 22 66
rect 30 61 32 66
rect 42 61 44 66
rect 52 61 54 66
rect 9 57 11 61
rect 9 35 11 39
rect 20 35 22 48
rect 30 45 32 48
rect 30 44 37 45
rect 30 40 32 44
rect 36 40 37 44
rect 30 39 37 40
rect 42 43 44 48
rect 42 42 48 43
rect 9 34 15 35
rect 9 30 10 34
rect 14 30 15 34
rect 9 29 15 30
rect 20 34 26 35
rect 20 30 21 34
rect 25 30 26 34
rect 20 29 26 30
rect 9 24 11 29
rect 24 24 26 29
rect 31 24 33 39
rect 42 38 43 42
rect 47 38 48 42
rect 42 37 48 38
rect 42 35 44 37
rect 38 33 44 35
rect 52 35 54 48
rect 52 34 58 35
rect 38 24 40 33
rect 52 30 53 34
rect 57 30 58 34
rect 52 29 58 30
rect 45 27 58 29
rect 45 24 47 27
rect 9 11 11 15
rect 24 3 26 8
rect 31 3 33 8
rect 38 3 40 8
rect 45 3 47 8
<< ndiffusion >>
rect 4 21 9 24
rect 2 20 9 21
rect 2 16 3 20
rect 7 16 9 20
rect 2 15 9 16
rect 11 15 24 24
rect 13 8 24 15
rect 26 8 31 24
rect 33 8 38 24
rect 40 8 45 24
rect 47 18 52 24
rect 47 17 54 18
rect 47 13 49 17
rect 53 13 54 17
rect 47 12 54 13
rect 47 8 52 12
rect 13 4 15 8
rect 19 4 22 8
rect 13 3 22 4
<< pdiffusion >>
rect 34 68 40 69
rect 34 64 35 68
rect 39 64 40 68
rect 34 61 40 64
rect 13 59 20 61
rect 13 57 14 59
rect 4 52 9 57
rect 2 51 9 52
rect 2 47 3 51
rect 7 47 9 51
rect 2 44 9 47
rect 2 40 3 44
rect 7 40 9 44
rect 2 39 9 40
rect 11 55 14 57
rect 18 55 20 59
rect 11 48 20 55
rect 22 59 30 61
rect 22 55 24 59
rect 28 55 30 59
rect 22 48 30 55
rect 32 48 42 61
rect 44 59 52 61
rect 44 55 46 59
rect 50 55 52 59
rect 44 48 52 55
rect 54 60 61 61
rect 54 56 56 60
rect 60 56 61 60
rect 54 53 61 56
rect 54 49 56 53
rect 60 49 61 53
rect 54 48 61 49
rect 11 39 18 48
<< metal1 >>
rect -2 68 66 72
rect -2 64 4 68
rect 8 64 35 68
rect 39 64 66 68
rect 14 59 18 64
rect 56 60 60 64
rect 2 51 7 59
rect 14 54 18 55
rect 22 55 24 59
rect 28 55 46 59
rect 50 55 51 59
rect 2 47 3 51
rect 22 50 26 55
rect 56 53 60 56
rect 2 44 7 47
rect 2 40 3 44
rect 2 39 7 40
rect 12 46 26 50
rect 2 21 6 39
rect 12 35 16 46
rect 34 44 38 51
rect 25 40 32 42
rect 36 40 38 44
rect 25 38 38 40
rect 42 42 46 51
rect 56 48 60 49
rect 42 38 43 42
rect 47 38 55 42
rect 10 34 16 35
rect 14 30 16 34
rect 20 30 21 34
rect 25 30 31 34
rect 41 30 53 34
rect 57 30 62 34
rect 10 29 16 30
rect 12 26 16 29
rect 27 26 31 30
rect 12 22 23 26
rect 27 22 47 26
rect 2 20 7 21
rect 2 16 3 20
rect 7 16 15 18
rect 2 13 15 16
rect 19 17 23 22
rect 19 13 49 17
rect 53 13 54 17
rect 58 13 62 30
rect -2 4 4 8
rect 8 4 15 8
rect 19 4 66 8
rect -2 0 66 4
<< ntransistor >>
rect 9 15 11 24
rect 24 8 26 24
rect 31 8 33 24
rect 38 8 40 24
rect 45 8 47 24
<< ptransistor >>
rect 9 39 11 57
rect 20 48 22 61
rect 30 48 32 61
rect 42 48 44 61
rect 52 48 54 61
<< polycontact >>
rect 32 40 36 44
rect 10 30 14 34
rect 21 30 25 34
rect 43 38 47 42
rect 53 30 57 34
<< ndcontact >>
rect 3 16 7 20
rect 49 13 53 17
rect 15 4 19 8
<< pdcontact >>
rect 35 64 39 68
rect 3 47 7 51
rect 3 40 7 44
rect 14 55 18 59
rect 24 55 28 59
rect 46 55 50 59
rect 56 56 60 60
rect 56 49 60 53
<< psubstratepcontact >>
rect 4 4 8 8
<< nsubstratencontact >>
rect 4 64 8 68
<< psubstratepdiff >>
rect 3 8 9 9
rect 3 4 4 8
rect 8 4 9 8
rect 3 3 9 4
<< nsubstratendiff >>
rect 3 68 9 69
rect 3 64 4 68
rect 8 64 9 68
rect 3 63 9 64
<< labels >>
rlabel polycontact 12 32 12 32 6 zn
rlabel metal1 12 16 12 16 6 z
rlabel metal1 4 36 4 36 6 z
rlabel metal1 28 32 28 32 6 a
rlabel metal1 28 40 28 40 6 b
rlabel metal1 14 36 14 36 6 zn
rlabel metal1 32 4 32 4 6 vss
rlabel metal1 36 24 36 24 6 a
rlabel metal1 44 24 44 24 6 a
rlabel metal1 44 32 44 32 6 d
rlabel metal1 36 48 36 48 6 b
rlabel metal1 44 48 44 48 6 c
rlabel metal1 32 68 32 68 6 vdd
rlabel metal1 36 15 36 15 6 zn
rlabel metal1 60 20 60 20 6 d
rlabel metal1 52 32 52 32 6 d
rlabel metal1 52 40 52 40 6 c
rlabel metal1 36 57 36 57 6 zn
<< end >>
