magic
tech scmos
timestamp 1179385079
<< checkpaint >>
rect -22 -25 78 105
<< ab >>
rect 0 0 56 80
<< pwell >>
rect -4 -7 60 36
<< nwell >>
rect -4 36 60 87
<< polysilicon >>
rect 9 70 11 74
rect 19 67 21 72
rect 29 67 31 72
rect 41 67 43 72
rect 9 39 11 42
rect 19 39 21 50
rect 29 47 31 50
rect 29 46 35 47
rect 29 42 30 46
rect 34 42 35 46
rect 29 41 35 42
rect 9 38 15 39
rect 9 34 10 38
rect 14 34 15 38
rect 9 33 15 34
rect 19 38 25 39
rect 19 34 20 38
rect 24 34 25 38
rect 19 33 25 34
rect 9 29 11 33
rect 22 29 24 33
rect 29 29 31 41
rect 41 39 43 50
rect 41 38 47 39
rect 41 35 42 38
rect 36 34 42 35
rect 46 34 47 38
rect 36 33 47 34
rect 36 29 38 33
rect 9 10 11 15
rect 22 7 24 12
rect 29 7 31 12
rect 36 7 38 12
<< ndiffusion >>
rect 4 23 9 29
rect 2 22 9 23
rect 2 18 3 22
rect 7 18 9 22
rect 2 17 9 18
rect 4 15 9 17
rect 11 15 22 29
rect 13 12 22 15
rect 24 12 29 29
rect 31 12 36 29
rect 38 22 43 29
rect 38 21 45 22
rect 38 17 40 21
rect 44 17 45 21
rect 38 16 45 17
rect 38 12 43 16
rect 13 8 15 12
rect 19 8 20 12
rect 13 7 20 8
<< pdiffusion >>
rect 33 72 39 73
rect 4 55 9 70
rect 2 54 9 55
rect 2 50 3 54
rect 7 50 9 54
rect 2 47 9 50
rect 2 43 3 47
rect 7 43 9 47
rect 2 42 9 43
rect 11 67 17 70
rect 33 68 34 72
rect 38 68 39 72
rect 33 67 39 68
rect 11 66 19 67
rect 11 62 13 66
rect 17 62 19 66
rect 11 50 19 62
rect 21 62 29 67
rect 21 58 23 62
rect 27 58 29 62
rect 21 55 29 58
rect 21 51 23 55
rect 27 51 29 55
rect 21 50 29 51
rect 31 50 41 67
rect 43 64 48 67
rect 43 63 50 64
rect 43 59 45 63
rect 49 59 50 63
rect 43 58 50 59
rect 43 50 48 58
rect 11 42 17 50
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect -2 72 58 78
rect -2 68 34 72
rect 38 68 58 72
rect 13 66 17 68
rect 13 61 17 62
rect 23 62 45 63
rect 27 59 45 62
rect 49 59 50 63
rect 27 58 28 59
rect 23 55 28 58
rect 2 54 7 55
rect 2 50 3 54
rect 2 47 7 50
rect 2 43 3 47
rect 2 42 7 43
rect 10 51 23 55
rect 27 51 28 55
rect 2 22 6 42
rect 10 38 14 51
rect 18 38 22 47
rect 42 46 46 55
rect 29 42 30 46
rect 34 42 46 46
rect 18 34 20 38
rect 24 34 31 38
rect 41 34 42 38
rect 46 34 47 38
rect 10 30 14 34
rect 41 30 47 34
rect 10 26 26 30
rect 33 26 47 30
rect 2 18 3 22
rect 7 18 15 22
rect 2 17 15 18
rect 22 21 26 26
rect 22 17 40 21
rect 44 17 45 21
rect -2 8 15 12
rect 19 8 58 12
rect -2 2 58 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
<< ntransistor >>
rect 9 15 11 29
rect 22 12 24 29
rect 29 12 31 29
rect 36 12 38 29
<< ptransistor >>
rect 9 42 11 70
rect 19 50 21 67
rect 29 50 31 67
rect 41 50 43 67
<< polycontact >>
rect 30 42 34 46
rect 10 34 14 38
rect 20 34 24 38
rect 42 34 46 38
<< ndcontact >>
rect 3 18 7 22
rect 40 17 44 21
rect 15 8 19 12
<< pdcontact >>
rect 3 50 7 54
rect 3 43 7 47
rect 34 68 38 72
rect 13 62 17 66
rect 23 58 27 62
rect 23 51 27 55
rect 45 59 49 63
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
<< psubstratepdiff >>
rect 0 2 56 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 56 2
rect 0 -3 56 -2
<< nsubstratendiff >>
rect 0 82 56 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 56 82
rect 0 77 56 78
<< labels >>
rlabel polycontact 12 36 12 36 6 zn
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 20 12 20 6 z
rlabel metal1 20 44 20 44 6 a
rlabel metal1 12 40 12 40 6 zn
rlabel metal1 28 6 28 6 6 vss
rlabel metal1 28 36 28 36 6 a
rlabel metal1 36 28 36 28 6 c
rlabel metal1 36 44 36 44 6 b
rlabel metal1 19 53 19 53 6 zn
rlabel metal1 25 57 25 57 6 zn
rlabel metal1 28 74 28 74 6 vdd
rlabel metal1 33 19 33 19 6 zn
rlabel metal1 44 32 44 32 6 c
rlabel metal1 44 52 44 52 6 b
rlabel metal1 36 61 36 61 6 zn
<< end >>
