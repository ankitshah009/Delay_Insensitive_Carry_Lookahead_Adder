magic
tech scmos
timestamp 1179385070
<< checkpaint >>
rect -22 -25 78 105
<< ab >>
rect 0 0 56 80
<< pwell >>
rect -4 -7 60 36
<< nwell >>
rect -4 36 60 87
<< polysilicon >>
rect 9 62 11 67
rect 19 62 21 67
rect 29 62 31 67
rect 41 61 43 66
rect 9 39 11 44
rect 19 39 21 49
rect 29 46 31 49
rect 29 45 35 46
rect 29 41 30 45
rect 34 41 35 45
rect 29 40 35 41
rect 9 38 15 39
rect 9 34 10 38
rect 14 34 15 38
rect 9 33 15 34
rect 19 38 25 39
rect 19 34 20 38
rect 24 34 25 38
rect 19 33 25 34
rect 9 29 11 33
rect 22 29 24 33
rect 29 29 31 40
rect 41 39 43 48
rect 41 38 47 39
rect 41 35 42 38
rect 36 34 42 35
rect 46 34 47 38
rect 36 33 47 34
rect 36 29 38 33
rect 9 15 11 20
rect 22 11 24 16
rect 29 11 31 16
rect 36 11 38 16
<< ndiffusion >>
rect 2 28 9 29
rect 2 24 3 28
rect 7 24 9 28
rect 2 23 9 24
rect 4 20 9 23
rect 11 20 22 29
rect 13 16 22 20
rect 24 16 29 29
rect 31 16 36 29
rect 38 22 43 29
rect 38 21 45 22
rect 38 17 40 21
rect 44 17 45 21
rect 38 16 45 17
rect 13 12 20 16
rect 13 8 14 12
rect 18 8 20 12
rect 13 7 20 8
<< pdiffusion >>
rect 33 72 39 73
rect 33 68 34 72
rect 38 68 39 72
rect 33 62 39 68
rect 4 57 9 62
rect 2 56 9 57
rect 2 52 3 56
rect 7 52 9 56
rect 2 49 9 52
rect 2 45 3 49
rect 7 45 9 49
rect 2 44 9 45
rect 11 61 19 62
rect 11 57 13 61
rect 17 57 19 61
rect 11 49 19 57
rect 21 61 29 62
rect 21 57 23 61
rect 27 57 29 61
rect 21 54 29 57
rect 21 50 23 54
rect 27 50 29 54
rect 21 49 29 50
rect 31 61 39 62
rect 31 49 41 61
rect 11 44 17 49
rect 36 48 41 49
rect 43 60 50 61
rect 43 56 45 60
rect 49 56 50 60
rect 43 53 50 56
rect 43 49 45 53
rect 49 49 50 53
rect 43 48 50 49
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect -2 72 58 78
rect -2 68 34 72
rect 38 68 58 72
rect 2 56 7 63
rect 12 61 18 68
rect 12 57 13 61
rect 17 57 18 61
rect 23 61 50 62
rect 27 60 50 61
rect 27 58 45 60
rect 2 52 3 56
rect 23 54 27 57
rect 44 56 45 58
rect 49 56 50 60
rect 7 52 15 54
rect 2 50 15 52
rect 18 50 23 53
rect 2 49 7 50
rect 2 45 3 49
rect 18 49 27 50
rect 18 46 22 49
rect 33 46 39 54
rect 44 53 50 56
rect 44 49 45 53
rect 49 49 50 53
rect 2 44 7 45
rect 2 29 6 44
rect 10 42 22 46
rect 25 45 47 46
rect 25 42 30 45
rect 10 38 14 42
rect 29 41 30 42
rect 34 42 47 45
rect 34 41 35 42
rect 17 34 20 38
rect 24 34 30 38
rect 10 29 14 34
rect 2 28 7 29
rect 2 24 3 28
rect 10 25 19 29
rect 26 25 30 34
rect 41 34 42 38
rect 46 34 47 38
rect 41 31 47 34
rect 34 25 47 31
rect 2 23 7 24
rect 2 17 6 23
rect 15 21 19 25
rect 15 17 40 21
rect 44 17 45 21
rect -2 8 14 12
rect 18 8 58 12
rect -2 2 58 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
<< ntransistor >>
rect 9 20 11 29
rect 22 16 24 29
rect 29 16 31 29
rect 36 16 38 29
<< ptransistor >>
rect 9 44 11 62
rect 19 49 21 62
rect 29 49 31 62
rect 41 48 43 61
<< polycontact >>
rect 30 41 34 45
rect 10 34 14 38
rect 20 34 24 38
rect 42 34 46 38
<< ndcontact >>
rect 3 24 7 28
rect 40 17 44 21
rect 14 8 18 12
<< pdcontact >>
rect 34 68 38 72
rect 3 52 7 56
rect 3 45 7 49
rect 13 57 17 61
rect 23 57 27 61
rect 23 50 27 54
rect 45 56 49 60
rect 45 49 49 53
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
<< psubstratepdiff >>
rect 0 2 56 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 56 2
rect 0 -3 56 -2
<< nsubstratendiff >>
rect 0 82 56 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 56 82
rect 0 77 56 78
<< labels >>
rlabel polycontact 12 36 12 36 6 zn
rlabel metal1 4 40 4 40 6 z
rlabel polycontact 12 35 12 35 6 zn
rlabel metal1 12 52 12 52 6 z
rlabel metal1 28 6 28 6 6 vss
rlabel metal1 28 28 28 28 6 a
rlabel metal1 20 36 20 36 6 a
rlabel metal1 28 44 28 44 6 b
rlabel metal1 25 55 25 55 6 zn
rlabel metal1 28 74 28 74 6 vdd
rlabel metal1 36 28 36 28 6 c
rlabel metal1 30 19 30 19 6 zn
rlabel metal1 44 32 44 32 6 c
rlabel metal1 44 44 44 44 6 b
rlabel polycontact 44 36 44 36 6 c
rlabel metal1 36 48 36 48 6 b
rlabel metal1 47 55 47 55 6 zn
<< end >>
