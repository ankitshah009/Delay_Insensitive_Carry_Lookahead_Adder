magic
tech scmos
timestamp 1179385424
<< checkpaint >>
rect -22 -25 94 105
<< ab >>
rect 0 0 72 80
<< pwell >>
rect -4 -7 76 36
<< nwell >>
rect -4 36 76 87
<< polysilicon >>
rect 9 67 11 72
rect 19 67 21 72
rect 29 67 31 72
rect 39 67 41 72
rect 49 67 51 72
rect 59 67 61 72
rect 9 39 11 50
rect 19 47 21 50
rect 29 47 31 50
rect 19 46 31 47
rect 19 45 26 46
rect 25 42 26 45
rect 30 42 31 46
rect 9 38 15 39
rect 9 34 10 38
rect 14 34 15 38
rect 25 38 31 42
rect 39 39 41 50
rect 49 39 51 42
rect 25 35 26 38
rect 9 33 15 34
rect 19 34 26 35
rect 30 34 31 38
rect 19 33 31 34
rect 35 38 41 39
rect 35 34 36 38
rect 40 34 41 38
rect 35 33 41 34
rect 45 38 51 39
rect 45 34 46 38
rect 50 34 51 38
rect 59 35 61 42
rect 45 33 51 34
rect 55 34 70 35
rect 55 33 65 34
rect 12 30 14 33
rect 19 30 21 33
rect 29 30 31 33
rect 36 30 38 33
rect 48 30 50 33
rect 55 30 57 33
rect 64 30 65 33
rect 69 30 70 34
rect 12 15 14 19
rect 19 15 21 19
rect 29 8 31 13
rect 36 8 38 13
rect 64 29 70 30
rect 48 6 50 10
rect 55 6 57 10
<< ndiffusion >>
rect 3 19 12 30
rect 14 19 19 30
rect 21 24 29 30
rect 21 20 23 24
rect 27 20 29 24
rect 21 19 29 20
rect 3 12 10 19
rect 24 13 29 19
rect 31 13 36 30
rect 38 15 48 30
rect 38 13 41 15
rect 3 8 5 12
rect 9 8 10 12
rect 40 11 41 13
rect 45 11 48 15
rect 40 10 48 11
rect 50 10 55 30
rect 57 23 62 30
rect 57 22 64 23
rect 57 18 59 22
rect 63 18 64 22
rect 57 17 64 18
rect 57 10 62 17
rect 3 7 10 8
<< pdiffusion >>
rect 2 66 9 67
rect 2 62 3 66
rect 7 62 9 66
rect 2 50 9 62
rect 11 62 19 67
rect 11 58 13 62
rect 17 58 19 62
rect 11 55 19 58
rect 11 51 13 55
rect 17 51 19 55
rect 11 50 19 51
rect 21 66 29 67
rect 21 62 23 66
rect 27 62 29 66
rect 21 50 29 62
rect 31 62 39 67
rect 31 58 33 62
rect 37 58 39 62
rect 31 55 39 58
rect 31 51 33 55
rect 37 51 39 55
rect 31 50 39 51
rect 41 66 49 67
rect 41 62 43 66
rect 47 62 49 66
rect 41 50 49 62
rect 43 42 49 50
rect 51 62 59 67
rect 51 58 53 62
rect 57 58 59 62
rect 51 55 59 58
rect 51 51 53 55
rect 57 51 59 55
rect 51 42 59 51
rect 61 66 69 67
rect 61 62 63 66
rect 67 62 69 66
rect 61 58 69 62
rect 61 54 63 58
rect 67 54 69 58
rect 61 42 69 54
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect -2 68 74 78
rect 3 66 7 68
rect 23 66 27 68
rect 3 61 7 62
rect 13 62 17 63
rect 43 66 47 68
rect 23 61 27 62
rect 33 62 38 63
rect 13 55 17 58
rect 2 51 13 55
rect 37 58 38 62
rect 63 66 67 68
rect 43 61 47 62
rect 53 62 57 63
rect 33 55 38 58
rect 17 51 33 54
rect 37 51 38 55
rect 53 55 57 58
rect 2 50 38 51
rect 42 51 53 54
rect 63 58 67 62
rect 63 53 67 54
rect 42 50 57 51
rect 2 22 6 50
rect 42 46 46 50
rect 17 42 26 46
rect 30 42 31 46
rect 10 38 14 39
rect 25 38 31 42
rect 25 34 26 38
rect 30 34 31 38
rect 36 42 46 46
rect 36 38 40 42
rect 50 41 62 47
rect 45 34 46 38
rect 10 31 14 34
rect 36 31 40 34
rect 10 27 40 31
rect 22 22 23 24
rect 2 20 23 22
rect 27 20 28 24
rect 2 18 28 20
rect 36 22 40 27
rect 50 25 54 41
rect 66 35 70 39
rect 65 34 70 35
rect 58 30 65 31
rect 69 30 70 34
rect 58 25 70 30
rect 36 18 59 22
rect 63 18 64 22
rect 40 12 41 15
rect -2 8 5 12
rect 9 11 41 12
rect 45 12 46 15
rect 45 11 74 12
rect 9 8 74 11
rect -2 2 74 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
<< ntransistor >>
rect 12 19 14 30
rect 19 19 21 30
rect 29 13 31 30
rect 36 13 38 30
rect 48 10 50 30
rect 55 10 57 30
<< ptransistor >>
rect 9 50 11 67
rect 19 50 21 67
rect 29 50 31 67
rect 39 50 41 67
rect 49 42 51 67
rect 59 42 61 67
<< polycontact >>
rect 26 42 30 46
rect 10 34 14 38
rect 26 34 30 38
rect 36 34 40 38
rect 46 34 50 38
rect 65 30 69 34
<< ndcontact >>
rect 23 20 27 24
rect 5 8 9 12
rect 41 11 45 15
rect 59 18 63 22
<< pdcontact >>
rect 3 62 7 66
rect 13 58 17 62
rect 13 51 17 55
rect 23 62 27 66
rect 33 58 37 62
rect 33 51 37 55
rect 43 62 47 66
rect 53 58 57 62
rect 53 51 57 55
rect 63 62 67 66
rect 63 54 67 58
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
<< psubstratepdiff >>
rect 0 2 72 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 72 2
rect 0 -3 72 -2
<< nsubstratendiff >>
rect 0 82 72 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 72 82
rect 0 77 72 78
<< labels >>
rlabel ntransistor 13 27 13 27 6 an
rlabel polycontact 38 36 38 36 6 an
rlabel metal1 4 40 4 40 6 z
rlabel metal1 12 20 12 20 6 z
rlabel metal1 20 20 20 20 6 z
rlabel metal1 12 33 12 33 6 an
rlabel metal1 20 44 20 44 6 b
rlabel metal1 20 52 20 52 6 z
rlabel metal1 12 52 12 52 6 z
rlabel metal1 36 6 36 6 6 vss
rlabel metal1 38 32 38 32 6 an
rlabel metal1 28 40 28 40 6 b
rlabel metal1 28 52 28 52 6 z
rlabel pdcontact 36 60 36 60 6 z
rlabel metal1 36 74 36 74 6 vdd
rlabel metal1 52 36 52 36 6 a1
rlabel metal1 55 56 55 56 6 an
rlabel metal1 60 28 60 28 6 a2
rlabel metal1 50 20 50 20 6 an
rlabel polycontact 68 32 68 32 6 a2
rlabel metal1 60 44 60 44 6 a1
<< end >>
