magic
tech scmos
timestamp 1185039059
<< checkpaint >>
rect -22 -24 152 124
<< ab >>
rect 0 0 130 100
<< pwell >>
rect -2 -4 132 49
<< nwell >>
rect -2 49 132 104
<< polysilicon >>
rect 11 95 13 98
rect 23 95 25 98
rect 35 95 37 98
rect 47 95 49 98
rect 69 95 71 98
rect 81 95 83 98
rect 93 95 95 98
rect 105 95 107 98
rect 117 75 119 78
rect 11 53 13 55
rect 23 53 25 55
rect 35 53 37 55
rect 47 53 49 55
rect 69 53 71 55
rect 81 53 83 55
rect 11 51 19 53
rect 23 51 29 53
rect 35 52 43 53
rect 35 51 38 52
rect 17 43 19 51
rect 27 43 29 51
rect 37 48 38 51
rect 42 48 43 52
rect 37 47 43 48
rect 47 52 53 53
rect 47 48 48 52
rect 52 48 53 52
rect 47 47 53 48
rect 67 52 73 53
rect 67 48 68 52
rect 72 48 73 52
rect 67 47 73 48
rect 77 52 83 53
rect 77 48 78 52
rect 82 48 83 52
rect 77 47 83 48
rect 17 42 23 43
rect 17 38 18 42
rect 22 38 23 42
rect 17 37 23 38
rect 27 42 33 43
rect 27 38 28 42
rect 32 38 33 42
rect 27 37 33 38
rect 17 29 19 37
rect 27 29 29 37
rect 37 29 39 47
rect 47 29 49 47
rect 15 27 19 29
rect 23 27 29 29
rect 35 27 39 29
rect 43 27 49 29
rect 69 29 71 47
rect 69 27 75 29
rect 15 25 17 27
rect 23 25 25 27
rect 35 25 37 27
rect 43 25 45 27
rect 73 25 75 27
rect 81 25 83 47
rect 93 41 95 55
rect 105 43 107 55
rect 105 42 113 43
rect 105 41 108 42
rect 93 39 108 41
rect 93 25 95 39
rect 105 38 108 39
rect 112 38 113 42
rect 105 37 113 38
rect 105 25 107 37
rect 117 33 119 55
rect 111 32 119 33
rect 111 28 112 32
rect 116 28 119 32
rect 111 27 119 28
rect 117 25 119 27
rect 117 12 119 15
rect 15 2 17 5
rect 23 2 25 5
rect 35 2 37 5
rect 43 2 45 5
rect 73 2 75 5
rect 81 2 83 5
rect 93 2 95 5
rect 105 2 107 5
<< ndiffusion >>
rect 97 32 103 33
rect 97 28 98 32
rect 102 28 103 32
rect 97 25 103 28
rect 7 12 15 25
rect 7 8 8 12
rect 12 8 15 12
rect 7 5 15 8
rect 17 5 23 25
rect 25 22 35 25
rect 25 18 28 22
rect 32 18 35 22
rect 25 5 35 18
rect 37 5 43 25
rect 45 12 53 25
rect 45 8 48 12
rect 52 8 53 12
rect 45 5 53 8
rect 65 22 73 25
rect 65 18 66 22
rect 70 18 73 22
rect 65 5 73 18
rect 75 5 81 25
rect 83 12 93 25
rect 83 8 86 12
rect 90 8 93 12
rect 83 5 93 8
rect 95 5 105 25
rect 107 15 117 25
rect 119 22 127 25
rect 119 18 122 22
rect 126 18 127 22
rect 119 15 127 18
rect 107 12 115 15
rect 107 8 110 12
rect 114 8 115 12
rect 107 5 115 8
<< pdiffusion >>
rect 3 82 11 95
rect 3 78 4 82
rect 8 78 11 82
rect 3 55 11 78
rect 13 72 23 95
rect 13 68 16 72
rect 20 68 23 72
rect 13 55 23 68
rect 25 82 35 95
rect 25 78 28 82
rect 32 78 35 82
rect 25 55 35 78
rect 37 72 47 95
rect 37 68 40 72
rect 44 68 47 72
rect 37 55 47 68
rect 49 83 53 95
rect 61 94 69 95
rect 61 90 62 94
rect 66 90 69 94
rect 61 89 69 90
rect 49 82 57 83
rect 49 78 52 82
rect 56 78 57 82
rect 49 55 57 78
rect 63 55 69 89
rect 71 82 81 95
rect 71 78 74 82
rect 78 78 81 82
rect 71 55 81 78
rect 83 92 93 95
rect 83 88 86 92
rect 90 88 93 92
rect 83 82 93 88
rect 83 78 86 82
rect 90 78 93 82
rect 83 72 93 78
rect 83 68 86 72
rect 90 68 93 72
rect 83 55 93 68
rect 95 82 105 95
rect 95 78 98 82
rect 102 78 105 82
rect 95 72 105 78
rect 95 68 98 72
rect 102 68 105 72
rect 95 62 105 68
rect 95 58 98 62
rect 102 58 105 62
rect 95 55 105 58
rect 107 92 115 95
rect 107 88 110 92
rect 114 88 115 92
rect 107 82 115 88
rect 107 78 110 82
rect 114 78 115 82
rect 107 75 115 78
rect 107 72 117 75
rect 107 68 110 72
rect 114 68 117 72
rect 107 55 117 68
rect 119 72 127 75
rect 119 68 122 72
rect 126 68 127 72
rect 119 62 127 68
rect 119 58 122 62
rect 126 58 127 62
rect 119 55 127 58
<< metal1 >>
rect -2 94 132 101
rect -2 90 62 94
rect 66 92 122 94
rect 66 90 86 92
rect -2 88 86 90
rect 90 88 110 92
rect 114 90 122 92
rect 126 90 132 94
rect 114 88 132 90
rect -2 87 132 88
rect 3 82 9 83
rect 27 82 33 83
rect 51 82 57 83
rect 3 78 4 82
rect 8 78 28 82
rect 32 78 52 82
rect 56 78 57 82
rect 3 77 9 78
rect 27 77 33 78
rect 51 77 57 78
rect 73 82 79 83
rect 73 78 74 82
rect 78 78 79 82
rect 73 77 79 78
rect 85 82 91 87
rect 85 78 86 82
rect 90 78 91 82
rect 15 72 21 73
rect 39 72 45 73
rect 74 72 78 77
rect 15 71 16 72
rect 8 68 16 71
rect 20 68 21 72
rect 8 67 21 68
rect 8 22 12 67
rect 17 42 23 62
rect 17 38 18 42
rect 22 38 23 42
rect 17 28 23 38
rect 27 42 33 72
rect 39 68 40 72
rect 44 68 78 72
rect 85 72 91 78
rect 85 68 86 72
rect 90 68 91 72
rect 39 67 45 68
rect 85 67 91 68
rect 97 82 103 83
rect 97 78 98 82
rect 102 78 103 82
rect 97 72 103 78
rect 97 68 98 72
rect 102 68 103 72
rect 97 62 103 68
rect 109 82 115 87
rect 109 78 110 82
rect 114 78 115 82
rect 109 72 115 78
rect 109 68 110 72
rect 114 68 115 72
rect 109 67 115 68
rect 121 72 127 73
rect 121 68 122 72
rect 126 68 127 72
rect 121 67 127 68
rect 122 63 126 67
rect 27 38 28 42
rect 32 38 33 42
rect 27 28 33 38
rect 37 52 43 62
rect 37 48 38 52
rect 42 48 43 52
rect 37 28 43 48
rect 47 52 53 62
rect 47 48 48 52
rect 52 48 53 52
rect 47 28 53 48
rect 67 52 73 62
rect 67 48 68 52
rect 72 48 73 52
rect 67 28 73 48
rect 77 52 83 62
rect 77 48 78 52
rect 82 48 83 52
rect 77 28 83 48
rect 97 58 98 62
rect 102 58 103 62
rect 97 32 103 58
rect 121 62 127 63
rect 121 58 122 62
rect 126 58 127 62
rect 121 57 127 58
rect 107 42 113 43
rect 122 42 126 57
rect 107 38 108 42
rect 112 38 126 42
rect 107 37 113 38
rect 97 28 98 32
rect 102 28 103 32
rect 97 27 103 28
rect 111 32 117 33
rect 111 28 112 32
rect 116 28 117 32
rect 111 27 117 28
rect 27 22 33 23
rect 65 22 71 23
rect 112 22 116 27
rect 122 23 126 38
rect 8 18 28 22
rect 32 18 66 22
rect 70 18 116 22
rect 121 22 127 23
rect 121 18 122 22
rect 126 18 127 22
rect 27 17 33 18
rect 65 17 71 18
rect 121 17 127 18
rect -2 12 132 13
rect -2 8 8 12
rect 12 8 48 12
rect 52 8 86 12
rect 90 8 110 12
rect 114 8 132 12
rect -2 -1 132 8
<< ntransistor >>
rect 15 5 17 25
rect 23 5 25 25
rect 35 5 37 25
rect 43 5 45 25
rect 73 5 75 25
rect 81 5 83 25
rect 93 5 95 25
rect 105 5 107 25
rect 117 15 119 25
<< ptransistor >>
rect 11 55 13 95
rect 23 55 25 95
rect 35 55 37 95
rect 47 55 49 95
rect 69 55 71 95
rect 81 55 83 95
rect 93 55 95 95
rect 105 55 107 95
rect 117 55 119 75
<< polycontact >>
rect 38 48 42 52
rect 48 48 52 52
rect 68 48 72 52
rect 78 48 82 52
rect 18 38 22 42
rect 28 38 32 42
rect 108 38 112 42
rect 112 28 116 32
<< ndcontact >>
rect 98 28 102 32
rect 8 8 12 12
rect 28 18 32 22
rect 48 8 52 12
rect 66 18 70 22
rect 86 8 90 12
rect 122 18 126 22
rect 110 8 114 12
<< pdcontact >>
rect 4 78 8 82
rect 16 68 20 72
rect 28 78 32 82
rect 40 68 44 72
rect 62 90 66 94
rect 52 78 56 82
rect 74 78 78 82
rect 86 88 90 92
rect 86 78 90 82
rect 86 68 90 72
rect 98 78 102 82
rect 98 68 102 72
rect 98 58 102 62
rect 110 88 114 92
rect 110 78 114 82
rect 110 68 114 72
rect 122 68 126 72
rect 122 58 126 62
<< nsubstratencontact >>
rect 122 90 126 94
<< nsubstratendiff >>
rect 121 94 127 95
rect 121 90 122 94
rect 126 90 127 94
rect 121 83 127 90
<< labels >>
rlabel metal1 20 45 20 45 6 i5
rlabel metal1 20 45 20 45 6 i5
rlabel metal1 40 45 40 45 6 i3
rlabel metal1 30 50 30 50 6 i4
rlabel metal1 30 50 30 50 6 i4
rlabel metal1 40 45 40 45 6 i3
rlabel metal1 65 6 65 6 6 vss
rlabel metal1 65 6 65 6 6 vss
rlabel metal1 50 45 50 45 6 i2
rlabel metal1 50 45 50 45 6 i2
rlabel metal1 70 45 70 45 6 i1
rlabel metal1 70 45 70 45 6 i1
rlabel metal1 65 94 65 94 6 vdd
rlabel metal1 65 94 65 94 6 vdd
rlabel metal1 80 45 80 45 6 i0
rlabel metal1 80 45 80 45 6 i0
rlabel metal1 100 55 100 55 6 nq
rlabel metal1 100 55 100 55 6 nq
<< end >>
