.subckt iv1v7x4 a vdd vss z
*   SPICE3 file   created from iv1v7x4.ext -      technology: scmos
m00 z      a      vdd    vdd p w=28u  l=2.3636u ad=176p     pd=50u      as=196p     ps=70u
m01 vdd    a      z      vdd p w=28u  l=2.3636u ad=196p     pd=70u      as=176p     ps=50u
m02 z      a      vss    vss n w=20u  l=2.3636u ad=136p     pd=42u      as=140p     ps=54u
m03 vss    a      z      vss n w=20u  l=2.3636u ad=140p     pd=54u      as=136p     ps=42u
C0  vss    z      0.123f
C1  z      a      0.218f
C2  vss    vdd    0.007f
C3  a      vdd    0.071f
C4  vss    a      0.063f
C5  z      vdd    0.076f
C7  z      vss    0.003f
C8  a      vss    0.091f
.ends
