magic
tech scmos
timestamp 1179387254
<< checkpaint >>
rect -22 -22 78 94
<< ab >>
rect 0 0 56 72
<< pwell >>
rect -4 -4 60 32
<< nwell >>
rect -4 32 60 76
<< polysilicon >>
rect 9 66 11 70
rect 22 66 24 70
rect 29 66 31 70
rect 36 66 38 70
rect 9 35 11 38
rect 22 35 24 38
rect 9 34 15 35
rect 9 30 10 34
rect 14 30 15 34
rect 9 29 15 30
rect 19 34 25 35
rect 19 30 20 34
rect 24 30 25 34
rect 19 29 25 30
rect 9 25 11 29
rect 19 19 21 29
rect 29 28 31 38
rect 36 35 38 38
rect 36 34 49 35
rect 36 33 44 34
rect 41 30 44 33
rect 48 30 49 34
rect 41 29 49 30
rect 29 27 37 28
rect 29 23 32 27
rect 36 23 37 27
rect 29 22 37 23
rect 29 19 31 22
rect 41 19 43 29
rect 9 6 11 11
rect 19 6 21 11
rect 29 6 31 11
rect 41 6 43 11
<< ndiffusion >>
rect 2 24 9 25
rect 2 20 3 24
rect 7 20 9 24
rect 2 19 9 20
rect 4 11 9 19
rect 11 19 16 25
rect 11 16 19 19
rect 11 12 13 16
rect 17 12 19 16
rect 11 11 19 12
rect 21 18 29 19
rect 21 14 23 18
rect 27 14 29 18
rect 21 11 29 14
rect 31 11 41 19
rect 43 18 50 19
rect 43 14 45 18
rect 49 14 50 18
rect 43 13 50 14
rect 43 11 48 13
rect 33 8 39 11
rect 33 4 34 8
rect 38 4 39 8
rect 33 3 39 4
<< pdiffusion >>
rect 13 68 20 69
rect 13 66 14 68
rect 4 60 9 66
rect 2 59 9 60
rect 2 55 3 59
rect 7 55 9 59
rect 2 52 9 55
rect 2 48 3 52
rect 7 48 9 52
rect 2 47 9 48
rect 4 38 9 47
rect 11 64 14 66
rect 18 66 20 68
rect 18 64 22 66
rect 11 38 22 64
rect 24 38 29 66
rect 31 38 36 66
rect 38 59 43 66
rect 38 58 45 59
rect 38 54 40 58
rect 44 54 45 58
rect 38 53 45 54
rect 38 38 43 53
<< metal1 >>
rect -2 68 58 72
rect -2 64 14 68
rect 18 64 48 68
rect 52 64 58 68
rect 2 55 3 59
rect 7 55 14 59
rect 2 53 14 55
rect 18 54 40 58
rect 44 54 45 58
rect 2 52 7 53
rect 2 48 3 52
rect 2 47 7 48
rect 2 25 6 47
rect 18 43 22 54
rect 34 45 46 51
rect 10 39 22 43
rect 10 34 14 39
rect 26 34 30 43
rect 17 30 20 34
rect 24 30 30 34
rect 10 25 14 30
rect 34 27 38 35
rect 42 34 46 45
rect 42 30 44 34
rect 48 30 49 34
rect 2 24 7 25
rect 2 20 3 24
rect 10 21 26 25
rect 31 23 32 27
rect 36 26 38 27
rect 36 23 47 26
rect 31 22 47 23
rect 2 19 7 20
rect 2 13 6 19
rect 22 18 26 21
rect 13 16 17 17
rect 22 14 23 18
rect 27 14 45 18
rect 49 14 50 18
rect 13 8 17 12
rect -2 4 34 8
rect 38 4 58 8
rect -2 0 58 4
<< ntransistor >>
rect 9 11 11 25
rect 19 11 21 19
rect 29 11 31 19
rect 41 11 43 19
<< ptransistor >>
rect 9 38 11 66
rect 22 38 24 66
rect 29 38 31 66
rect 36 38 38 66
<< polycontact >>
rect 10 30 14 34
rect 20 30 24 34
rect 44 30 48 34
rect 32 23 36 27
<< ndcontact >>
rect 3 20 7 24
rect 13 12 17 16
rect 23 14 27 18
rect 45 14 49 18
rect 34 4 38 8
<< pdcontact >>
rect 3 55 7 59
rect 3 48 7 52
rect 14 64 18 68
rect 40 54 44 58
<< nsubstratencontact >>
rect 48 64 52 68
<< nsubstratendiff >>
rect 47 68 53 69
rect 47 64 48 68
rect 52 64 53 68
rect 47 63 53 64
<< labels >>
rlabel polycontact 12 32 12 32 6 zn
rlabel metal1 4 36 4 36 6 z
rlabel metal1 20 32 20 32 6 a
rlabel polycontact 12 32 12 32 6 zn
rlabel metal1 12 56 12 56 6 z
rlabel metal1 28 4 28 4 6 vss
rlabel metal1 36 28 36 28 6 b
rlabel metal1 28 40 28 40 6 a
rlabel metal1 36 48 36 48 6 c
rlabel metal1 28 68 28 68 6 vdd
rlabel metal1 36 16 36 16 6 zn
rlabel metal1 44 24 44 24 6 b
rlabel metal1 44 44 44 44 6 c
rlabel metal1 31 56 31 56 6 zn
<< end >>
