.subckt oai23av0x05 a3 b1 b2 vdd vss z
*   SPICE3 file   created from oai23av0x05.ext -      technology: scmos
m00 w1     b      vdd    vdd p w=16u  l=2.3636u ad=40p      pd=21u      as=137.931p ps=47.4483u
m01 z      a3     w1     vdd p w=16u  l=2.3636u ad=64p      pd=24u      as=40p      ps=21u
m02 w2     b2     z      vdd p w=16u  l=2.3636u ad=40p      pd=21u      as=64p      ps=24u
m03 vdd    b1     w2     vdd p w=16u  l=2.3636u ad=137.931p pd=47.4483u as=40p      ps=21u
m04 b      b1     vdd    vdd p w=13u  l=2.3636u ad=52p      pd=21u      as=112.069p ps=38.5517u
m05 vdd    b2     b      vdd p w=13u  l=2.3636u ad=112.069p pd=38.5517u as=52p      ps=21u
m06 n4     a3     vss    vss n w=7u   l=2.3636u ad=28p      pd=15u      as=72.52p   ps=28.56u
m07 z      b2     n4     vss n w=7u   l=2.3636u ad=28p      pd=15u      as=28p      ps=15u
m08 n4     b1     z      vss n w=7u   l=2.3636u ad=28p      pd=15u      as=28p      ps=15u
m09 vss    b      n4     vss n w=7u   l=2.3636u ad=72.52p   pd=28.56u   as=28p      ps=15u
m10 w3     b1     vss    vss n w=11u  l=2.3636u ad=27.5p    pd=16u      as=113.96p  ps=44.88u
m11 b      b2     w3     vss n w=11u  l=2.3636u ad=67p      pd=36u      as=27.5p    ps=16u
C0  n4     z      0.145f
C1  b2     b      0.437f
C2  b1     vdd    0.026f
C3  n4     b1     0.003f
C4  a3     vdd    0.016f
C5  z      w1     0.003f
C6  w3     b      0.006f
C7  vss    b2     0.035f
C8  n4     a3     0.060f
C9  z      b2     0.134f
C10 n4     vdd    0.006f
C11 vss    b      0.137f
C12 b1     b2     0.395f
C13 z      b      0.261f
C14 b1     b      0.347f
C15 b2     a3     0.081f
C16 vss    z      0.031f
C17 a3     b      0.123f
C18 b2     vdd    0.096f
C19 n4     b2     0.026f
C20 vss    b1     0.026f
C21 b      vdd    0.553f
C22 w2     b2     0.004f
C23 vss    a3     0.068f
C24 z      b1     0.016f
C25 n4     b      0.048f
C26 vss    vdd    0.003f
C27 z      a3     0.076f
C28 w2     b      0.010f
C29 n4     vss    0.178f
C30 z      vdd    0.038f
C31 b1     a3     0.049f
C32 w1     b      0.015f
C33 n4     vss    0.011f
C35 z      vss    0.012f
C36 b1     vss    0.045f
C37 b2     vss    0.051f
C38 a3     vss    0.027f
C39 b      vss    0.044f
.ends
