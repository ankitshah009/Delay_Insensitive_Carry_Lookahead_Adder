magic
tech scmos
timestamp 1179387537
<< checkpaint >>
rect -22 -25 94 105
<< ab >>
rect 0 0 72 80
<< pwell >>
rect -4 -7 76 36
<< nwell >>
rect -4 36 76 87
<< polysilicon >>
rect 9 54 11 59
rect 41 72 63 74
rect 21 62 27 63
rect 21 58 22 62
rect 26 58 27 62
rect 21 57 27 58
rect 31 62 37 63
rect 31 58 32 62
rect 36 58 37 62
rect 31 57 37 58
rect 21 54 23 57
rect 31 54 33 57
rect 41 54 43 72
rect 61 63 63 72
rect 51 54 53 59
rect 9 38 11 42
rect 9 37 15 38
rect 9 33 10 37
rect 14 33 15 37
rect 21 35 23 42
rect 31 39 33 42
rect 31 37 37 39
rect 41 38 43 42
rect 51 39 53 42
rect 61 39 63 51
rect 48 38 54 39
rect 9 32 15 33
rect 19 32 23 35
rect 35 34 37 37
rect 48 34 49 38
rect 53 34 54 38
rect 9 29 11 32
rect 19 29 21 32
rect 29 29 31 33
rect 35 32 41 34
rect 48 33 54 34
rect 58 38 64 39
rect 58 34 59 38
rect 63 34 64 38
rect 58 33 64 34
rect 39 29 41 32
rect 50 30 52 33
rect 9 18 11 23
rect 19 18 21 23
rect 29 8 31 23
rect 39 18 41 23
rect 50 19 52 24
rect 61 23 63 33
rect 61 8 63 17
rect 29 6 63 8
<< ndiffusion >>
rect 43 29 50 30
rect 2 28 9 29
rect 2 24 3 28
rect 7 24 9 28
rect 2 23 9 24
rect 11 23 19 29
rect 21 28 29 29
rect 21 24 23 28
rect 27 24 29 28
rect 21 23 29 24
rect 31 28 39 29
rect 31 24 33 28
rect 37 24 39 28
rect 31 23 39 24
rect 41 25 44 29
rect 48 25 50 29
rect 41 24 50 25
rect 52 24 59 30
rect 41 23 46 24
rect 13 13 17 23
rect 11 12 17 13
rect 11 8 12 12
rect 16 8 17 12
rect 11 7 17 8
rect 54 23 59 24
rect 54 17 61 23
rect 63 22 70 23
rect 63 18 65 22
rect 69 18 70 22
rect 63 17 70 18
rect 54 16 59 17
rect 53 15 59 16
rect 53 11 54 15
rect 58 11 59 15
rect 53 10 59 11
<< pdiffusion >>
rect 13 72 19 73
rect 13 68 14 72
rect 18 68 19 72
rect 13 54 19 68
rect 53 69 59 70
rect 53 65 54 69
rect 58 65 59 69
rect 53 63 59 65
rect 53 61 61 63
rect 55 54 61 61
rect 4 48 9 54
rect 2 47 9 48
rect 2 43 3 47
rect 7 43 9 47
rect 2 42 9 43
rect 11 42 21 54
rect 23 53 31 54
rect 23 49 25 53
rect 29 49 31 53
rect 23 42 31 49
rect 33 47 41 54
rect 33 43 35 47
rect 39 43 41 47
rect 33 42 41 43
rect 43 47 51 54
rect 43 43 45 47
rect 49 43 51 47
rect 43 42 51 43
rect 53 51 61 54
rect 63 62 70 63
rect 63 58 65 62
rect 69 58 70 62
rect 63 57 70 58
rect 63 51 68 57
rect 53 42 59 51
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect -2 72 74 78
rect -2 68 14 72
rect 18 69 74 72
rect 18 68 54 69
rect 53 65 54 68
rect 58 68 74 69
rect 58 65 59 68
rect 9 58 22 62
rect 26 58 27 62
rect 31 58 32 62
rect 36 58 65 62
rect 69 58 70 62
rect 18 49 22 58
rect 25 53 56 55
rect 29 51 56 53
rect 2 43 3 47
rect 7 43 14 47
rect 2 41 14 43
rect 2 29 6 41
rect 9 33 10 37
rect 14 33 16 37
rect 2 28 7 29
rect 2 24 3 28
rect 2 23 7 24
rect 12 21 16 33
rect 25 28 29 49
rect 22 24 23 28
rect 27 24 29 28
rect 33 47 39 48
rect 33 43 35 47
rect 33 42 39 43
rect 42 47 49 48
rect 42 43 45 47
rect 42 42 49 43
rect 33 28 37 42
rect 42 29 46 42
rect 52 39 56 51
rect 49 38 56 39
rect 53 34 56 38
rect 49 33 56 34
rect 59 38 63 39
rect 59 30 63 34
rect 42 25 44 29
rect 48 25 49 29
rect 57 26 63 30
rect 33 21 37 24
rect 57 22 61 26
rect 66 23 70 58
rect 12 17 37 21
rect 49 18 61 22
rect 65 22 70 23
rect 69 18 70 22
rect 65 17 70 18
rect 53 12 54 15
rect -2 8 12 12
rect 16 11 54 12
rect 58 12 59 15
rect 58 11 74 12
rect 16 8 74 11
rect -2 2 74 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
<< ntransistor >>
rect 9 23 11 29
rect 19 23 21 29
rect 29 23 31 29
rect 39 23 41 29
rect 50 24 52 30
rect 61 17 63 23
<< ptransistor >>
rect 9 42 11 54
rect 21 42 23 54
rect 31 42 33 54
rect 41 42 43 54
rect 51 42 53 54
rect 61 51 63 63
<< polycontact >>
rect 22 58 26 62
rect 32 58 36 62
rect 10 33 14 37
rect 49 34 53 38
rect 59 34 63 38
<< ndcontact >>
rect 3 24 7 28
rect 23 24 27 28
rect 33 24 37 28
rect 44 25 48 29
rect 12 8 16 12
rect 65 18 69 22
rect 54 11 58 15
<< pdcontact >>
rect 14 68 18 72
rect 54 65 58 69
rect 3 43 7 47
rect 25 49 29 53
rect 35 43 39 47
rect 45 43 49 47
rect 65 58 69 62
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
<< psubstratepdiff >>
rect 0 2 72 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 72 2
rect 0 -3 72 -2
<< nsubstratendiff >>
rect 0 82 72 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 72 82
rect 0 77 72 78
<< labels >>
rlabel polycontact 12 35 12 35 6 zn
rlabel polycontact 34 60 34 60 6 bn
rlabel polycontact 51 36 51 36 6 an
rlabel metal1 4 36 4 36 6 z
rlabel metal1 14 27 14 27 6 zn
rlabel metal1 12 44 12 44 6 z
rlabel metal1 12 60 12 60 6 a
rlabel metal1 20 56 20 56 6 a
rlabel metal1 36 6 36 6 6 vss
rlabel metal1 27 39 27 39 6 an
rlabel metal1 35 32 35 32 6 zn
rlabel metal1 36 74 36 74 6 vdd
rlabel metal1 52 20 52 20 6 b
rlabel metal1 44 36 44 36 6 ai
rlabel metal1 54 44 54 44 6 an
rlabel metal1 60 28 60 28 6 b
rlabel metal1 68 39 68 39 6 bn
rlabel metal1 50 60 50 60 6 bn
<< end >>
