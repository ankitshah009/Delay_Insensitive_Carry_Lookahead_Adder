magic
tech scmos
timestamp 1179386744
<< checkpaint >>
rect -22 -25 70 105
<< ab >>
rect 0 0 48 80
<< pwell >>
rect -4 -7 52 36
<< nwell >>
rect -4 36 52 87
<< polysilicon >>
rect 9 70 11 74
rect 16 70 18 74
rect 26 70 28 74
rect 33 70 35 74
rect 9 34 11 43
rect 16 40 18 43
rect 26 40 28 43
rect 16 38 28 40
rect 21 34 23 38
rect 27 34 28 38
rect 9 33 17 34
rect 9 31 12 33
rect 11 29 12 31
rect 16 29 17 33
rect 11 28 17 29
rect 21 33 28 34
rect 11 25 13 28
rect 21 25 23 33
rect 33 31 35 43
rect 33 30 39 31
rect 33 26 34 30
rect 38 26 39 30
rect 33 25 39 26
rect 11 6 13 10
rect 21 6 23 10
<< ndiffusion >>
rect 3 15 11 25
rect 3 11 5 15
rect 9 11 11 15
rect 3 10 11 11
rect 13 22 21 25
rect 13 18 15 22
rect 19 18 21 22
rect 13 10 21 18
rect 23 22 31 25
rect 23 18 25 22
rect 29 18 31 22
rect 23 15 31 18
rect 23 11 25 15
rect 29 11 31 15
rect 23 10 31 11
<< pdiffusion >>
rect 2 69 9 70
rect 2 65 3 69
rect 7 65 9 69
rect 2 62 9 65
rect 2 58 3 62
rect 7 58 9 62
rect 2 43 9 58
rect 11 43 16 70
rect 18 55 26 70
rect 18 51 20 55
rect 24 51 26 55
rect 18 48 26 51
rect 18 44 20 48
rect 24 44 26 48
rect 18 43 26 44
rect 28 43 33 70
rect 35 69 42 70
rect 35 65 37 69
rect 41 65 42 69
rect 35 62 42 65
rect 35 58 37 62
rect 41 58 42 62
rect 35 43 42 58
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect -2 69 50 78
rect -2 68 3 69
rect 2 65 3 68
rect 7 68 37 69
rect 7 65 8 68
rect 2 62 8 65
rect 2 58 3 62
rect 7 58 8 62
rect 36 65 37 68
rect 41 68 50 69
rect 41 65 42 68
rect 36 62 42 65
rect 36 58 37 62
rect 41 58 42 62
rect 18 55 24 56
rect 18 51 20 55
rect 18 48 24 51
rect 18 46 20 48
rect 2 44 20 46
rect 2 42 24 44
rect 2 22 6 42
rect 34 38 39 47
rect 22 34 23 38
rect 27 34 39 38
rect 12 33 16 34
rect 16 29 34 30
rect 12 26 34 29
rect 38 26 39 30
rect 2 18 15 22
rect 19 18 20 22
rect 24 18 25 22
rect 29 18 30 22
rect 24 15 30 18
rect 34 17 39 26
rect 4 12 5 15
rect -2 11 5 12
rect 9 12 10 15
rect 24 12 25 15
rect 9 11 25 12
rect 29 12 30 15
rect 29 11 50 12
rect -2 2 50 11
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
<< ntransistor >>
rect 11 10 13 25
rect 21 10 23 25
<< ptransistor >>
rect 9 43 11 70
rect 16 43 18 70
rect 26 43 28 70
rect 33 43 35 70
<< polycontact >>
rect 23 34 27 38
rect 12 29 16 33
rect 34 26 38 30
<< ndcontact >>
rect 5 11 9 15
rect 15 18 19 22
rect 25 18 29 22
rect 25 11 29 15
<< pdcontact >>
rect 3 65 7 69
rect 3 58 7 62
rect 20 51 24 55
rect 20 44 24 48
rect 37 65 41 69
rect 37 58 41 62
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
<< psubstratepdiff >>
rect 0 2 48 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 48 2
rect 0 -3 48 -2
<< nsubstratendiff >>
rect 0 82 48 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 48 82
rect 0 77 48 78
<< labels >>
rlabel metal1 4 32 4 32 6 z
rlabel metal1 12 20 12 20 6 z
rlabel metal1 20 28 20 28 6 a
rlabel metal1 12 44 12 44 6 z
rlabel metal1 20 48 20 48 6 z
rlabel metal1 24 6 24 6 6 vss
rlabel metal1 28 28 28 28 6 a
rlabel metal1 28 36 28 36 6 b
rlabel metal1 24 74 24 74 6 vdd
rlabel metal1 36 24 36 24 6 a
rlabel metal1 36 40 36 40 6 b
<< end >>
