magic
tech scmos
timestamp 1180600703
<< checkpaint >>
rect -22 -22 142 122
<< ab >>
rect 0 0 120 100
<< pwell >>
rect -4 -4 124 48
<< nwell >>
rect -4 48 124 104
<< polysilicon >>
rect 11 85 13 89
rect 93 94 95 98
rect 105 94 107 98
rect 23 85 25 89
rect 31 85 33 89
rect 47 85 49 89
rect 55 85 57 89
rect 67 85 69 89
rect 11 41 13 65
rect 23 63 25 66
rect 17 62 25 63
rect 17 58 18 62
rect 22 61 25 62
rect 22 58 23 61
rect 17 57 23 58
rect 31 43 33 66
rect 47 57 49 66
rect 55 63 57 66
rect 55 62 63 63
rect 55 61 58 62
rect 57 58 58 61
rect 62 58 63 62
rect 57 57 63 58
rect 47 56 53 57
rect 47 52 48 56
rect 52 52 53 56
rect 47 51 53 52
rect 37 50 43 51
rect 37 46 38 50
rect 42 47 43 50
rect 67 47 69 65
rect 73 52 79 53
rect 73 48 74 52
rect 78 51 79 52
rect 93 51 95 55
rect 105 51 107 55
rect 78 49 107 51
rect 78 48 79 49
rect 73 47 79 48
rect 42 46 69 47
rect 37 45 69 46
rect 27 42 33 43
rect 27 41 28 42
rect 11 39 28 41
rect 11 15 13 39
rect 27 38 28 39
rect 32 41 33 42
rect 32 39 49 41
rect 32 38 33 39
rect 27 37 33 38
rect 17 32 23 33
rect 17 28 18 32
rect 22 29 23 32
rect 22 28 25 29
rect 17 27 25 28
rect 23 14 25 27
rect 29 22 35 23
rect 29 18 30 22
rect 34 18 35 22
rect 29 17 35 18
rect 31 14 33 17
rect 47 15 49 39
rect 57 32 63 33
rect 57 29 58 32
rect 55 28 58 29
rect 62 28 63 32
rect 55 27 63 28
rect 55 15 57 27
rect 67 15 69 45
rect 93 25 95 49
rect 105 25 107 49
rect 11 2 13 6
rect 23 2 25 6
rect 31 2 33 6
rect 47 2 49 6
rect 55 2 57 6
rect 67 2 69 6
rect 93 2 95 6
rect 105 2 107 6
<< ndiffusion >>
rect 3 22 9 23
rect 3 18 4 22
rect 8 18 9 22
rect 3 15 9 18
rect 37 32 45 33
rect 3 6 11 15
rect 13 14 18 15
rect 37 28 38 32
rect 42 28 45 32
rect 37 15 45 28
rect 71 22 77 23
rect 71 18 72 22
rect 76 18 77 22
rect 71 15 77 18
rect 37 14 47 15
rect 13 12 23 14
rect 13 8 16 12
rect 20 8 23 12
rect 13 6 23 8
rect 25 6 31 14
rect 33 6 47 14
rect 49 6 55 15
rect 57 12 67 15
rect 57 8 60 12
rect 64 8 67 12
rect 57 6 67 8
rect 69 6 77 15
rect 85 22 93 25
rect 85 18 86 22
rect 90 18 93 22
rect 85 12 93 18
rect 85 8 86 12
rect 90 8 93 12
rect 85 6 93 8
rect 95 22 105 25
rect 95 18 98 22
rect 102 18 105 22
rect 95 6 105 18
rect 107 22 115 25
rect 107 18 110 22
rect 114 18 115 22
rect 107 12 115 18
rect 107 8 110 12
rect 114 8 115 12
rect 107 6 115 8
<< pdiffusion >>
rect 15 92 21 93
rect 15 88 16 92
rect 20 88 21 92
rect 59 92 65 93
rect 15 85 21 88
rect 59 88 60 92
rect 64 88 65 92
rect 85 92 93 94
rect 59 85 65 88
rect 85 88 86 92
rect 90 88 93 92
rect 3 82 11 85
rect 3 78 4 82
rect 8 78 11 82
rect 3 72 11 78
rect 3 68 4 72
rect 8 68 11 72
rect 3 65 11 68
rect 13 66 23 85
rect 25 66 31 85
rect 33 82 47 85
rect 33 78 38 82
rect 42 78 47 82
rect 33 72 47 78
rect 33 68 38 72
rect 42 68 47 72
rect 33 66 47 68
rect 49 66 55 85
rect 57 66 67 85
rect 13 65 18 66
rect 62 65 67 66
rect 69 82 77 85
rect 69 78 72 82
rect 76 78 77 82
rect 69 70 77 78
rect 69 66 72 70
rect 76 66 77 70
rect 69 65 77 66
rect 85 82 93 88
rect 85 78 86 82
rect 90 78 93 82
rect 85 72 93 78
rect 85 68 86 72
rect 90 68 93 72
rect 85 62 93 68
rect 85 58 86 62
rect 90 58 93 62
rect 85 55 93 58
rect 95 82 105 94
rect 95 78 98 82
rect 102 78 105 82
rect 95 72 105 78
rect 95 68 98 72
rect 102 68 105 72
rect 95 62 105 68
rect 95 58 98 62
rect 102 58 105 62
rect 95 55 105 58
rect 107 92 115 94
rect 107 88 110 92
rect 114 88 115 92
rect 107 82 115 88
rect 107 78 110 82
rect 114 78 115 82
rect 107 72 115 78
rect 107 68 110 72
rect 114 68 115 72
rect 107 62 115 68
rect 107 58 110 62
rect 114 58 115 62
rect 107 55 115 58
<< metal1 >>
rect -2 96 122 100
rect -2 92 28 96
rect 32 92 38 96
rect 42 92 48 96
rect 52 92 122 96
rect -2 88 16 92
rect 20 88 60 92
rect 64 88 86 92
rect 90 88 110 92
rect 114 88 122 92
rect 4 82 8 83
rect 4 72 8 78
rect 4 22 8 68
rect 18 62 22 83
rect 18 32 22 58
rect 18 27 22 28
rect 28 42 32 83
rect 28 27 32 38
rect 38 82 42 83
rect 38 72 42 78
rect 38 50 42 68
rect 58 62 62 83
rect 38 32 42 46
rect 38 27 42 28
rect 48 56 52 57
rect 48 22 52 52
rect 8 18 30 22
rect 34 18 52 22
rect 58 32 62 58
rect 4 17 8 18
rect 58 17 62 28
rect 72 82 76 83
rect 72 70 76 78
rect 72 52 76 66
rect 86 82 90 88
rect 86 72 90 78
rect 86 62 90 68
rect 86 57 90 58
rect 98 82 102 83
rect 98 72 102 78
rect 98 62 102 68
rect 72 48 74 52
rect 78 48 79 52
rect 72 22 76 48
rect 72 17 76 18
rect 86 22 90 23
rect 86 12 90 18
rect 98 22 102 58
rect 110 82 114 88
rect 110 72 114 78
rect 110 62 114 68
rect 110 57 114 58
rect 98 17 102 18
rect 110 22 114 23
rect 110 12 114 18
rect -2 8 16 12
rect 20 8 60 12
rect 64 8 86 12
rect 90 8 110 12
rect 114 8 122 12
rect -2 0 122 8
<< ntransistor >>
rect 11 6 13 15
rect 23 6 25 14
rect 31 6 33 14
rect 47 6 49 15
rect 55 6 57 15
rect 67 6 69 15
rect 93 6 95 25
rect 105 6 107 25
<< ptransistor >>
rect 11 65 13 85
rect 23 66 25 85
rect 31 66 33 85
rect 47 66 49 85
rect 55 66 57 85
rect 67 65 69 85
rect 93 55 95 94
rect 105 55 107 94
<< polycontact >>
rect 18 58 22 62
rect 58 58 62 62
rect 48 52 52 56
rect 38 46 42 50
rect 74 48 78 52
rect 28 38 32 42
rect 18 28 22 32
rect 30 18 34 22
rect 58 28 62 32
<< ndcontact >>
rect 4 18 8 22
rect 38 28 42 32
rect 72 18 76 22
rect 16 8 20 12
rect 60 8 64 12
rect 86 18 90 22
rect 86 8 90 12
rect 98 18 102 22
rect 110 18 114 22
rect 110 8 114 12
<< pdcontact >>
rect 16 88 20 92
rect 60 88 64 92
rect 86 88 90 92
rect 4 78 8 82
rect 4 68 8 72
rect 38 78 42 82
rect 38 68 42 72
rect 72 78 76 82
rect 72 66 76 70
rect 86 78 90 82
rect 86 68 90 72
rect 86 58 90 62
rect 98 78 102 82
rect 98 68 102 72
rect 98 58 102 62
rect 110 88 114 92
rect 110 78 114 82
rect 110 68 114 72
rect 110 58 114 62
<< nsubstratencontact >>
rect 28 92 32 96
rect 38 92 42 96
rect 48 92 52 96
<< nsubstratendiff >>
rect 27 96 53 97
rect 27 92 28 96
rect 32 92 38 96
rect 42 92 48 96
rect 52 92 53 96
rect 27 91 53 92
<< labels >>
rlabel metal1 20 55 20 55 6 i0
rlabel metal1 30 55 30 55 6 cmd
rlabel metal1 60 6 60 6 6 vss
rlabel metal1 60 50 60 50 6 i1
rlabel metal1 60 94 60 94 6 vdd
rlabel metal1 100 50 100 50 6 nq
<< end >>
