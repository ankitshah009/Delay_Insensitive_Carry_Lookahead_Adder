magic
tech scmos
timestamp 1179387654
<< checkpaint >>
rect -22 -25 158 105
<< ab >>
rect 0 0 136 80
<< pwell >>
rect -4 -7 140 36
<< nwell >>
rect -4 36 140 87
<< polysilicon >>
rect 20 70 22 74
rect 30 70 32 74
rect 45 70 47 74
rect 55 70 57 74
rect 85 70 87 74
rect 95 70 97 74
rect 105 70 107 74
rect 115 70 117 74
rect 125 70 127 74
rect 71 63 77 64
rect 65 55 67 60
rect 71 59 72 63
rect 76 59 77 63
rect 71 58 77 59
rect 75 55 77 58
rect 20 39 22 42
rect 30 39 32 42
rect 45 39 47 42
rect 55 39 57 42
rect 9 38 51 39
rect 9 34 10 38
rect 14 37 51 38
rect 14 34 21 37
rect 9 33 21 34
rect 9 30 11 33
rect 19 30 21 33
rect 39 30 41 37
rect 49 30 51 37
rect 55 38 61 39
rect 55 34 56 38
rect 60 34 61 38
rect 65 37 67 42
rect 75 37 77 42
rect 85 39 87 42
rect 95 39 97 42
rect 105 39 107 42
rect 85 38 97 39
rect 65 35 80 37
rect 55 33 61 34
rect 59 30 61 33
rect 66 30 68 35
rect 78 30 80 35
rect 85 34 86 38
rect 90 37 97 38
rect 101 38 107 39
rect 90 34 91 37
rect 85 33 91 34
rect 101 34 102 38
rect 106 34 107 38
rect 101 33 107 34
rect 115 39 117 42
rect 125 39 127 42
rect 115 38 127 39
rect 115 34 122 38
rect 126 34 127 38
rect 115 33 127 34
rect 85 30 87 33
rect 115 30 117 33
rect 125 30 127 33
rect 9 15 11 19
rect 19 8 21 13
rect 39 11 41 16
rect 49 11 51 16
rect 59 6 61 11
rect 66 6 68 11
rect 115 12 117 16
rect 125 12 127 16
rect 78 6 80 11
rect 85 6 87 11
<< ndiffusion >>
rect 2 24 9 30
rect 2 20 3 24
rect 7 20 9 24
rect 2 19 9 20
rect 11 29 19 30
rect 11 25 13 29
rect 17 25 19 29
rect 11 19 19 25
rect 14 13 19 19
rect 21 18 28 30
rect 21 14 23 18
rect 27 14 28 18
rect 32 29 39 30
rect 32 25 33 29
rect 37 25 39 29
rect 32 22 39 25
rect 32 18 33 22
rect 37 18 39 22
rect 32 16 39 18
rect 41 29 49 30
rect 41 25 43 29
rect 47 25 49 29
rect 41 16 49 25
rect 51 29 59 30
rect 51 25 53 29
rect 57 25 59 29
rect 51 22 59 25
rect 51 18 53 22
rect 57 18 59 22
rect 51 16 59 18
rect 21 13 28 14
rect 54 11 59 16
rect 61 11 66 30
rect 68 12 78 30
rect 68 11 71 12
rect 70 8 71 11
rect 75 11 78 12
rect 80 11 85 30
rect 87 23 92 30
rect 87 22 94 23
rect 87 18 89 22
rect 93 18 94 22
rect 87 17 94 18
rect 108 21 115 30
rect 108 17 109 21
rect 113 17 115 21
rect 87 11 92 17
rect 108 16 115 17
rect 117 29 125 30
rect 117 25 119 29
rect 123 25 125 29
rect 117 22 125 25
rect 117 18 119 22
rect 123 18 125 22
rect 117 16 125 18
rect 127 21 134 30
rect 127 17 129 21
rect 133 17 134 21
rect 127 16 134 17
rect 75 8 76 11
rect 70 7 76 8
<< pdiffusion >>
rect 13 69 20 70
rect 13 65 14 69
rect 18 65 20 69
rect 13 62 20 65
rect 13 58 14 62
rect 18 58 20 62
rect 13 42 20 58
rect 22 54 30 70
rect 22 50 24 54
rect 28 50 30 54
rect 22 47 30 50
rect 22 43 24 47
rect 28 43 30 47
rect 22 42 30 43
rect 32 69 45 70
rect 32 65 36 69
rect 40 65 45 69
rect 32 62 45 65
rect 32 58 36 62
rect 40 58 45 62
rect 32 42 45 58
rect 47 62 55 70
rect 47 58 49 62
rect 53 58 55 62
rect 47 55 55 58
rect 47 51 49 55
rect 53 51 55 55
rect 47 42 55 51
rect 57 55 62 70
rect 80 55 85 70
rect 57 54 65 55
rect 57 50 59 54
rect 63 50 65 54
rect 57 47 65 50
rect 57 43 59 47
rect 63 43 65 47
rect 57 42 65 43
rect 67 47 75 55
rect 67 43 69 47
rect 73 43 75 47
rect 67 42 75 43
rect 77 54 85 55
rect 77 50 79 54
rect 83 50 85 54
rect 77 42 85 50
rect 87 63 95 70
rect 87 59 89 63
rect 93 59 95 63
rect 87 47 95 59
rect 87 43 89 47
rect 93 43 95 47
rect 87 42 95 43
rect 97 62 105 70
rect 97 58 99 62
rect 103 58 105 62
rect 97 55 105 58
rect 97 51 99 55
rect 103 51 105 55
rect 97 42 105 51
rect 107 54 115 70
rect 107 50 109 54
rect 113 50 115 54
rect 107 47 115 50
rect 107 43 109 47
rect 113 43 115 47
rect 107 42 115 43
rect 117 69 125 70
rect 117 65 119 69
rect 123 65 125 69
rect 117 62 125 65
rect 117 58 119 62
rect 123 58 125 62
rect 117 42 125 58
rect 127 55 132 70
rect 127 54 134 55
rect 127 50 129 54
rect 133 50 134 54
rect 127 47 134 50
rect 127 43 129 47
rect 133 43 134 47
rect 127 42 134 43
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect 118 78 122 82
rect 126 78 130 82
rect 134 78 138 82
rect -2 69 138 78
rect -2 68 14 69
rect 18 68 36 69
rect 14 62 18 65
rect 35 65 36 68
rect 40 68 119 69
rect 40 65 41 68
rect 35 62 41 65
rect 123 68 138 69
rect 35 58 36 62
rect 40 58 41 62
rect 49 62 72 63
rect 53 59 72 62
rect 76 59 89 63
rect 93 59 94 63
rect 98 62 103 63
rect 14 57 18 58
rect 49 55 53 58
rect 23 50 24 54
rect 28 51 49 54
rect 98 58 99 62
rect 98 55 103 58
rect 119 62 123 65
rect 119 57 123 58
rect 98 54 99 55
rect 28 50 53 51
rect 58 50 59 54
rect 63 50 79 54
rect 83 51 99 54
rect 83 50 103 51
rect 108 54 113 55
rect 108 50 109 54
rect 23 47 28 50
rect 2 39 6 47
rect 23 43 24 47
rect 58 47 63 50
rect 108 47 113 50
rect 129 54 134 55
rect 133 50 134 54
rect 129 47 134 50
rect 58 46 59 47
rect 23 42 28 43
rect 34 43 59 46
rect 34 42 63 43
rect 68 43 69 47
rect 73 43 74 47
rect 2 38 14 39
rect 2 34 10 38
rect 2 33 14 34
rect 23 29 27 42
rect 34 29 38 42
rect 68 38 74 43
rect 88 43 89 47
rect 93 46 94 47
rect 93 43 103 46
rect 108 43 109 47
rect 113 43 129 47
rect 133 43 134 47
rect 88 42 103 43
rect 99 38 103 42
rect 12 25 13 29
rect 17 25 27 29
rect 32 25 33 29
rect 37 25 38 29
rect 42 34 56 38
rect 60 34 86 38
rect 90 34 93 38
rect 99 34 102 38
rect 106 34 107 38
rect 42 29 48 34
rect 89 30 93 34
rect 112 30 116 43
rect 121 38 134 39
rect 121 34 122 38
rect 126 34 134 38
rect 42 25 43 29
rect 47 25 48 29
rect 53 29 57 30
rect 89 29 123 30
rect 89 26 119 29
rect 3 24 7 25
rect 3 12 7 20
rect 32 22 38 25
rect 53 22 57 25
rect 130 25 134 34
rect 119 22 123 25
rect 23 18 27 19
rect 32 18 33 22
rect 37 18 53 22
rect 57 18 89 22
rect 93 18 95 22
rect 109 21 113 22
rect 23 12 27 14
rect 119 17 123 18
rect 128 17 129 21
rect 133 17 134 21
rect 109 12 113 17
rect 128 12 134 17
rect -2 8 71 12
rect 75 8 138 12
rect -2 2 138 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 122 2
rect 126 -2 130 2
rect 134 -2 138 2
<< ntransistor >>
rect 9 19 11 30
rect 19 13 21 30
rect 39 16 41 30
rect 49 16 51 30
rect 59 11 61 30
rect 66 11 68 30
rect 78 11 80 30
rect 85 11 87 30
rect 115 16 117 30
rect 125 16 127 30
<< ptransistor >>
rect 20 42 22 70
rect 30 42 32 70
rect 45 42 47 70
rect 55 42 57 70
rect 65 42 67 55
rect 75 42 77 55
rect 85 42 87 70
rect 95 42 97 70
rect 105 42 107 70
rect 115 42 117 70
rect 125 42 127 70
<< polycontact >>
rect 72 59 76 63
rect 10 34 14 38
rect 56 34 60 38
rect 86 34 90 38
rect 102 34 106 38
rect 122 34 126 38
<< ndcontact >>
rect 3 20 7 24
rect 13 25 17 29
rect 23 14 27 18
rect 33 25 37 29
rect 33 18 37 22
rect 43 25 47 29
rect 53 25 57 29
rect 53 18 57 22
rect 71 8 75 12
rect 89 18 93 22
rect 109 17 113 21
rect 119 25 123 29
rect 119 18 123 22
rect 129 17 133 21
<< pdcontact >>
rect 14 65 18 69
rect 14 58 18 62
rect 24 50 28 54
rect 24 43 28 47
rect 36 65 40 69
rect 36 58 40 62
rect 49 58 53 62
rect 49 51 53 55
rect 59 50 63 54
rect 59 43 63 47
rect 69 43 73 47
rect 79 50 83 54
rect 89 59 93 63
rect 89 43 93 47
rect 99 58 103 62
rect 99 51 103 55
rect 109 50 113 54
rect 109 43 113 47
rect 119 65 123 69
rect 119 58 123 62
rect 129 50 133 54
rect 129 43 133 47
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
rect 90 -2 94 2
rect 98 -2 102 2
rect 106 -2 110 2
rect 114 -2 118 2
rect 122 -2 126 2
rect 130 -2 134 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
rect 90 78 94 82
rect 98 78 102 82
rect 106 78 110 82
rect 114 78 118 82
rect 122 78 126 82
rect 130 78 134 82
<< psubstratepdiff >>
rect 0 2 136 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 122 2
rect 126 -2 130 2
rect 134 -2 136 2
rect 0 -3 136 -2
<< nsubstratendiff >>
rect 0 82 136 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect 118 78 122 82
rect 126 78 130 82
rect 134 78 136 82
rect 0 77 136 78
<< labels >>
rlabel polycontact 88 36 88 36 6 an
rlabel polycontact 74 61 74 61 6 bn
rlabel polycontact 104 36 104 36 6 bn
rlabel metal1 4 40 4 40 6 b
rlabel polycontact 12 36 12 36 6 b
rlabel metal1 19 27 19 27 6 bn
rlabel ndcontact 36 28 36 28 6 z
rlabel metal1 44 20 44 20 6 z
rlabel metal1 45 31 45 31 6 an
rlabel metal1 44 44 44 44 6 z
rlabel metal1 51 56 51 56 6 bn
rlabel metal1 38 52 38 52 6 bn
rlabel metal1 25 48 25 48 6 bn
rlabel metal1 68 6 68 6 6 vss
rlabel metal1 52 20 52 20 6 z
rlabel metal1 76 20 76 20 6 z
rlabel metal1 68 20 68 20 6 z
rlabel metal1 60 20 60 20 6 z
rlabel metal1 52 44 52 44 6 z
rlabel metal1 71 40 71 40 6 an
rlabel pdcontact 60 44 60 44 6 z
rlabel metal1 76 52 76 52 6 z
rlabel metal1 68 52 68 52 6 z
rlabel metal1 68 74 68 74 6 vdd
rlabel metal1 84 20 84 20 6 z
rlabel ndcontact 92 20 92 20 6 z
rlabel metal1 67 36 67 36 6 an
rlabel metal1 95 44 95 44 6 bn
rlabel polycontact 103 36 103 36 6 bn
rlabel metal1 92 52 92 52 6 z
rlabel metal1 84 52 84 52 6 z
rlabel metal1 71 61 71 61 6 bn
rlabel metal1 100 56 100 56 6 z
rlabel metal1 121 23 121 23 6 an
rlabel metal1 132 32 132 32 6 a
rlabel metal1 121 45 121 45 6 an
rlabel polycontact 124 36 124 36 6 a
rlabel metal1 131 49 131 49 6 an
rlabel metal1 110 49 110 49 6 an
<< end >>
