magic
tech scmos
timestamp 1185094763
<< checkpaint >>
rect -22 -22 72 122
<< ab >>
rect 0 0 50 100
<< pwell >>
rect -4 -4 54 48
<< nwell >>
rect -4 48 54 104
<< polysilicon >>
rect 15 94 17 98
rect 23 94 25 98
rect 37 77 39 82
rect 15 43 17 55
rect 23 52 25 55
rect 37 52 39 55
rect 23 49 27 52
rect 13 42 21 43
rect 13 38 16 42
rect 20 38 21 42
rect 13 37 21 38
rect 25 42 27 49
rect 32 51 39 52
rect 32 47 33 51
rect 37 47 39 51
rect 32 46 39 47
rect 25 41 32 42
rect 25 37 27 41
rect 31 37 32 41
rect 13 28 15 37
rect 25 36 32 37
rect 25 28 27 36
rect 37 28 39 46
rect 13 12 15 17
rect 25 12 27 17
rect 37 12 39 17
<< ndiffusion >>
rect 4 17 13 28
rect 15 22 25 28
rect 15 18 18 22
rect 22 18 25 22
rect 15 17 25 18
rect 27 22 37 28
rect 27 18 30 22
rect 34 18 37 22
rect 27 17 37 18
rect 39 27 47 28
rect 39 23 42 27
rect 46 23 47 27
rect 39 22 47 23
rect 39 17 44 22
rect 4 12 11 17
rect 4 8 6 12
rect 10 8 11 12
rect 4 7 11 8
<< pdiffusion >>
rect 10 69 15 94
rect 7 68 15 69
rect 7 64 8 68
rect 12 64 15 68
rect 7 60 15 64
rect 7 56 8 60
rect 12 56 15 60
rect 7 55 15 56
rect 17 55 23 94
rect 25 92 35 94
rect 25 88 28 92
rect 32 88 35 92
rect 25 82 35 88
rect 25 78 28 82
rect 32 78 35 82
rect 25 77 35 78
rect 25 72 37 77
rect 25 68 28 72
rect 32 68 37 72
rect 25 55 37 68
rect 39 69 44 77
rect 39 68 47 69
rect 39 64 42 68
rect 46 64 47 68
rect 39 60 47 64
rect 39 56 42 60
rect 46 56 47 60
rect 39 55 47 56
<< metal1 >>
rect -2 96 52 100
rect -2 92 42 96
rect 46 92 52 96
rect -2 88 28 92
rect 32 88 52 92
rect 28 82 32 88
rect 8 68 12 73
rect 8 60 12 64
rect 18 63 22 73
rect 28 72 32 78
rect 28 67 32 68
rect 42 68 46 69
rect 18 57 32 63
rect 8 23 12 56
rect 18 44 22 53
rect 28 51 32 57
rect 42 60 46 64
rect 28 47 33 51
rect 37 47 38 51
rect 16 42 22 44
rect 20 38 22 42
rect 42 41 46 56
rect 18 32 22 38
rect 26 37 27 41
rect 31 37 46 41
rect 18 27 33 32
rect 42 27 46 37
rect 8 22 22 23
rect 8 18 18 22
rect 8 17 22 18
rect 30 22 34 23
rect 42 22 46 23
rect 30 12 34 18
rect -2 8 6 12
rect 10 8 52 12
rect -2 4 18 8
rect 22 4 28 8
rect 32 4 52 8
rect -2 0 52 4
<< ntransistor >>
rect 13 17 15 28
rect 25 17 27 28
rect 37 17 39 28
<< ptransistor >>
rect 15 55 17 94
rect 23 55 25 94
rect 37 55 39 77
<< polycontact >>
rect 16 38 20 42
rect 33 47 37 51
rect 27 37 31 41
<< ndcontact >>
rect 18 18 22 22
rect 30 18 34 22
rect 42 23 46 27
rect 6 8 10 12
<< pdcontact >>
rect 8 64 12 68
rect 8 56 12 60
rect 28 88 32 92
rect 28 78 32 82
rect 28 68 32 72
rect 42 64 46 68
rect 42 56 46 60
<< psubstratepcontact >>
rect 18 4 22 8
rect 28 4 32 8
<< nsubstratencontact >>
rect 42 92 46 96
<< psubstratepdiff >>
rect 17 8 33 9
rect 17 4 18 8
rect 22 4 28 8
rect 32 4 33 8
rect 17 3 33 4
<< nsubstratendiff >>
rect 41 96 47 97
rect 41 92 42 96
rect 46 92 47 96
rect 41 91 47 92
<< labels >>
rlabel polycontact 28 39 28 39 6 an
rlabel ndcontact 20 20 20 20 6 z
rlabel metal1 10 45 10 45 6 z
rlabel metal1 20 40 20 40 6 b
rlabel metal1 20 65 20 65 6 a
rlabel metal1 25 6 25 6 6 vss
rlabel metal1 30 30 30 30 6 b
rlabel metal1 30 55 30 55 6 a
rlabel metal1 25 94 25 94 6 vdd
rlabel metal1 36 39 36 39 6 an
rlabel metal1 44 45 44 45 6 an
<< end >>
