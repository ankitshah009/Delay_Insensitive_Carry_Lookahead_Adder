magic
tech scmos
timestamp 1179385689
<< checkpaint >>
rect -22 -25 94 105
<< ab >>
rect 0 0 72 80
<< pwell >>
rect -4 -7 76 36
<< nwell >>
rect -4 36 76 87
<< polysilicon >>
rect 26 69 48 71
rect 56 69 58 74
rect 9 58 11 63
rect 19 58 21 63
rect 26 58 28 69
rect 46 66 48 69
rect 36 58 38 63
rect 9 37 11 42
rect 19 37 21 42
rect 26 39 28 42
rect 36 39 38 42
rect 9 35 21 37
rect 9 32 11 35
rect 5 31 11 32
rect 5 27 6 31
rect 10 27 11 31
rect 19 30 21 35
rect 25 38 31 39
rect 25 34 26 38
rect 30 34 31 38
rect 25 33 31 34
rect 36 38 42 39
rect 36 34 37 38
rect 41 34 42 38
rect 36 33 42 34
rect 26 30 28 33
rect 36 30 38 33
rect 46 30 48 50
rect 56 47 58 50
rect 56 46 63 47
rect 56 42 58 46
rect 62 42 63 46
rect 56 41 63 42
rect 56 30 58 41
rect 5 26 11 27
rect 9 23 11 26
rect 19 18 21 23
rect 26 18 28 23
rect 36 18 38 23
rect 46 18 48 23
rect 9 11 11 16
rect 56 15 58 20
<< ndiffusion >>
rect 13 23 19 30
rect 21 23 26 30
rect 28 29 36 30
rect 28 25 30 29
rect 34 25 36 29
rect 28 23 36 25
rect 38 28 46 30
rect 38 24 40 28
rect 44 24 46 28
rect 38 23 46 24
rect 48 28 56 30
rect 48 24 50 28
rect 54 24 56 28
rect 48 23 56 24
rect 2 21 9 23
rect 2 17 3 21
rect 7 17 9 21
rect 2 16 9 17
rect 11 16 17 23
rect 50 20 56 23
rect 58 29 65 30
rect 58 25 60 29
rect 64 25 65 29
rect 58 24 65 25
rect 58 20 63 24
rect 13 12 19 16
rect 13 8 14 12
rect 18 8 19 12
rect 13 7 19 8
<< pdiffusion >>
rect 13 72 19 73
rect 13 68 14 72
rect 18 68 19 72
rect 13 65 19 68
rect 13 58 17 65
rect 50 66 56 69
rect 41 58 46 66
rect 2 57 9 58
rect 2 53 3 57
rect 7 53 9 57
rect 2 50 9 53
rect 2 46 3 50
rect 7 46 9 50
rect 2 45 9 46
rect 4 42 9 45
rect 11 42 19 58
rect 21 42 26 58
rect 28 55 36 58
rect 28 51 30 55
rect 34 51 36 55
rect 28 42 36 51
rect 38 57 46 58
rect 38 53 40 57
rect 44 53 46 57
rect 38 50 46 53
rect 48 65 56 66
rect 48 61 50 65
rect 54 61 56 65
rect 48 50 56 61
rect 58 63 63 69
rect 58 62 65 63
rect 58 58 60 62
rect 64 58 65 62
rect 58 55 65 58
rect 58 51 60 55
rect 64 51 65 55
rect 58 50 65 51
rect 38 42 43 50
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect -2 72 74 78
rect -2 68 14 72
rect 18 68 74 72
rect 50 65 54 68
rect 3 59 44 63
rect 50 60 54 61
rect 60 62 64 63
rect 3 57 7 59
rect 40 57 44 59
rect 3 50 7 53
rect 10 51 30 55
rect 34 51 35 55
rect 60 55 64 58
rect 40 52 44 53
rect 50 51 60 54
rect 10 49 22 51
rect 3 45 7 46
rect 2 27 6 39
rect 10 27 14 31
rect 2 25 14 27
rect 18 29 22 49
rect 50 50 64 51
rect 26 41 38 47
rect 26 38 30 41
rect 50 38 54 50
rect 58 46 70 47
rect 62 42 70 46
rect 58 41 70 42
rect 36 34 37 38
rect 41 34 62 38
rect 26 33 30 34
rect 58 29 62 34
rect 66 33 70 41
rect 18 25 30 29
rect 34 25 35 29
rect 40 28 44 29
rect 40 21 44 24
rect 2 17 3 21
rect 7 17 44 21
rect 50 28 54 29
rect 58 25 60 29
rect 64 25 65 29
rect 50 12 54 24
rect -2 8 14 12
rect 18 8 74 12
rect -2 2 74 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
<< ntransistor >>
rect 19 23 21 30
rect 26 23 28 30
rect 36 23 38 30
rect 46 23 48 30
rect 9 16 11 23
rect 56 20 58 30
<< ptransistor >>
rect 9 42 11 58
rect 19 42 21 58
rect 26 42 28 58
rect 36 42 38 58
rect 46 50 48 66
rect 56 50 58 69
<< polycontact >>
rect 6 27 10 31
rect 26 34 30 38
rect 37 34 41 38
rect 58 42 62 46
<< ndcontact >>
rect 30 25 34 29
rect 40 24 44 28
rect 50 24 54 28
rect 3 17 7 21
rect 60 25 64 29
rect 14 8 18 12
<< pdcontact >>
rect 14 68 18 72
rect 3 53 7 57
rect 3 46 7 50
rect 30 51 34 55
rect 40 53 44 57
rect 50 61 54 65
rect 60 58 64 62
rect 60 51 64 55
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
<< psubstratepdiff >>
rect 0 2 72 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 72 2
rect 0 -3 72 -2
<< nsubstratendiff >>
rect 0 82 72 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 72 82
rect 0 77 72 78
<< labels >>
rlabel polycontact 39 36 39 36 6 cn
rlabel metal1 4 32 4 32 6 a
rlabel pdcontact 5 54 5 54 6 n1
rlabel metal1 12 28 12 28 6 a
rlabel metal1 20 40 20 40 6 z
rlabel metal1 12 52 12 52 6 z
rlabel metal1 36 6 36 6 6 vss
rlabel metal1 28 40 28 40 6 b
rlabel metal1 36 44 36 44 6 b
rlabel metal1 36 74 36 74 6 vdd
rlabel metal1 42 23 42 23 6 n3
rlabel metal1 23 19 23 19 6 n3
rlabel metal1 42 57 42 57 6 n1
rlabel metal1 60 31 60 31 6 cn
rlabel polycontact 60 44 60 44 6 c
rlabel metal1 49 36 49 36 6 cn
rlabel metal1 68 40 68 40 6 c
rlabel metal1 62 56 62 56 6 cn
<< end >>
