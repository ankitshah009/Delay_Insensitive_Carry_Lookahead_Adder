magic
tech scmos
timestamp 1179386436
<< checkpaint >>
rect -22 -25 134 105
<< ab >>
rect 0 0 112 80
<< pwell >>
rect -4 -7 116 36
<< nwell >>
rect -4 36 116 87
<< polysilicon >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 39 70 41 74
rect 49 70 51 74
rect 59 70 61 74
rect 69 70 71 74
rect 79 70 81 74
rect 90 60 92 65
rect 100 60 102 65
rect 9 39 11 43
rect 19 39 21 43
rect 29 39 31 43
rect 39 39 41 43
rect 49 39 51 43
rect 59 39 61 43
rect 69 39 71 43
rect 9 38 15 39
rect 9 34 10 38
rect 14 34 15 38
rect 9 33 15 34
rect 19 38 33 39
rect 19 34 26 38
rect 30 34 33 38
rect 19 33 33 34
rect 12 30 14 33
rect 19 30 21 33
rect 31 30 33 33
rect 38 38 51 39
rect 38 34 42 38
rect 46 34 51 38
rect 38 33 51 34
rect 55 38 71 39
rect 55 34 58 38
rect 62 37 71 38
rect 79 39 81 43
rect 90 39 92 43
rect 100 39 102 43
rect 79 38 92 39
rect 79 37 82 38
rect 62 34 63 37
rect 55 33 63 34
rect 81 34 82 37
rect 86 37 92 38
rect 96 38 102 39
rect 86 34 87 37
rect 81 33 87 34
rect 96 34 97 38
rect 101 34 102 38
rect 96 33 102 34
rect 38 30 40 33
rect 48 30 50 33
rect 55 30 57 33
rect 12 11 14 16
rect 19 11 21 16
rect 31 6 33 11
rect 38 6 40 11
rect 48 6 50 11
rect 55 6 57 11
<< ndiffusion >>
rect 5 29 12 30
rect 5 25 6 29
rect 10 25 12 29
rect 5 22 12 25
rect 5 18 6 22
rect 10 18 12 22
rect 5 16 12 18
rect 14 16 19 30
rect 21 16 31 30
rect 23 12 31 16
rect 23 8 24 12
rect 28 11 31 12
rect 33 11 38 30
rect 40 22 48 30
rect 40 18 42 22
rect 46 18 48 22
rect 40 11 48 18
rect 50 11 55 30
rect 57 12 66 30
rect 57 11 60 12
rect 28 8 29 11
rect 23 7 29 8
rect 59 8 60 11
rect 64 8 66 12
rect 59 7 66 8
<< pdiffusion >>
rect 2 69 9 70
rect 2 65 3 69
rect 7 65 9 69
rect 2 62 9 65
rect 2 58 3 62
rect 7 58 9 62
rect 2 43 9 58
rect 11 61 19 70
rect 11 57 13 61
rect 17 57 19 61
rect 11 54 19 57
rect 11 50 13 54
rect 17 50 19 54
rect 11 43 19 50
rect 21 69 29 70
rect 21 65 23 69
rect 27 65 29 69
rect 21 62 29 65
rect 21 58 23 62
rect 27 58 29 62
rect 21 43 29 58
rect 31 62 39 70
rect 31 58 33 62
rect 37 58 39 62
rect 31 54 39 58
rect 31 50 33 54
rect 37 50 39 54
rect 31 43 39 50
rect 41 69 49 70
rect 41 65 43 69
rect 47 65 49 69
rect 41 62 49 65
rect 41 58 43 62
rect 47 58 49 62
rect 41 43 49 58
rect 51 61 59 70
rect 51 57 53 61
rect 57 57 59 61
rect 51 54 59 57
rect 51 50 53 54
rect 57 50 59 54
rect 51 43 59 50
rect 61 69 69 70
rect 61 65 63 69
rect 67 65 69 69
rect 61 62 69 65
rect 61 58 63 62
rect 67 58 69 62
rect 61 43 69 58
rect 71 62 79 70
rect 71 58 73 62
rect 77 58 79 62
rect 71 54 79 58
rect 71 50 73 54
rect 77 50 79 54
rect 71 43 79 50
rect 81 69 88 70
rect 81 65 83 69
rect 87 65 88 69
rect 81 62 88 65
rect 81 58 83 62
rect 87 60 88 62
rect 87 58 90 60
rect 81 43 90 58
rect 92 54 100 60
rect 92 50 94 54
rect 98 50 100 54
rect 92 43 100 50
rect 102 59 110 60
rect 102 55 104 59
rect 108 55 110 59
rect 102 51 110 55
rect 102 47 104 51
rect 108 47 110 51
rect 102 43 110 47
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect -2 69 114 78
rect -2 68 3 69
rect 2 65 3 68
rect 7 68 23 69
rect 7 65 8 68
rect 2 62 8 65
rect 22 65 23 68
rect 27 68 43 69
rect 27 65 28 68
rect 22 62 28 65
rect 42 65 43 68
rect 47 68 63 69
rect 47 65 48 68
rect 2 58 3 62
rect 7 58 8 62
rect 13 61 17 62
rect 22 58 23 62
rect 27 58 28 62
rect 33 62 38 63
rect 37 58 38 62
rect 42 62 48 65
rect 62 65 63 68
rect 67 68 83 69
rect 67 65 68 68
rect 62 62 68 65
rect 82 65 83 68
rect 87 68 114 69
rect 87 65 88 68
rect 42 58 43 62
rect 47 58 48 62
rect 53 61 57 62
rect 13 54 17 57
rect 33 54 38 58
rect 62 58 63 62
rect 67 58 68 62
rect 73 62 78 63
rect 77 58 78 62
rect 82 62 88 65
rect 82 58 83 62
rect 87 58 88 62
rect 104 59 108 68
rect 53 54 57 57
rect 73 54 78 58
rect 2 50 13 54
rect 17 50 33 54
rect 37 50 53 54
rect 57 50 73 54
rect 77 50 94 54
rect 98 50 99 54
rect 104 51 108 55
rect 2 25 6 50
rect 104 46 108 47
rect 25 42 97 46
rect 10 38 20 39
rect 14 34 20 38
rect 25 38 31 42
rect 57 38 63 42
rect 25 34 26 38
rect 30 34 31 38
rect 41 34 42 38
rect 46 34 47 38
rect 57 34 58 38
rect 62 34 63 38
rect 81 34 82 38
rect 86 34 87 38
rect 93 34 97 42
rect 101 34 103 38
rect 10 33 20 34
rect 16 30 20 33
rect 41 30 47 34
rect 81 30 87 34
rect 10 25 11 29
rect 16 26 87 30
rect 5 22 11 25
rect 5 18 6 22
rect 10 18 42 22
rect 46 18 47 22
rect -2 8 24 12
rect 28 8 60 12
rect 64 8 114 12
rect -2 2 114 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
<< ntransistor >>
rect 12 16 14 30
rect 19 16 21 30
rect 31 11 33 30
rect 38 11 40 30
rect 48 11 50 30
rect 55 11 57 30
<< ptransistor >>
rect 9 43 11 70
rect 19 43 21 70
rect 29 43 31 70
rect 39 43 41 70
rect 49 43 51 70
rect 59 43 61 70
rect 69 43 71 70
rect 79 43 81 70
rect 90 43 92 60
rect 100 43 102 60
<< polycontact >>
rect 10 34 14 38
rect 26 34 30 38
rect 42 34 46 38
rect 58 34 62 38
rect 82 34 86 38
rect 97 34 101 38
<< ndcontact >>
rect 6 25 10 29
rect 6 18 10 22
rect 24 8 28 12
rect 42 18 46 22
rect 60 8 64 12
<< pdcontact >>
rect 3 65 7 69
rect 3 58 7 62
rect 13 57 17 61
rect 13 50 17 54
rect 23 65 27 69
rect 23 58 27 62
rect 33 58 37 62
rect 33 50 37 54
rect 43 65 47 69
rect 43 58 47 62
rect 53 57 57 61
rect 53 50 57 54
rect 63 65 67 69
rect 63 58 67 62
rect 73 58 77 62
rect 73 50 77 54
rect 83 65 87 69
rect 83 58 87 62
rect 94 50 98 54
rect 104 55 108 59
rect 104 47 108 51
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
rect 90 -2 94 2
rect 98 -2 102 2
rect 106 -2 110 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
rect 90 78 94 82
rect 98 78 102 82
rect 106 78 110 82
<< psubstratepdiff >>
rect 0 2 112 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 112 2
rect 0 -3 112 -2
<< nsubstratendiff >>
rect 0 82 112 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 112 82
rect 0 77 112 78
<< labels >>
rlabel metal1 12 20 12 20 6 z
rlabel polycontact 12 36 12 36 6 b
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 52 12 52 6 z
rlabel metal1 20 20 20 20 6 z
rlabel metal1 20 28 20 28 6 b
rlabel metal1 28 20 28 20 6 z
rlabel metal1 28 28 28 28 6 b
rlabel metal1 36 20 36 20 6 z
rlabel metal1 36 28 36 28 6 b
rlabel polycontact 28 36 28 36 6 a
rlabel metal1 28 40 28 40 6 a
rlabel metal1 36 44 36 44 6 a
rlabel metal1 28 52 28 52 6 z
rlabel metal1 20 52 20 52 6 z
rlabel metal1 36 56 36 56 6 z
rlabel metal1 56 6 56 6 6 vss
rlabel ndcontact 44 20 44 20 6 z
rlabel metal1 52 28 52 28 6 b
rlabel metal1 60 28 60 28 6 b
rlabel metal1 44 32 44 32 6 b
rlabel metal1 44 44 44 44 6 a
rlabel metal1 52 44 52 44 6 a
rlabel metal1 60 40 60 40 6 a
rlabel metal1 52 52 52 52 6 z
rlabel metal1 60 52 60 52 6 z
rlabel metal1 44 52 44 52 6 z
rlabel metal1 56 74 56 74 6 vdd
rlabel metal1 68 28 68 28 6 b
rlabel metal1 76 28 76 28 6 b
rlabel metal1 84 32 84 32 6 b
rlabel metal1 68 44 68 44 6 a
rlabel metal1 76 44 76 44 6 a
rlabel metal1 84 44 84 44 6 a
rlabel metal1 84 52 84 52 6 z
rlabel metal1 68 52 68 52 6 z
rlabel metal1 76 56 76 56 6 z
rlabel metal1 92 44 92 44 6 a
rlabel polycontact 100 36 100 36 6 a
rlabel metal1 92 52 92 52 6 z
<< end >>
