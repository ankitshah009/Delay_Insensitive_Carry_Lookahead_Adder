magic
tech scmos
timestamp 1179387145
<< checkpaint >>
rect -22 -25 86 105
<< ab >>
rect 0 0 64 80
<< pwell >>
rect -4 -7 68 36
<< nwell >>
rect -4 36 68 87
<< polysilicon >>
rect 39 69 41 74
rect 46 69 48 74
rect 29 62 31 67
rect 9 54 11 59
rect 29 47 31 54
rect 29 46 35 47
rect 29 42 30 46
rect 34 42 35 46
rect 9 39 11 42
rect 29 41 35 42
rect 9 38 18 39
rect 9 34 13 38
rect 17 34 18 38
rect 9 33 18 34
rect 9 30 11 33
rect 29 30 31 41
rect 39 39 41 54
rect 46 47 48 54
rect 46 46 57 47
rect 46 45 52 46
rect 51 42 52 45
rect 56 42 57 46
rect 51 41 57 42
rect 39 38 47 39
rect 39 34 42 38
rect 46 34 47 38
rect 39 33 47 34
rect 39 30 41 33
rect 9 19 11 24
rect 51 23 53 41
rect 29 18 31 23
rect 39 18 41 23
rect 51 11 53 16
<< ndiffusion >>
rect 2 29 9 30
rect 2 25 3 29
rect 7 25 9 29
rect 2 24 9 25
rect 11 29 18 30
rect 11 25 13 29
rect 17 25 18 29
rect 11 24 18 25
rect 22 29 29 30
rect 22 25 23 29
rect 27 25 29 29
rect 22 23 29 25
rect 31 28 39 30
rect 31 24 33 28
rect 37 24 39 28
rect 31 23 39 24
rect 41 23 49 30
rect 43 16 51 23
rect 53 21 60 23
rect 53 17 55 21
rect 59 17 60 21
rect 53 16 60 17
rect 43 12 49 16
rect 43 8 44 12
rect 48 8 49 12
rect 43 7 49 8
<< pdiffusion >>
rect 13 63 27 64
rect 13 59 14 63
rect 18 62 27 63
rect 34 62 39 69
rect 18 59 29 62
rect 13 55 29 59
rect 13 54 14 55
rect 4 48 9 54
rect 2 47 9 48
rect 2 43 3 47
rect 7 43 9 47
rect 2 42 9 43
rect 11 51 14 54
rect 18 54 29 55
rect 31 61 39 62
rect 31 57 33 61
rect 37 57 39 61
rect 31 54 39 57
rect 41 54 46 69
rect 48 68 56 69
rect 48 64 50 68
rect 54 64 56 68
rect 48 61 56 64
rect 48 57 50 61
rect 54 57 56 61
rect 48 54 56 57
rect 18 51 27 54
rect 11 42 27 51
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect -2 68 66 78
rect 13 63 19 68
rect 13 59 14 63
rect 18 59 19 63
rect 50 61 54 64
rect 13 55 19 59
rect 13 51 14 55
rect 18 51 19 55
rect 23 57 33 61
rect 37 57 38 61
rect 2 43 3 47
rect 7 43 15 47
rect 2 42 15 43
rect 2 30 6 42
rect 23 38 27 57
rect 50 56 54 57
rect 42 50 46 55
rect 34 47 46 50
rect 30 46 46 47
rect 50 46 62 47
rect 34 42 38 46
rect 30 41 38 42
rect 50 42 52 46
rect 56 42 62 46
rect 50 41 62 42
rect 12 34 13 38
rect 17 34 27 38
rect 2 29 7 30
rect 2 25 3 29
rect 2 24 7 25
rect 13 29 17 30
rect 2 17 6 24
rect 13 12 17 25
rect 23 29 27 34
rect 42 38 46 39
rect 42 31 46 34
rect 58 33 62 41
rect 23 24 27 25
rect 33 28 37 29
rect 42 25 54 31
rect 33 21 37 24
rect 33 17 55 21
rect 59 17 60 21
rect -2 8 44 12
rect 48 8 66 12
rect -2 2 66 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
<< ntransistor >>
rect 9 24 11 30
rect 29 23 31 30
rect 39 23 41 30
rect 51 16 53 23
<< ptransistor >>
rect 9 42 11 54
rect 29 54 31 62
rect 39 54 41 69
rect 46 54 48 69
<< polycontact >>
rect 30 42 34 46
rect 13 34 17 38
rect 52 42 56 46
rect 42 34 46 38
<< ndcontact >>
rect 3 25 7 29
rect 13 25 17 29
rect 23 25 27 29
rect 33 24 37 28
rect 55 17 59 21
rect 44 8 48 12
<< pdcontact >>
rect 14 59 18 63
rect 3 43 7 47
rect 14 51 18 55
rect 33 57 37 61
rect 50 64 54 68
rect 50 57 54 61
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
<< psubstratepdiff >>
rect 0 2 64 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 64 2
rect 0 -3 64 -2
<< nsubstratendiff >>
rect 0 82 64 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 64 82
rect 0 77 64 78
<< labels >>
rlabel polysilicon 13 36 13 36 6 zn
rlabel metal1 4 32 4 32 6 z
rlabel metal1 12 44 12 44 6 z
rlabel metal1 19 36 19 36 6 zn
rlabel metal1 25 42 25 42 6 zn
rlabel metal1 32 6 32 6 6 vss
rlabel metal1 35 23 35 23 6 n1
rlabel metal1 44 32 44 32 6 a2
rlabel metal1 36 44 36 44 6 b
rlabel metal1 30 59 30 59 6 zn
rlabel metal1 44 52 44 52 6 b
rlabel metal1 32 74 32 74 6 vdd
rlabel metal1 46 19 46 19 6 n1
rlabel metal1 52 28 52 28 6 a2
rlabel metal1 60 40 60 40 6 a1
rlabel metal1 52 44 52 44 6 a1
<< end >>
