.subckt nd2ab_x1 a b vdd vss z
*   SPICE3 file   created from nd2ab_x1.ext -      technology: scmos
m00 vdd    b      bn     vdd p w=18u  l=2.3636u ad=115.579p pd=36u      as=108p     ps=52u
m01 z      bn     vdd    vdd p w=20u  l=2.3636u ad=100p     pd=30u      as=128.421p ps=40u
m02 vdd    an     z      vdd p w=20u  l=2.3636u ad=128.421p pd=40u      as=100p     ps=30u
m03 an     a      vdd    vdd p w=18u  l=2.3636u ad=108p     pd=52u      as=115.579p ps=36u
m04 bn     b      vss    vss n w=9u   l=2.3636u ad=63p      pd=34u      as=72p      ps=27.2571u
m05 an     a      vss    vss n w=9u   l=2.3636u ad=63p      pd=34u      as=72p      ps=27.2571u
m06 w1     bn     z      vss n w=17u  l=2.3636u ad=51p      pd=23u      as=103p     ps=50u
m07 vss    an     w1     vss n w=17u  l=2.3636u ad=136p     pd=51.4857u as=51p      ps=23u
C0  vss    z      0.192f
C1  a      an     0.212f
C2  vss    bn     0.044f
C3  z      bn     0.138f
C4  a      b      0.041f
C5  an     b      0.024f
C6  z      vdd    0.008f
C7  w1     vss    0.010f
C8  bn     vdd    0.018f
C9  w1     z      0.010f
C10 vss    a      0.016f
C11 vss    an     0.079f
C12 a      z      0.131f
C13 z      an     0.070f
C14 a      bn     0.041f
C15 a      vdd    0.103f
C16 z      b      0.084f
C17 an     bn     0.121f
C18 an     vdd    0.008f
C19 bn     b      0.118f
C20 b      vdd    0.169f
C22 a      vss    0.024f
C23 z      vss    0.013f
C24 an     vss    0.039f
C25 bn     vss    0.037f
C26 b      vss    0.020f
.ends
