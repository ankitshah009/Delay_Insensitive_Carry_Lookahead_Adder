magic
tech scmos
timestamp 1179386772
<< checkpaint >>
rect -22 -25 150 105
<< ab >>
rect 0 0 128 80
<< pwell >>
rect -4 -7 132 36
<< nwell >>
rect -4 36 132 87
<< polysilicon >>
rect 9 70 11 74
rect 16 70 18 74
rect 26 70 28 74
rect 33 70 35 74
rect 43 70 45 74
rect 50 70 52 74
rect 60 70 62 74
rect 67 70 69 74
rect 77 70 79 74
rect 84 70 86 74
rect 94 70 96 74
rect 101 70 103 74
rect 9 33 11 42
rect 16 39 18 42
rect 26 39 28 42
rect 33 39 35 42
rect 43 39 45 42
rect 50 39 52 42
rect 60 39 62 42
rect 67 39 69 42
rect 77 39 79 42
rect 16 38 29 39
rect 16 37 24 38
rect 23 34 24 37
rect 28 34 29 38
rect 33 38 45 39
rect 33 37 38 38
rect 23 33 29 34
rect 37 34 38 37
rect 42 37 45 38
rect 49 38 63 39
rect 42 34 43 37
rect 37 33 43 34
rect 49 34 50 38
rect 54 37 63 38
rect 67 38 79 39
rect 67 37 74 38
rect 54 34 55 37
rect 49 33 55 34
rect 9 32 19 33
rect 9 31 14 32
rect 13 28 14 31
rect 18 28 19 32
rect 13 27 19 28
rect 17 24 19 27
rect 27 24 29 33
rect 39 30 41 33
rect 49 30 51 33
rect 61 30 63 37
rect 71 34 74 37
rect 78 34 79 38
rect 84 39 86 42
rect 94 39 96 42
rect 84 38 96 39
rect 84 37 88 38
rect 71 33 79 34
rect 87 34 88 37
rect 92 37 96 38
rect 92 34 93 37
rect 87 33 93 34
rect 71 30 73 33
rect 101 31 103 42
rect 97 30 103 31
rect 97 26 98 30
rect 102 26 103 30
rect 97 25 103 26
rect 17 8 19 13
rect 27 8 29 13
rect 39 8 41 13
rect 49 8 51 13
rect 61 8 63 13
rect 71 8 73 13
<< ndiffusion >>
rect 31 24 39 30
rect 8 13 17 24
rect 19 22 27 24
rect 19 18 21 22
rect 25 18 27 22
rect 19 13 27 18
rect 29 13 39 24
rect 41 22 49 30
rect 41 18 43 22
rect 47 18 49 22
rect 41 13 49 18
rect 51 13 61 30
rect 63 22 71 30
rect 63 18 65 22
rect 69 18 71 22
rect 63 13 71 18
rect 73 18 81 30
rect 73 14 75 18
rect 79 14 81 18
rect 73 13 81 14
rect 8 12 15 13
rect 8 8 10 12
rect 14 8 15 12
rect 31 12 37 13
rect 31 8 32 12
rect 36 8 37 12
rect 53 12 59 13
rect 53 8 54 12
rect 58 8 59 12
rect 8 7 15 8
rect 31 7 37 8
rect 53 7 59 8
<< pdiffusion >>
rect 2 69 9 70
rect 2 65 3 69
rect 7 65 9 69
rect 2 62 9 65
rect 2 58 3 62
rect 7 58 9 62
rect 2 42 9 58
rect 11 42 16 70
rect 18 62 26 70
rect 18 58 20 62
rect 24 58 26 62
rect 18 54 26 58
rect 18 50 20 54
rect 24 50 26 54
rect 18 42 26 50
rect 28 42 33 70
rect 35 69 43 70
rect 35 65 37 69
rect 41 65 43 69
rect 35 62 43 65
rect 35 58 37 62
rect 41 58 43 62
rect 35 42 43 58
rect 45 42 50 70
rect 52 61 60 70
rect 52 57 54 61
rect 58 57 60 61
rect 52 54 60 57
rect 52 50 54 54
rect 58 50 60 54
rect 52 42 60 50
rect 62 42 67 70
rect 69 69 77 70
rect 69 65 71 69
rect 75 65 77 69
rect 69 62 77 65
rect 69 58 71 62
rect 75 58 77 62
rect 69 42 77 58
rect 79 42 84 70
rect 86 62 94 70
rect 86 58 88 62
rect 92 58 94 62
rect 86 54 94 58
rect 86 50 88 54
rect 92 50 94 54
rect 86 42 94 50
rect 96 42 101 70
rect 103 69 110 70
rect 103 65 105 69
rect 109 65 110 69
rect 103 62 110 65
rect 103 58 105 62
rect 109 58 110 62
rect 103 42 110 58
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect 118 78 122 82
rect 126 78 130 82
rect -2 69 130 78
rect -2 68 3 69
rect 2 65 3 68
rect 7 68 37 69
rect 7 65 8 68
rect 2 62 8 65
rect 36 65 37 68
rect 41 68 71 69
rect 41 65 42 68
rect 2 58 3 62
rect 7 58 8 62
rect 18 62 24 63
rect 18 58 20 62
rect 36 62 42 65
rect 70 65 71 68
rect 75 68 105 69
rect 75 65 76 68
rect 70 62 76 65
rect 104 65 105 68
rect 109 68 130 69
rect 109 65 110 68
rect 36 58 37 62
rect 41 58 42 62
rect 54 61 58 62
rect 18 54 24 58
rect 70 58 71 62
rect 75 58 76 62
rect 88 62 94 63
rect 92 58 94 62
rect 104 62 110 65
rect 104 58 105 62
rect 109 58 110 62
rect 54 54 58 57
rect 88 54 94 58
rect 2 50 20 54
rect 24 50 54 54
rect 58 50 88 54
rect 92 50 95 54
rect 2 22 6 50
rect 27 42 88 46
rect 27 38 31 42
rect 49 38 55 42
rect 23 34 24 38
rect 28 34 31 38
rect 37 34 38 38
rect 42 34 43 38
rect 49 34 50 38
rect 54 34 55 38
rect 73 34 74 38
rect 78 34 79 38
rect 84 34 88 42
rect 92 34 95 38
rect 14 32 18 33
rect 37 30 43 34
rect 73 30 79 34
rect 18 28 98 30
rect 14 26 98 28
rect 102 26 103 30
rect 2 18 21 22
rect 25 18 43 22
rect 47 18 65 22
rect 69 18 71 22
rect 75 18 79 19
rect 75 12 79 14
rect -2 8 10 12
rect 14 8 32 12
rect 36 8 54 12
rect 58 8 130 12
rect -2 2 130 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 122 2
rect 126 -2 130 2
<< ntransistor >>
rect 17 13 19 24
rect 27 13 29 24
rect 39 13 41 30
rect 49 13 51 30
rect 61 13 63 30
rect 71 13 73 30
<< ptransistor >>
rect 9 42 11 70
rect 16 42 18 70
rect 26 42 28 70
rect 33 42 35 70
rect 43 42 45 70
rect 50 42 52 70
rect 60 42 62 70
rect 67 42 69 70
rect 77 42 79 70
rect 84 42 86 70
rect 94 42 96 70
rect 101 42 103 70
<< polycontact >>
rect 24 34 28 38
rect 38 34 42 38
rect 50 34 54 38
rect 14 28 18 32
rect 74 34 78 38
rect 88 34 92 38
rect 98 26 102 30
<< ndcontact >>
rect 21 18 25 22
rect 43 18 47 22
rect 65 18 69 22
rect 75 14 79 18
rect 10 8 14 12
rect 32 8 36 12
rect 54 8 58 12
<< pdcontact >>
rect 3 65 7 69
rect 3 58 7 62
rect 20 58 24 62
rect 20 50 24 54
rect 37 65 41 69
rect 37 58 41 62
rect 54 57 58 61
rect 54 50 58 54
rect 71 65 75 69
rect 71 58 75 62
rect 88 58 92 62
rect 88 50 92 54
rect 105 65 109 69
rect 105 58 109 62
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
rect 90 -2 94 2
rect 98 -2 102 2
rect 106 -2 110 2
rect 114 -2 118 2
rect 122 -2 126 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
rect 90 78 94 82
rect 98 78 102 82
rect 106 78 110 82
rect 114 78 118 82
rect 122 78 126 82
<< psubstratepdiff >>
rect 0 2 128 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 122 2
rect 126 -2 128 2
rect 0 -3 128 -2
<< nsubstratendiff >>
rect 0 82 128 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect 118 78 122 82
rect 126 78 128 82
rect 0 77 128 78
<< labels >>
rlabel metal1 12 20 12 20 6 z
rlabel metal1 20 20 20 20 6 z
rlabel metal1 20 28 20 28 6 a
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 52 12 52 6 z
rlabel metal1 20 56 20 56 6 z
rlabel metal1 28 20 28 20 6 z
rlabel metal1 28 28 28 28 6 a
rlabel metal1 36 20 36 20 6 z
rlabel metal1 36 28 36 28 6 a
rlabel ndcontact 44 20 44 20 6 z
rlabel metal1 44 28 44 28 6 a
rlabel metal1 28 36 28 36 6 b
rlabel metal1 36 44 36 44 6 b
rlabel metal1 44 44 44 44 6 b
rlabel metal1 28 52 28 52 6 z
rlabel metal1 36 52 36 52 6 z
rlabel metal1 44 52 44 52 6 z
rlabel metal1 64 6 64 6 6 vss
rlabel metal1 52 20 52 20 6 z
rlabel metal1 52 28 52 28 6 a
rlabel metal1 60 20 60 20 6 z
rlabel metal1 60 28 60 28 6 a
rlabel ndcontact 68 20 68 20 6 z
rlabel metal1 68 28 68 28 6 a
rlabel metal1 52 40 52 40 6 b
rlabel metal1 60 44 60 44 6 b
rlabel metal1 68 44 68 44 6 b
rlabel metal1 60 52 60 52 6 z
rlabel metal1 68 52 68 52 6 z
rlabel metal1 52 52 52 52 6 z
rlabel metal1 64 74 64 74 6 vdd
rlabel polycontact 100 28 100 28 6 a
rlabel metal1 84 28 84 28 6 a
rlabel metal1 92 28 92 28 6 a
rlabel metal1 76 32 76 32 6 a
rlabel metal1 76 44 76 44 6 b
rlabel metal1 84 44 84 44 6 b
rlabel metal1 92 36 92 36 6 b
rlabel metal1 84 52 84 52 6 z
rlabel metal1 76 52 76 52 6 z
rlabel metal1 92 56 92 56 6 z
<< end >>
