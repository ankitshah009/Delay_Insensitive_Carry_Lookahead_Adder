magic
tech scmos
timestamp 1179386783
<< checkpaint >>
rect -22 -25 174 105
<< ab >>
rect 0 0 152 80
<< pwell >>
rect -4 -7 156 36
<< nwell >>
rect -4 36 156 87
<< polysilicon >>
rect 9 70 11 74
rect 16 70 18 74
rect 26 70 28 74
rect 33 70 35 74
rect 43 70 45 74
rect 50 70 52 74
rect 60 70 62 74
rect 67 70 69 74
rect 77 70 79 74
rect 84 70 86 74
rect 94 70 96 74
rect 101 70 103 74
rect 111 70 113 74
rect 118 70 120 74
rect 128 61 130 65
rect 135 61 137 65
rect 9 33 11 42
rect 16 39 18 42
rect 26 39 28 42
rect 33 39 35 42
rect 43 39 45 42
rect 50 39 52 42
rect 60 39 62 42
rect 16 38 29 39
rect 16 37 24 38
rect 23 34 24 37
rect 28 34 29 38
rect 33 38 45 39
rect 33 37 38 38
rect 23 33 29 34
rect 9 32 15 33
rect 9 28 10 32
rect 14 28 15 32
rect 27 30 29 33
rect 37 34 38 37
rect 42 36 45 38
rect 49 38 62 39
rect 42 34 43 36
rect 37 33 43 34
rect 49 34 50 38
rect 54 37 62 38
rect 67 39 69 42
rect 77 39 79 42
rect 67 38 79 39
rect 54 34 56 37
rect 49 33 56 34
rect 67 34 74 38
rect 78 34 79 38
rect 84 39 86 42
rect 94 39 96 42
rect 84 38 96 39
rect 84 36 90 38
rect 67 33 79 34
rect 86 34 90 36
rect 94 36 96 38
rect 94 34 95 36
rect 86 33 95 34
rect 37 30 39 33
rect 9 27 15 28
rect 54 28 56 33
rect 64 31 69 33
rect 64 28 66 31
rect 76 30 78 33
rect 86 30 88 33
rect 101 31 103 42
rect 111 31 113 42
rect 118 39 120 42
rect 128 39 130 42
rect 118 38 130 39
rect 118 34 119 38
rect 123 37 130 38
rect 123 34 124 37
rect 118 33 124 34
rect 135 31 137 42
rect 101 30 113 31
rect 101 29 105 30
rect 104 26 105 29
rect 109 29 113 30
rect 129 30 137 31
rect 109 26 110 29
rect 104 25 110 26
rect 129 26 130 30
rect 134 26 137 30
rect 129 25 137 26
rect 27 6 29 10
rect 37 6 39 10
rect 54 6 56 10
rect 64 6 66 10
rect 76 6 78 10
rect 86 6 88 10
<< ndiffusion >>
rect 19 15 27 30
rect 19 11 21 15
rect 25 11 27 15
rect 19 10 27 11
rect 29 22 37 30
rect 29 18 31 22
rect 35 18 37 22
rect 29 10 37 18
rect 39 28 51 30
rect 71 28 76 30
rect 39 15 54 28
rect 39 11 44 15
rect 48 11 54 15
rect 39 10 54 11
rect 56 22 64 28
rect 56 18 58 22
rect 62 18 64 22
rect 56 10 64 18
rect 66 15 76 28
rect 66 11 69 15
rect 73 11 76 15
rect 66 10 76 11
rect 78 22 86 30
rect 78 18 80 22
rect 84 18 86 22
rect 78 10 86 18
rect 88 22 96 30
rect 88 18 90 22
rect 94 18 96 22
rect 88 15 96 18
rect 88 11 90 15
rect 94 11 96 15
rect 88 10 96 11
<< pdiffusion >>
rect 2 69 9 70
rect 2 65 3 69
rect 7 65 9 69
rect 2 62 9 65
rect 2 58 3 62
rect 7 58 9 62
rect 2 42 9 58
rect 11 42 16 70
rect 18 62 26 70
rect 18 58 20 62
rect 24 58 26 62
rect 18 54 26 58
rect 18 50 20 54
rect 24 50 26 54
rect 18 42 26 50
rect 28 42 33 70
rect 35 69 43 70
rect 35 65 37 69
rect 41 65 43 69
rect 35 62 43 65
rect 35 58 37 62
rect 41 58 43 62
rect 35 42 43 58
rect 45 42 50 70
rect 52 61 60 70
rect 52 57 54 61
rect 58 57 60 61
rect 52 54 60 57
rect 52 50 54 54
rect 58 50 60 54
rect 52 42 60 50
rect 62 42 67 70
rect 69 69 77 70
rect 69 65 71 69
rect 75 65 77 69
rect 69 62 77 65
rect 69 58 71 62
rect 75 58 77 62
rect 69 42 77 58
rect 79 42 84 70
rect 86 62 94 70
rect 86 58 88 62
rect 92 58 94 62
rect 86 54 94 58
rect 86 50 88 54
rect 92 50 94 54
rect 86 42 94 50
rect 96 42 101 70
rect 103 69 111 70
rect 103 65 105 69
rect 109 65 111 69
rect 103 62 111 65
rect 103 58 105 62
rect 109 58 111 62
rect 103 42 111 58
rect 113 42 118 70
rect 120 61 125 70
rect 120 54 128 61
rect 120 50 122 54
rect 126 50 128 54
rect 120 47 128 50
rect 120 43 122 47
rect 126 43 128 47
rect 120 42 128 43
rect 130 42 135 61
rect 137 60 145 61
rect 137 56 139 60
rect 143 56 145 60
rect 137 53 145 56
rect 137 49 139 53
rect 143 49 145 53
rect 137 42 145 49
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect 118 78 122 82
rect 126 78 130 82
rect 134 78 138 82
rect 142 78 146 82
rect 150 78 154 82
rect -2 69 154 78
rect -2 68 3 69
rect 2 65 3 68
rect 7 68 37 69
rect 7 65 8 68
rect 2 62 8 65
rect 36 65 37 68
rect 41 68 71 69
rect 41 65 42 68
rect 2 58 3 62
rect 7 58 8 62
rect 18 62 24 63
rect 18 58 20 62
rect 36 62 42 65
rect 70 65 71 68
rect 75 68 105 69
rect 75 65 76 68
rect 70 62 76 65
rect 104 65 105 68
rect 109 68 154 69
rect 109 65 110 68
rect 36 58 37 62
rect 41 58 42 62
rect 54 61 58 62
rect 18 54 24 58
rect 70 58 71 62
rect 75 58 76 62
rect 88 62 94 63
rect 92 58 94 62
rect 104 62 110 65
rect 104 58 105 62
rect 109 58 110 62
rect 138 60 144 68
rect 54 54 58 57
rect 88 54 94 58
rect 138 56 139 60
rect 143 56 144 60
rect 2 50 20 54
rect 24 50 54 54
rect 58 50 88 54
rect 92 50 122 54
rect 126 50 127 54
rect 2 22 6 50
rect 121 47 127 50
rect 138 53 144 56
rect 138 49 139 53
rect 143 49 144 53
rect 25 42 95 46
rect 121 43 122 47
rect 126 43 127 47
rect 121 42 127 43
rect 25 38 31 42
rect 49 38 55 42
rect 89 38 95 42
rect 23 34 24 38
rect 28 34 31 38
rect 37 34 38 38
rect 42 34 43 38
rect 49 34 50 38
rect 54 34 55 38
rect 73 34 74 38
rect 78 34 79 38
rect 89 34 90 38
rect 94 34 119 38
rect 123 34 127 38
rect 10 32 14 33
rect 37 30 43 34
rect 73 30 79 34
rect 14 28 105 30
rect 10 26 105 28
rect 109 26 130 30
rect 134 26 135 30
rect 2 18 31 22
rect 35 18 58 22
rect 62 18 80 22
rect 84 18 85 22
rect 89 18 90 22
rect 94 18 95 22
rect 89 15 95 18
rect 20 12 21 15
rect -2 11 21 12
rect 25 12 26 15
rect 43 12 44 15
rect 25 11 44 12
rect 48 12 49 15
rect 68 12 69 15
rect 48 11 69 12
rect 73 12 74 15
rect 89 12 90 15
rect 73 11 90 12
rect 94 12 95 15
rect 94 11 154 12
rect -2 2 154 11
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 122 2
rect 126 -2 130 2
rect 134 -2 138 2
rect 142 -2 146 2
rect 150 -2 154 2
<< ntransistor >>
rect 27 10 29 30
rect 37 10 39 30
rect 54 10 56 28
rect 64 10 66 28
rect 76 10 78 30
rect 86 10 88 30
<< ptransistor >>
rect 9 42 11 70
rect 16 42 18 70
rect 26 42 28 70
rect 33 42 35 70
rect 43 42 45 70
rect 50 42 52 70
rect 60 42 62 70
rect 67 42 69 70
rect 77 42 79 70
rect 84 42 86 70
rect 94 42 96 70
rect 101 42 103 70
rect 111 42 113 70
rect 118 42 120 70
rect 128 42 130 61
rect 135 42 137 61
<< polycontact >>
rect 24 34 28 38
rect 10 28 14 32
rect 38 34 42 38
rect 50 34 54 38
rect 74 34 78 38
rect 90 34 94 38
rect 119 34 123 38
rect 105 26 109 30
rect 130 26 134 30
<< ndcontact >>
rect 21 11 25 15
rect 31 18 35 22
rect 44 11 48 15
rect 58 18 62 22
rect 69 11 73 15
rect 80 18 84 22
rect 90 18 94 22
rect 90 11 94 15
<< pdcontact >>
rect 3 65 7 69
rect 3 58 7 62
rect 20 58 24 62
rect 20 50 24 54
rect 37 65 41 69
rect 37 58 41 62
rect 54 57 58 61
rect 54 50 58 54
rect 71 65 75 69
rect 71 58 75 62
rect 88 58 92 62
rect 88 50 92 54
rect 105 65 109 69
rect 105 58 109 62
rect 122 50 126 54
rect 122 43 126 47
rect 139 56 143 60
rect 139 49 143 53
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
rect 90 -2 94 2
rect 98 -2 102 2
rect 106 -2 110 2
rect 114 -2 118 2
rect 122 -2 126 2
rect 130 -2 134 2
rect 138 -2 142 2
rect 146 -2 150 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
rect 90 78 94 82
rect 98 78 102 82
rect 106 78 110 82
rect 114 78 118 82
rect 122 78 126 82
rect 130 78 134 82
rect 138 78 142 82
rect 146 78 150 82
<< psubstratepdiff >>
rect 0 2 152 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 122 2
rect 126 -2 130 2
rect 134 -2 138 2
rect 142 -2 146 2
rect 150 -2 152 2
rect 0 -3 152 -2
<< nsubstratendiff >>
rect 0 82 152 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect 118 78 122 82
rect 126 78 130 82
rect 134 78 138 82
rect 142 78 146 82
rect 150 78 152 82
rect 0 77 152 78
<< labels >>
rlabel metal1 20 20 20 20 6 z
rlabel metal1 12 20 12 20 6 z
rlabel metal1 20 28 20 28 6 a
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 52 12 52 6 z
rlabel metal1 20 56 20 56 6 z
rlabel metal1 44 20 44 20 6 z
rlabel metal1 36 20 36 20 6 z
rlabel metal1 28 20 28 20 6 z
rlabel metal1 28 28 28 28 6 a
rlabel metal1 36 28 36 28 6 a
rlabel metal1 44 28 44 28 6 a
rlabel metal1 28 36 28 36 6 b
rlabel metal1 36 44 36 44 6 b
rlabel metal1 44 44 44 44 6 b
rlabel metal1 28 52 28 52 6 z
rlabel metal1 36 52 36 52 6 z
rlabel metal1 44 52 44 52 6 z
rlabel metal1 52 20 52 20 6 z
rlabel metal1 68 20 68 20 6 z
rlabel ndcontact 60 20 60 20 6 z
rlabel metal1 60 28 60 28 6 a
rlabel metal1 68 28 68 28 6 a
rlabel metal1 52 28 52 28 6 a
rlabel metal1 60 44 60 44 6 b
rlabel metal1 68 44 68 44 6 b
rlabel metal1 52 40 52 40 6 b
rlabel metal1 52 52 52 52 6 z
rlabel metal1 60 52 60 52 6 z
rlabel metal1 68 52 68 52 6 z
rlabel metal1 76 6 76 6 6 vss
rlabel metal1 76 20 76 20 6 z
rlabel metal1 84 28 84 28 6 a
rlabel metal1 92 28 92 28 6 a
rlabel metal1 100 28 100 28 6 a
rlabel metal1 76 32 76 32 6 a
rlabel metal1 100 36 100 36 6 b
rlabel metal1 84 44 84 44 6 b
rlabel metal1 92 40 92 40 6 b
rlabel metal1 76 44 76 44 6 b
rlabel metal1 76 52 76 52 6 z
rlabel metal1 100 52 100 52 6 z
rlabel metal1 84 52 84 52 6 z
rlabel metal1 92 56 92 56 6 z
rlabel metal1 76 74 76 74 6 vdd
rlabel polycontact 108 28 108 28 6 a
rlabel metal1 116 28 116 28 6 a
rlabel metal1 124 28 124 28 6 a
rlabel metal1 124 36 124 36 6 b
rlabel metal1 116 36 116 36 6 b
rlabel metal1 108 36 108 36 6 b
rlabel metal1 124 48 124 48 6 z
rlabel metal1 108 52 108 52 6 z
rlabel metal1 116 52 116 52 6 z
rlabel polycontact 132 28 132 28 6 a
<< end >>
