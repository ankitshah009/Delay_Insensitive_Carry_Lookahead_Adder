magic
tech scmos
timestamp 1179386130
<< checkpaint >>
rect -22 -22 246 94
<< ab >>
rect 0 0 224 72
<< pwell >>
rect -4 -4 228 32
<< nwell >>
rect -4 32 228 76
<< polysilicon >>
rect 9 66 11 70
rect 19 66 21 70
rect 29 66 31 70
rect 39 66 41 70
rect 59 67 81 69
rect 59 61 61 67
rect 69 64 71 67
rect 79 64 81 67
rect 139 68 205 70
rect 139 65 141 68
rect 49 59 61 61
rect 49 56 51 59
rect 59 56 61 59
rect 89 60 91 65
rect 99 63 141 65
rect 99 60 101 63
rect 109 60 111 63
rect 119 60 121 63
rect 129 60 131 63
rect 139 60 141 63
rect 149 60 151 64
rect 163 60 165 64
rect 173 60 175 64
rect 183 60 185 64
rect 193 60 195 64
rect 203 60 205 68
rect 213 54 215 59
rect 9 35 11 38
rect 19 35 21 38
rect 29 35 31 38
rect 39 35 41 38
rect 9 34 41 35
rect 49 34 51 38
rect 59 34 61 38
rect 69 34 71 38
rect 79 35 81 38
rect 89 35 91 38
rect 79 34 91 35
rect 99 34 101 38
rect 109 34 111 38
rect 119 35 121 38
rect 119 34 125 35
rect 9 30 10 34
rect 14 30 18 34
rect 22 30 41 34
rect 79 30 84 34
rect 88 30 91 34
rect 119 30 120 34
rect 124 30 125 34
rect 129 33 131 38
rect 139 33 141 38
rect 149 35 151 38
rect 163 35 165 38
rect 173 35 175 38
rect 183 35 185 38
rect 193 35 195 38
rect 149 34 195 35
rect 9 29 41 30
rect 19 26 21 29
rect 29 26 31 29
rect 39 26 41 29
rect 49 26 51 30
rect 59 26 61 30
rect 69 26 71 30
rect 79 29 91 30
rect 79 26 81 29
rect 89 26 91 29
rect 99 26 101 30
rect 109 26 111 30
rect 119 29 125 30
rect 149 30 150 34
rect 154 30 158 34
rect 162 33 195 34
rect 203 35 205 38
rect 213 35 215 38
rect 162 30 181 33
rect 149 29 181 30
rect 79 9 81 13
rect 89 10 91 13
rect 99 10 101 13
rect 109 10 111 13
rect 89 8 111 10
rect 19 3 21 8
rect 29 3 31 8
rect 39 3 41 8
rect 49 4 51 8
rect 59 4 61 8
rect 69 4 71 8
rect 120 4 122 29
rect 149 26 151 29
rect 159 26 161 29
rect 169 26 171 29
rect 179 26 181 29
rect 203 29 215 35
rect 203 26 205 29
rect 213 26 215 29
rect 49 2 122 4
rect 149 7 151 12
rect 159 7 161 12
rect 169 7 171 12
rect 179 7 181 12
rect 203 10 205 15
rect 213 11 215 15
<< ndiffusion >>
rect 11 21 19 26
rect 11 17 13 21
rect 17 17 19 21
rect 11 13 19 17
rect 11 9 13 13
rect 17 9 19 13
rect 11 8 19 9
rect 21 25 29 26
rect 21 21 23 25
rect 27 21 29 25
rect 21 18 29 21
rect 21 14 23 18
rect 27 14 29 18
rect 21 8 29 14
rect 31 13 39 26
rect 31 9 33 13
rect 37 9 39 13
rect 31 8 39 9
rect 41 25 49 26
rect 41 21 43 25
rect 47 21 49 25
rect 41 18 49 21
rect 41 14 43 18
rect 47 14 49 18
rect 41 8 49 14
rect 51 25 59 26
rect 51 21 53 25
rect 57 21 59 25
rect 51 8 59 21
rect 61 17 69 26
rect 61 13 63 17
rect 67 13 69 17
rect 61 8 69 13
rect 71 25 79 26
rect 71 21 73 25
rect 77 21 79 25
rect 71 18 79 21
rect 71 14 73 18
rect 77 14 79 18
rect 71 13 79 14
rect 81 18 89 26
rect 81 14 83 18
rect 87 14 89 18
rect 81 13 89 14
rect 91 25 99 26
rect 91 21 93 25
rect 97 21 99 25
rect 91 13 99 21
rect 101 18 109 26
rect 101 14 103 18
rect 107 14 109 18
rect 101 13 109 14
rect 111 25 118 26
rect 111 21 113 25
rect 117 21 118 25
rect 111 20 118 21
rect 111 13 116 20
rect 71 8 76 13
rect 141 12 149 26
rect 151 25 159 26
rect 151 21 153 25
rect 157 21 159 25
rect 151 18 159 21
rect 151 14 153 18
rect 157 14 159 18
rect 151 12 159 14
rect 161 17 169 26
rect 161 13 163 17
rect 167 13 169 17
rect 161 12 169 13
rect 171 25 179 26
rect 171 21 173 25
rect 177 21 179 25
rect 171 18 179 21
rect 171 14 173 18
rect 177 14 179 18
rect 171 12 179 14
rect 181 25 189 26
rect 181 21 183 25
rect 187 21 189 25
rect 181 17 189 21
rect 181 13 183 17
rect 187 13 189 17
rect 195 20 203 26
rect 195 16 197 20
rect 201 16 203 20
rect 195 15 203 16
rect 205 25 213 26
rect 205 21 207 25
rect 211 21 213 25
rect 205 15 213 21
rect 215 20 222 26
rect 215 16 217 20
rect 221 16 222 20
rect 215 15 222 16
rect 181 12 189 13
rect 141 8 147 12
rect 141 4 142 8
rect 146 4 147 8
rect 141 3 147 4
<< pdiffusion >>
rect 4 51 9 66
rect 2 50 9 51
rect 2 46 3 50
rect 7 46 9 50
rect 2 43 9 46
rect 2 39 3 43
rect 7 39 9 43
rect 2 38 9 39
rect 11 65 19 66
rect 11 61 13 65
rect 17 61 19 65
rect 11 58 19 61
rect 11 54 13 58
rect 17 54 19 58
rect 11 38 19 54
rect 21 50 29 66
rect 21 46 23 50
rect 27 46 29 50
rect 21 43 29 46
rect 21 39 23 43
rect 27 39 29 43
rect 21 38 29 39
rect 31 65 39 66
rect 31 61 33 65
rect 37 61 39 65
rect 31 58 39 61
rect 31 54 33 58
rect 37 54 39 58
rect 31 38 39 54
rect 41 56 46 66
rect 64 56 69 64
rect 41 50 49 56
rect 41 46 43 50
rect 47 46 49 50
rect 41 43 49 46
rect 41 39 43 43
rect 47 39 49 43
rect 41 38 49 39
rect 51 50 59 56
rect 51 46 53 50
rect 57 46 59 50
rect 51 43 59 46
rect 51 39 53 43
rect 57 39 59 43
rect 51 38 59 39
rect 61 55 69 56
rect 61 51 63 55
rect 67 51 69 55
rect 61 48 69 51
rect 61 44 63 48
rect 67 44 69 48
rect 61 38 69 44
rect 71 50 79 64
rect 71 46 73 50
rect 77 46 79 50
rect 71 43 79 46
rect 71 39 73 43
rect 77 39 79 43
rect 71 38 79 39
rect 81 60 86 64
rect 81 59 89 60
rect 81 55 83 59
rect 87 55 89 59
rect 81 38 89 55
rect 91 43 99 60
rect 91 39 93 43
rect 97 39 99 43
rect 91 38 99 39
rect 101 51 109 60
rect 101 47 103 51
rect 107 47 109 51
rect 101 38 109 47
rect 111 43 119 60
rect 111 39 113 43
rect 117 39 119 43
rect 111 38 119 39
rect 121 51 129 60
rect 121 47 123 51
rect 127 47 129 51
rect 121 38 129 47
rect 131 43 139 60
rect 131 39 133 43
rect 137 39 139 43
rect 131 38 139 39
rect 141 50 149 60
rect 141 46 143 50
rect 147 46 149 50
rect 141 43 149 46
rect 141 39 143 43
rect 147 39 149 43
rect 141 38 149 39
rect 151 59 163 60
rect 151 55 157 59
rect 161 55 163 59
rect 151 38 163 55
rect 165 43 173 60
rect 165 39 167 43
rect 171 39 173 43
rect 165 38 173 39
rect 175 59 183 60
rect 175 55 177 59
rect 181 55 183 59
rect 175 38 183 55
rect 185 43 193 60
rect 185 39 187 43
rect 191 39 193 43
rect 185 38 193 39
rect 195 59 203 60
rect 195 55 197 59
rect 201 55 203 59
rect 195 38 203 55
rect 205 54 210 60
rect 205 50 213 54
rect 205 46 207 50
rect 211 46 213 50
rect 205 43 213 46
rect 205 39 207 43
rect 211 39 213 43
rect 205 38 213 39
rect 215 53 222 54
rect 215 49 217 53
rect 221 49 222 53
rect 215 45 222 49
rect 215 41 217 45
rect 221 41 222 45
rect 215 38 222 41
<< metal1 >>
rect -2 68 226 72
rect -2 65 51 68
rect -2 64 13 65
rect 17 64 33 65
rect 13 58 17 61
rect 13 53 17 54
rect 37 64 51 65
rect 55 64 216 68
rect 220 64 226 68
rect 33 58 37 61
rect 157 59 161 64
rect 33 53 37 54
rect 43 55 83 59
rect 87 55 88 59
rect 93 55 154 59
rect 3 50 7 51
rect 3 43 7 46
rect 23 50 27 51
rect 23 43 27 46
rect 7 39 23 42
rect 43 50 47 55
rect 43 43 47 46
rect 27 39 43 42
rect 3 38 47 39
rect 2 34 22 35
rect 2 30 10 34
rect 14 30 18 34
rect 2 29 22 30
rect 2 13 6 29
rect 43 26 47 38
rect 23 25 47 26
rect 13 21 17 22
rect 13 13 17 17
rect 27 22 43 25
rect 23 18 27 21
rect 43 18 47 21
rect 53 50 57 51
rect 53 43 57 46
rect 63 48 67 51
rect 63 43 67 44
rect 73 50 78 52
rect 93 51 97 55
rect 150 51 154 55
rect 157 54 161 55
rect 177 59 181 64
rect 196 59 202 64
rect 196 55 197 59
rect 201 55 202 59
rect 177 54 181 55
rect 217 53 221 64
rect 77 46 78 50
rect 73 43 78 46
rect 53 26 57 39
rect 77 39 78 43
rect 73 26 78 39
rect 84 47 97 51
rect 102 47 103 51
rect 107 47 123 51
rect 127 50 147 51
rect 127 47 143 50
rect 84 34 88 47
rect 142 46 143 47
rect 150 50 211 51
rect 150 47 207 50
rect 142 43 147 46
rect 207 43 211 46
rect 92 39 93 43
rect 97 42 98 43
rect 112 42 113 43
rect 97 39 113 42
rect 117 42 118 43
rect 132 42 133 43
rect 117 39 133 42
rect 137 39 138 43
rect 142 39 143 43
rect 147 39 167 43
rect 171 39 187 43
rect 191 39 192 43
rect 217 45 221 49
rect 217 40 221 41
rect 92 38 138 39
rect 84 29 88 30
rect 98 26 102 38
rect 146 34 166 35
rect 119 30 120 34
rect 124 30 135 34
rect 53 25 119 26
rect 57 22 73 25
rect 53 20 57 21
rect 77 22 93 25
rect 77 21 78 22
rect 92 21 93 22
rect 97 22 113 25
rect 97 21 98 22
rect 112 21 113 22
rect 117 21 119 25
rect 129 22 135 30
rect 146 30 150 34
rect 154 30 158 34
rect 162 30 166 34
rect 146 29 166 30
rect 146 21 150 29
rect 173 26 177 39
rect 153 25 177 26
rect 157 22 173 25
rect 157 21 158 22
rect 73 18 78 21
rect 153 18 158 21
rect 173 18 177 21
rect 47 14 63 17
rect 23 13 27 14
rect 33 13 37 14
rect 43 13 63 14
rect 67 13 68 17
rect 77 14 78 18
rect 82 14 83 18
rect 87 14 103 18
rect 107 14 153 18
rect 157 14 158 18
rect 163 17 167 18
rect 73 13 78 14
rect 173 13 177 14
rect 183 25 187 26
rect 207 25 211 39
rect 183 17 187 21
rect 13 8 17 9
rect 33 8 37 9
rect 163 8 167 13
rect 183 8 187 13
rect 197 20 201 21
rect 207 20 211 21
rect 217 20 221 21
rect 197 8 201 16
rect 217 8 221 16
rect -2 4 125 8
rect 129 4 132 8
rect 136 4 142 8
rect 146 4 208 8
rect 212 4 216 8
rect 220 4 226 8
rect -2 0 226 4
<< ntransistor >>
rect 19 8 21 26
rect 29 8 31 26
rect 39 8 41 26
rect 49 8 51 26
rect 59 8 61 26
rect 69 8 71 26
rect 79 13 81 26
rect 89 13 91 26
rect 99 13 101 26
rect 109 13 111 26
rect 149 12 151 26
rect 159 12 161 26
rect 169 12 171 26
rect 179 12 181 26
rect 203 15 205 26
rect 213 15 215 26
<< ptransistor >>
rect 9 38 11 66
rect 19 38 21 66
rect 29 38 31 66
rect 39 38 41 66
rect 49 38 51 56
rect 59 38 61 56
rect 69 38 71 64
rect 79 38 81 64
rect 89 38 91 60
rect 99 38 101 60
rect 109 38 111 60
rect 119 38 121 60
rect 129 38 131 60
rect 139 38 141 60
rect 149 38 151 60
rect 163 38 165 60
rect 173 38 175 60
rect 183 38 185 60
rect 193 38 195 60
rect 203 38 205 60
rect 213 38 215 54
<< polycontact >>
rect 10 30 14 34
rect 18 30 22 34
rect 84 30 88 34
rect 120 30 124 34
rect 150 30 154 34
rect 158 30 162 34
<< ndcontact >>
rect 13 17 17 21
rect 13 9 17 13
rect 23 21 27 25
rect 23 14 27 18
rect 33 9 37 13
rect 43 21 47 25
rect 43 14 47 18
rect 53 21 57 25
rect 63 13 67 17
rect 73 21 77 25
rect 73 14 77 18
rect 83 14 87 18
rect 93 21 97 25
rect 103 14 107 18
rect 113 21 117 25
rect 153 21 157 25
rect 153 14 157 18
rect 163 13 167 17
rect 173 21 177 25
rect 173 14 177 18
rect 183 21 187 25
rect 183 13 187 17
rect 197 16 201 20
rect 207 21 211 25
rect 217 16 221 20
rect 142 4 146 8
<< pdcontact >>
rect 3 46 7 50
rect 3 39 7 43
rect 13 61 17 65
rect 13 54 17 58
rect 23 46 27 50
rect 23 39 27 43
rect 33 61 37 65
rect 33 54 37 58
rect 43 46 47 50
rect 43 39 47 43
rect 53 46 57 50
rect 53 39 57 43
rect 63 51 67 55
rect 63 44 67 48
rect 73 46 77 50
rect 73 39 77 43
rect 83 55 87 59
rect 93 39 97 43
rect 103 47 107 51
rect 113 39 117 43
rect 123 47 127 51
rect 133 39 137 43
rect 143 46 147 50
rect 143 39 147 43
rect 157 55 161 59
rect 167 39 171 43
rect 177 55 181 59
rect 187 39 191 43
rect 197 55 201 59
rect 207 46 211 50
rect 207 39 211 43
rect 217 49 221 53
rect 217 41 221 45
<< psubstratepcontact >>
rect 125 4 129 8
rect 132 4 136 8
rect 208 4 212 8
rect 216 4 220 8
<< nsubstratencontact >>
rect 51 64 55 68
rect 216 64 220 68
<< psubstratepdiff >>
rect 124 8 137 9
rect 124 4 125 8
rect 129 4 132 8
rect 136 4 137 8
rect 124 3 137 4
rect 207 8 221 9
rect 207 4 208 8
rect 212 4 216 8
rect 220 4 221 8
rect 207 3 221 4
<< nsubstratendiff >>
rect 50 68 56 69
rect 50 64 51 68
rect 55 64 56 68
rect 50 63 56 64
rect 215 68 221 69
rect 215 64 216 68
rect 220 64 221 68
rect 215 63 221 64
<< labels >>
rlabel metal1 25 19 25 19 6 a1n
rlabel metal1 4 24 4 24 6 a1
rlabel polycontact 12 32 12 32 6 a1
rlabel polycontact 20 32 20 32 6 a1
rlabel metal1 5 44 5 44 6 a1n
rlabel metal1 25 44 25 44 6 a1n
rlabel metal1 55 15 55 15 6 a1n
rlabel metal1 60 24 60 24 6 z
rlabel metal1 68 24 68 24 6 z
rlabel metal1 84 24 84 24 6 z
rlabel metal1 76 32 76 32 6 z
rlabel metal1 86 40 86 40 6 sn
rlabel metal1 45 36 45 36 6 a1n
rlabel metal1 65 51 65 51 6 a1n
rlabel metal1 112 4 112 4 6 vss
rlabel metal1 92 24 92 24 6 z
rlabel metal1 108 24 108 24 6 z
rlabel ndcontact 116 24 116 24 6 z
rlabel metal1 100 32 100 32 6 z
rlabel metal1 124 32 124 32 6 s
rlabel metal1 132 28 132 28 6 s
rlabel metal1 108 40 108 40 6 z
rlabel pdcontact 116 40 116 40 6 z
rlabel metal1 124 40 124 40 6 z
rlabel metal1 132 40 132 40 6 z
rlabel metal1 112 68 112 68 6 vdd
rlabel metal1 155 20 155 20 6 a0n
rlabel metal1 120 16 120 16 6 a0n
rlabel metal1 164 32 164 32 6 a0
rlabel metal1 156 32 156 32 6 a0
rlabel metal1 148 28 148 28 6 a0
rlabel metal1 144 45 144 45 6 a0n
rlabel metal1 175 28 175 28 6 a0n
rlabel pdcontact 124 49 124 49 6 a0n
rlabel metal1 167 41 167 41 6 a0n
rlabel metal1 209 35 209 35 6 sn
<< end >>
