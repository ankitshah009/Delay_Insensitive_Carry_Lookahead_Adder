.subckt nr2_x1 a b vdd vss z
*   SPICE3 file   created from nr2_x1.ext -      technology: scmos
m00 w1     b      z      vdd p w=39u  l=2.3636u ad=117p     pd=45u      as=237p     ps=94u
m01 vdd    a      w1     vdd p w=39u  l=2.3636u ad=351p     pd=96u      as=117p     ps=45u
m02 z      b      vss    vss n w=11u  l=2.3636u ad=55p      pd=21u      as=99p      ps=40u
m03 vss    a      z      vss n w=11u  l=2.3636u ad=99p      pd=40u      as=55p      ps=21u
C0  z      b      0.148f
C1  vdd    w1     0.011f
C2  vss    z      0.113f
C3  vss    b      0.025f
C4  vdd    a      0.090f
C5  z      a      0.073f
C6  a      b      0.209f
C7  vdd    z      0.018f
C8  vss    a      0.009f
C9  w1     a      0.012f
C10 vdd    b      0.012f
C13 z      vss    0.019f
C14 a      vss    0.026f
C15 b      vss    0.034f
.ends
