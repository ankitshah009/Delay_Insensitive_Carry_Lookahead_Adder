.subckt an12_x4 i0 i1 q vdd vss
*   SPICE3 file   created from an12_x4.ext -      technology: scmos
m00 vdd    i0     w1     vdd p w=20u  l=2.3636u ad=164.571p pd=41.1429u as=160p     ps=56u
m01 w2     w1     vdd    vdd p w=20u  l=2.3636u ad=100p     pd=30u      as=164.571p ps=41.1429u
m02 vdd    i1     w2     vdd p w=20u  l=2.3636u ad=164.571p pd=41.1429u as=100p     ps=30u
m03 q      w2     vdd    vdd p w=40u  l=2.3636u ad=200p     pd=50u      as=329.143p ps=82.2857u
m04 vdd    w2     q      vdd p w=40u  l=2.3636u ad=329.143p pd=82.2857u as=200p     ps=50u
m05 vss    i0     w1     vss n w=10u  l=2.3636u ad=64.5714p pd=22.2857u as=104p     ps=44u
m06 w3     w1     w2     vss n w=20u  l=2.3636u ad=60p      pd=26u      as=160p     ps=56u
m07 vss    i1     w3     vss n w=20u  l=2.3636u ad=129.143p pd=44.5714u as=60p      ps=26u
m08 q      w2     vss    vss n w=20u  l=2.3636u ad=100p     pd=30u      as=129.143p ps=44.5714u
m09 vss    w2     q      vss n w=20u  l=2.3636u ad=129.143p pd=44.5714u as=100p     ps=30u
C0  w1     w2     0.153f
C1  i0     vdd    0.083f
C2  vdd    w2     0.086f
C3  vss    i1     0.076f
C4  vss    i0     0.044f
C5  vss    w2     0.132f
C6  i1     i0     0.092f
C7  q      vdd    0.209f
C8  w1     vdd    0.054f
C9  i1     w2     0.501f
C10 w3     vss    0.014f
C11 i0     w2     0.173f
C12 vss    q      0.111f
C13 q      i1     0.485f
C14 vss    w1     0.064f
C15 w3     w2     0.012f
C16 i1     w1     0.113f
C17 q      i0     0.057f
C18 vss    vdd    0.005f
C19 i1     vdd    0.146f
C20 w1     i0     0.288f
C21 q      w2     0.200f
C23 q      vss    0.020f
C24 i1     vss    0.043f
C25 w1     vss    0.055f
C26 i0     vss    0.048f
C28 w2     vss    0.064f
.ends
