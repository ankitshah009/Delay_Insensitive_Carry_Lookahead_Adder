magic
tech scmos
timestamp 1179386022
<< checkpaint >>
rect -22 -25 62 105
<< ab >>
rect 0 0 40 80
<< pwell >>
rect -4 -7 44 36
<< nwell >>
rect -4 36 44 87
<< polysilicon >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 9 38 31 39
rect 9 34 16 38
rect 20 37 31 38
rect 20 34 21 37
rect 9 33 21 34
rect 9 30 11 33
rect 19 30 21 33
rect 9 9 11 14
rect 19 9 21 14
<< ndiffusion >>
rect 2 19 9 30
rect 2 15 3 19
rect 7 15 9 19
rect 2 14 9 15
rect 11 29 19 30
rect 11 25 13 29
rect 17 25 19 29
rect 11 22 19 25
rect 11 18 13 22
rect 17 18 19 22
rect 11 14 19 18
rect 21 22 28 30
rect 21 18 23 22
rect 27 18 28 22
rect 21 17 28 18
rect 21 14 27 17
<< pdiffusion >>
rect 4 55 9 70
rect 2 54 9 55
rect 2 50 3 54
rect 7 50 9 54
rect 2 47 9 50
rect 2 43 3 47
rect 7 43 9 47
rect 2 42 9 43
rect 11 69 19 70
rect 11 65 13 69
rect 17 65 19 69
rect 11 62 19 65
rect 11 58 13 62
rect 17 58 19 62
rect 11 42 19 58
rect 21 54 29 70
rect 21 50 23 54
rect 27 50 29 54
rect 21 47 29 50
rect 21 43 23 47
rect 27 43 29 47
rect 21 42 29 43
rect 31 69 38 70
rect 31 65 33 69
rect 37 65 38 69
rect 31 62 38 65
rect 31 58 33 62
rect 37 58 38 62
rect 31 42 38 58
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect -2 69 42 78
rect -2 68 13 69
rect 17 68 33 69
rect 13 62 17 65
rect 32 65 33 68
rect 37 68 42 69
rect 37 65 38 68
rect 32 62 38 65
rect 32 58 33 62
rect 37 58 38 62
rect 13 57 17 58
rect 2 54 7 55
rect 2 50 3 54
rect 2 47 7 50
rect 2 43 3 47
rect 23 54 27 55
rect 23 47 27 50
rect 7 43 23 46
rect 27 43 31 46
rect 2 42 31 43
rect 2 30 6 42
rect 15 34 16 38
rect 20 34 31 38
rect 2 29 17 30
rect 2 25 13 29
rect 25 26 31 34
rect 13 22 17 25
rect 3 19 7 20
rect 13 17 17 18
rect 22 18 23 22
rect 27 18 28 22
rect 3 12 7 15
rect 22 12 28 18
rect -2 2 42 12
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
<< ntransistor >>
rect 9 14 11 30
rect 19 14 21 30
<< ptransistor >>
rect 9 42 11 70
rect 19 42 21 70
rect 29 42 31 70
<< polycontact >>
rect 16 34 20 38
<< ndcontact >>
rect 3 15 7 19
rect 13 25 17 29
rect 13 18 17 22
rect 23 18 27 22
<< pdcontact >>
rect 3 50 7 54
rect 3 43 7 47
rect 13 65 17 69
rect 13 58 17 62
rect 23 50 27 54
rect 23 43 27 47
rect 33 65 37 69
rect 33 58 37 62
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
<< psubstratepdiff >>
rect 0 2 40 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 40 2
rect 0 -3 40 -2
<< nsubstratendiff >>
rect 0 82 40 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 40 82
rect 0 77 40 78
<< labels >>
rlabel metal1 4 40 4 40 6 z
rlabel metal1 12 28 12 28 6 z
rlabel metal1 12 44 12 44 6 z
rlabel metal1 20 6 20 6 6 vss
rlabel metal1 20 36 20 36 6 a
rlabel metal1 28 32 28 32 6 a
rlabel metal1 28 44 28 44 6 z
rlabel metal1 20 44 20 44 6 z
rlabel metal1 20 74 20 74 6 vdd
<< end >>
