magic
tech scmos
timestamp 1180600666
<< checkpaint >>
rect -22 -22 112 122
<< ab >>
rect 0 0 90 100
<< pwell >>
rect -4 -4 94 48
<< nwell >>
rect -4 48 94 104
<< polysilicon >>
rect 11 85 13 89
rect 75 94 77 98
rect 23 85 25 89
rect 31 85 33 89
rect 47 85 49 89
rect 55 85 57 89
rect 11 41 13 65
rect 23 63 25 66
rect 17 62 25 63
rect 17 58 18 62
rect 22 61 25 62
rect 22 58 23 61
rect 17 57 23 58
rect 31 43 33 66
rect 47 57 49 66
rect 55 63 57 66
rect 55 62 63 63
rect 55 61 58 62
rect 57 58 58 61
rect 62 58 63 62
rect 57 57 63 58
rect 47 56 53 57
rect 47 52 48 56
rect 52 52 53 56
rect 47 51 53 52
rect 37 50 43 51
rect 37 46 38 50
rect 42 47 43 50
rect 75 47 77 55
rect 42 46 77 47
rect 37 45 77 46
rect 27 42 33 43
rect 27 41 28 42
rect 11 39 28 41
rect 11 15 13 39
rect 27 38 28 39
rect 32 41 33 42
rect 32 39 49 41
rect 32 38 33 39
rect 27 37 33 38
rect 17 32 23 33
rect 17 28 18 32
rect 22 29 23 32
rect 22 28 25 29
rect 17 27 25 28
rect 23 14 25 27
rect 29 22 35 23
rect 29 18 30 22
rect 34 18 35 22
rect 29 17 35 18
rect 31 14 33 17
rect 47 15 49 39
rect 57 32 63 33
rect 57 29 58 32
rect 55 28 58 29
rect 62 28 63 32
rect 55 27 63 28
rect 55 15 57 27
rect 75 25 77 45
rect 11 2 13 6
rect 23 2 25 6
rect 31 2 33 6
rect 47 2 49 6
rect 55 2 57 6
rect 75 2 77 6
<< ndiffusion >>
rect 3 22 9 25
rect 3 18 4 22
rect 8 18 9 22
rect 3 15 9 18
rect 37 32 45 33
rect 3 6 11 15
rect 13 14 18 15
rect 37 28 38 32
rect 42 28 45 32
rect 37 15 45 28
rect 59 22 75 25
rect 59 18 68 22
rect 72 18 75 22
rect 59 15 75 18
rect 37 14 47 15
rect 13 12 23 14
rect 13 8 16 12
rect 20 8 23 12
rect 13 6 23 8
rect 25 6 31 14
rect 33 6 47 14
rect 49 6 55 15
rect 57 12 75 15
rect 57 8 68 12
rect 72 8 75 12
rect 57 6 75 8
rect 77 22 85 25
rect 77 18 80 22
rect 84 18 85 22
rect 77 6 85 18
<< pdiffusion >>
rect 15 92 21 93
rect 15 88 16 92
rect 20 88 21 92
rect 59 92 75 94
rect 15 85 21 88
rect 59 88 68 92
rect 72 88 75 92
rect 59 85 75 88
rect 3 82 11 85
rect 3 78 4 82
rect 8 78 11 82
rect 3 72 11 78
rect 3 68 4 72
rect 8 68 11 72
rect 3 65 11 68
rect 13 66 23 85
rect 25 66 31 85
rect 33 82 47 85
rect 33 78 38 82
rect 42 78 47 82
rect 33 72 47 78
rect 33 68 38 72
rect 42 68 47 72
rect 33 66 47 68
rect 49 66 55 85
rect 57 82 75 85
rect 57 78 68 82
rect 72 78 75 82
rect 57 72 75 78
rect 57 68 68 72
rect 72 68 75 72
rect 57 66 75 68
rect 13 65 18 66
rect 59 65 75 66
rect 67 62 75 65
rect 67 58 68 62
rect 72 58 75 62
rect 67 55 75 58
rect 77 82 85 94
rect 77 78 80 82
rect 84 78 85 82
rect 77 72 85 78
rect 77 68 80 72
rect 84 68 85 72
rect 77 62 85 68
rect 77 58 80 62
rect 84 58 85 62
rect 77 55 85 58
<< metal1 >>
rect -2 96 92 100
rect -2 92 28 96
rect 32 92 38 96
rect 42 92 48 96
rect 52 92 92 96
rect -2 88 16 92
rect 20 88 68 92
rect 72 88 92 92
rect 4 82 8 83
rect 4 72 8 78
rect 4 22 8 68
rect 18 62 22 83
rect 18 32 22 58
rect 18 27 22 28
rect 28 42 32 83
rect 28 27 32 38
rect 38 82 42 83
rect 38 72 42 78
rect 38 50 42 68
rect 58 62 62 83
rect 38 32 42 46
rect 38 27 42 28
rect 48 56 52 57
rect 48 22 52 52
rect 8 18 30 22
rect 34 18 52 22
rect 58 32 62 58
rect 68 82 72 88
rect 68 72 72 78
rect 68 62 72 68
rect 68 57 72 58
rect 78 82 82 83
rect 78 78 80 82
rect 84 78 85 82
rect 78 72 82 78
rect 78 68 80 72
rect 84 68 85 72
rect 78 62 82 68
rect 78 58 80 62
rect 84 58 85 62
rect 4 17 8 18
rect 58 17 62 28
rect 68 22 72 23
rect 68 12 72 18
rect 78 22 82 58
rect 78 18 80 22
rect 84 18 85 22
rect 78 17 82 18
rect -2 8 16 12
rect 20 8 68 12
rect 72 8 92 12
rect -2 0 92 8
<< ntransistor >>
rect 11 6 13 15
rect 23 6 25 14
rect 31 6 33 14
rect 47 6 49 15
rect 55 6 57 15
rect 75 6 77 25
<< ptransistor >>
rect 11 65 13 85
rect 23 66 25 85
rect 31 66 33 85
rect 47 66 49 85
rect 55 66 57 85
rect 75 55 77 94
<< polycontact >>
rect 18 58 22 62
rect 58 58 62 62
rect 48 52 52 56
rect 38 46 42 50
rect 28 38 32 42
rect 18 28 22 32
rect 30 18 34 22
rect 58 28 62 32
<< ndcontact >>
rect 4 18 8 22
rect 38 28 42 32
rect 68 18 72 22
rect 16 8 20 12
rect 68 8 72 12
rect 80 18 84 22
<< pdcontact >>
rect 16 88 20 92
rect 68 88 72 92
rect 4 78 8 82
rect 4 68 8 72
rect 38 78 42 82
rect 38 68 42 72
rect 68 78 72 82
rect 68 68 72 72
rect 68 58 72 62
rect 80 78 84 82
rect 80 68 84 72
rect 80 58 84 62
<< nsubstratencontact >>
rect 28 92 32 96
rect 38 92 42 96
rect 48 92 52 96
<< nsubstratendiff >>
rect 27 96 53 97
rect 27 92 28 96
rect 32 92 38 96
rect 42 92 48 96
rect 52 92 53 96
rect 27 91 53 92
<< labels >>
rlabel metal1 20 55 20 55 6 i0
rlabel metal1 30 55 30 55 6 cmd
rlabel metal1 45 6 45 6 6 vss
rlabel metal1 60 50 60 50 6 i1
rlabel metal1 45 94 45 94 6 vdd
rlabel metal1 80 50 80 50 6 q
<< end >>
