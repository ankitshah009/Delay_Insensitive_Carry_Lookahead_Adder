magic
tech scmos
timestamp 1179387511
<< checkpaint >>
rect -22 -25 158 105
<< ab >>
rect 0 0 136 80
<< pwell >>
rect -4 -7 140 36
<< nwell >>
rect -4 36 140 87
<< polysilicon >>
rect 18 70 20 74
rect 25 70 27 74
rect 35 70 37 74
rect 42 70 44 74
rect 52 70 54 74
rect 59 70 61 74
rect 73 70 75 74
rect 83 70 85 74
rect 93 70 95 74
rect 103 70 105 74
rect 115 70 117 74
rect 125 70 127 74
rect 18 22 20 42
rect 25 39 27 42
rect 35 39 37 42
rect 42 39 44 42
rect 52 39 54 42
rect 25 38 38 39
rect 25 37 33 38
rect 32 34 33 37
rect 37 34 38 38
rect 32 33 38 34
rect 42 37 54 39
rect 59 39 61 42
rect 73 39 75 42
rect 83 39 85 42
rect 93 39 95 42
rect 59 38 68 39
rect 59 37 63 38
rect 32 30 34 33
rect 42 30 44 37
rect 52 30 54 37
rect 62 34 63 37
rect 67 34 68 38
rect 62 33 68 34
rect 72 38 79 39
rect 72 34 74 38
rect 78 34 79 38
rect 83 38 99 39
rect 83 37 94 38
rect 72 33 79 34
rect 93 34 94 37
rect 98 34 99 38
rect 93 33 99 34
rect 62 30 64 33
rect 72 30 74 33
rect 103 30 105 42
rect 115 39 117 42
rect 125 39 127 42
rect 109 38 127 39
rect 109 34 110 38
rect 114 34 127 38
rect 109 33 127 34
rect 115 30 117 33
rect 125 30 127 33
rect 17 21 23 22
rect 17 17 18 21
rect 22 17 23 21
rect 17 16 23 17
rect 21 8 23 16
rect 32 12 34 16
rect 42 8 44 16
rect 52 11 54 16
rect 62 11 64 16
rect 21 6 44 8
rect 72 8 74 16
rect 103 8 105 16
rect 115 11 117 16
rect 125 11 127 16
rect 72 6 105 8
<< ndiffusion >>
rect 27 22 32 30
rect 25 21 32 22
rect 25 17 26 21
rect 30 17 32 21
rect 25 16 32 17
rect 34 29 42 30
rect 34 25 36 29
rect 40 25 42 29
rect 34 16 42 25
rect 44 29 52 30
rect 44 25 46 29
rect 50 25 52 29
rect 44 16 52 25
rect 54 29 62 30
rect 54 25 56 29
rect 60 25 62 29
rect 54 16 62 25
rect 64 22 72 30
rect 64 18 66 22
rect 70 18 72 22
rect 64 16 72 18
rect 74 16 82 30
rect 96 29 103 30
rect 96 25 97 29
rect 101 25 103 29
rect 96 22 103 25
rect 96 18 97 22
rect 101 18 103 22
rect 96 16 103 18
rect 105 28 115 30
rect 105 24 108 28
rect 112 24 115 28
rect 105 21 115 24
rect 105 17 108 21
rect 112 17 115 21
rect 105 16 115 17
rect 117 29 125 30
rect 117 25 119 29
rect 123 25 125 29
rect 117 22 125 25
rect 117 18 119 22
rect 123 18 125 22
rect 117 16 125 18
rect 127 28 134 30
rect 127 24 129 28
rect 133 24 134 28
rect 127 21 134 24
rect 127 17 129 21
rect 133 17 134 21
rect 127 16 134 17
rect 76 15 82 16
rect 76 11 77 15
rect 81 11 82 15
rect 76 10 82 11
<< pdiffusion >>
rect 13 55 18 70
rect 11 54 18 55
rect 11 50 12 54
rect 16 50 18 54
rect 11 47 18 50
rect 11 43 12 47
rect 16 43 18 47
rect 11 42 18 43
rect 20 42 25 70
rect 27 69 35 70
rect 27 65 29 69
rect 33 65 35 69
rect 27 42 35 65
rect 37 42 42 70
rect 44 62 52 70
rect 44 58 46 62
rect 50 58 52 62
rect 44 47 52 58
rect 44 43 46 47
rect 50 43 52 47
rect 44 42 52 43
rect 54 42 59 70
rect 61 69 73 70
rect 61 65 65 69
rect 69 65 73 69
rect 61 42 73 65
rect 75 47 83 70
rect 75 43 77 47
rect 81 43 83 47
rect 75 42 83 43
rect 85 62 93 70
rect 85 58 87 62
rect 91 58 93 62
rect 85 42 93 58
rect 95 47 103 70
rect 95 43 97 47
rect 101 43 103 47
rect 95 42 103 43
rect 105 69 115 70
rect 105 65 108 69
rect 112 65 115 69
rect 105 62 115 65
rect 105 58 108 62
rect 112 58 115 62
rect 105 42 115 58
rect 117 55 125 70
rect 117 51 119 55
rect 123 51 125 55
rect 117 47 125 51
rect 117 43 119 47
rect 123 43 125 47
rect 117 42 125 43
rect 127 69 134 70
rect 127 65 129 69
rect 133 65 134 69
rect 127 62 134 65
rect 127 58 129 62
rect 133 58 134 62
rect 127 42 134 58
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect 118 78 122 82
rect 126 78 130 82
rect 134 78 138 82
rect -2 69 138 78
rect -2 68 29 69
rect 28 65 29 68
rect 33 68 65 69
rect 33 65 34 68
rect 64 65 65 68
rect 69 68 108 69
rect 69 65 70 68
rect 107 65 108 68
rect 112 68 129 69
rect 112 65 113 68
rect 107 62 113 65
rect 26 58 46 62
rect 50 58 87 62
rect 91 58 92 62
rect 107 58 108 62
rect 112 58 113 62
rect 128 65 129 68
rect 133 68 138 69
rect 133 65 134 68
rect 128 62 134 65
rect 128 58 129 62
rect 133 58 134 62
rect 10 54 16 55
rect 10 50 12 54
rect 10 47 16 50
rect 10 43 12 47
rect 26 46 30 58
rect 119 55 123 56
rect 16 43 30 46
rect 10 42 30 43
rect 26 29 30 42
rect 37 51 119 54
rect 37 50 123 51
rect 37 39 41 50
rect 45 43 46 47
rect 50 46 51 47
rect 50 43 58 46
rect 45 42 58 43
rect 33 38 41 39
rect 37 37 41 38
rect 37 34 50 37
rect 33 33 50 34
rect 46 29 50 33
rect 26 25 36 29
rect 40 25 41 29
rect 54 29 58 42
rect 63 38 67 50
rect 119 47 123 50
rect 76 43 77 47
rect 81 46 82 47
rect 96 46 97 47
rect 81 43 97 46
rect 101 43 102 47
rect 76 42 102 43
rect 63 33 67 34
rect 73 34 74 38
rect 78 34 79 38
rect 73 30 79 34
rect 54 25 56 29
rect 60 25 61 29
rect 65 26 79 30
rect 83 26 87 42
rect 106 38 110 47
rect 93 34 94 38
rect 98 34 110 38
rect 114 34 115 38
rect 97 29 101 30
rect 119 29 123 43
rect 83 25 97 26
rect 46 24 50 25
rect 83 22 101 25
rect 65 21 66 22
rect 17 17 18 21
rect 22 17 26 21
rect 30 18 66 21
rect 70 18 87 22
rect 30 17 70 18
rect 97 17 101 18
rect 108 28 112 29
rect 108 21 112 24
rect 119 22 123 25
rect 119 17 123 18
rect 129 28 133 29
rect 129 21 133 24
rect 76 12 77 15
rect -2 11 77 12
rect 81 12 82 15
rect 86 12 92 15
rect 108 12 112 17
rect 129 12 133 17
rect 81 11 138 12
rect -2 2 138 11
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 122 2
rect 126 -2 130 2
rect 134 -2 138 2
<< ntransistor >>
rect 32 16 34 30
rect 42 16 44 30
rect 52 16 54 30
rect 62 16 64 30
rect 72 16 74 30
rect 103 16 105 30
rect 115 16 117 30
rect 125 16 127 30
<< ptransistor >>
rect 18 42 20 70
rect 25 42 27 70
rect 35 42 37 70
rect 42 42 44 70
rect 52 42 54 70
rect 59 42 61 70
rect 73 42 75 70
rect 83 42 85 70
rect 93 42 95 70
rect 103 42 105 70
rect 115 42 117 70
rect 125 42 127 70
<< polycontact >>
rect 33 34 37 38
rect 63 34 67 38
rect 74 34 78 38
rect 94 34 98 38
rect 110 34 114 38
rect 18 17 22 21
<< ndcontact >>
rect 26 17 30 21
rect 36 25 40 29
rect 46 25 50 29
rect 56 25 60 29
rect 66 18 70 22
rect 97 25 101 29
rect 97 18 101 22
rect 108 24 112 28
rect 108 17 112 21
rect 119 25 123 29
rect 119 18 123 22
rect 129 24 133 28
rect 129 17 133 21
rect 77 11 81 15
<< pdcontact >>
rect 12 50 16 54
rect 12 43 16 47
rect 29 65 33 69
rect 46 58 50 62
rect 46 43 50 47
rect 65 65 69 69
rect 77 43 81 47
rect 87 58 91 62
rect 97 43 101 47
rect 108 65 112 69
rect 108 58 112 62
rect 119 51 123 55
rect 119 43 123 47
rect 129 65 133 69
rect 129 58 133 62
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
rect 90 -2 94 2
rect 98 -2 102 2
rect 106 -2 110 2
rect 114 -2 118 2
rect 122 -2 126 2
rect 130 -2 134 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
rect 90 78 94 82
rect 98 78 102 82
rect 106 78 110 82
rect 114 78 118 82
rect 122 78 126 82
rect 130 78 134 82
<< psubstratepdiff >>
rect 0 2 136 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 122 2
rect 126 -2 130 2
rect 134 -2 136 2
rect 0 -3 136 -2
<< nsubstratendiff >>
rect 0 82 136 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect 118 78 122 82
rect 126 78 130 82
rect 134 78 136 82
rect 0 77 136 78
<< labels >>
rlabel ptransistor 19 45 19 45 6 an
rlabel ptransistor 36 53 36 53 6 bn
rlabel polycontact 65 36 65 36 6 bn
rlabel metal1 20 44 20 44 6 z
rlabel metal1 12 52 12 52 6 z
rlabel metal1 48 30 48 30 6 bn
rlabel metal1 28 40 28 40 6 z
rlabel metal1 39 43 39 43 6 bn
rlabel metal1 36 60 36 60 6 z
rlabel metal1 44 60 44 60 6 z
rlabel metal1 68 6 68 6 6 vss
rlabel metal1 43 19 43 19 6 an
rlabel metal1 68 28 68 28 6 a
rlabel metal1 76 32 76 32 6 a
rlabel metal1 65 43 65 43 6 bn
rlabel metal1 52 60 52 60 6 z
rlabel metal1 68 60 68 60 6 z
rlabel metal1 76 60 76 60 6 z
rlabel metal1 60 60 60 60 6 z
rlabel metal1 68 74 68 74 6 vdd
rlabel metal1 76 20 76 20 6 an
rlabel metal1 99 23 99 23 6 an
rlabel metal1 89 44 89 44 6 an
rlabel pdcontact 99 44 99 44 6 an
rlabel metal1 108 40 108 40 6 b
rlabel metal1 100 36 100 36 6 b
rlabel metal1 84 60 84 60 6 z
rlabel metal1 121 36 121 36 6 bn
<< end >>
