magic
tech scmos
timestamp 1179385068
<< checkpaint >>
rect -22 -22 78 94
<< ab >>
rect 0 0 56 72
<< pwell >>
rect -4 -4 60 32
<< nwell >>
rect -4 32 60 76
<< polysilicon >>
rect 9 58 11 63
rect 19 58 21 63
rect 29 58 31 63
rect 41 57 43 62
rect 9 35 11 40
rect 19 35 21 45
rect 29 42 31 45
rect 29 41 35 42
rect 29 37 30 41
rect 34 37 35 41
rect 29 36 35 37
rect 9 34 15 35
rect 9 30 10 34
rect 14 30 15 34
rect 9 29 15 30
rect 19 34 25 35
rect 19 30 20 34
rect 24 30 25 34
rect 19 29 25 30
rect 9 25 11 29
rect 22 25 24 29
rect 29 25 31 36
rect 41 35 43 44
rect 41 34 47 35
rect 41 31 42 34
rect 36 30 42 31
rect 46 30 47 34
rect 36 29 47 30
rect 36 25 38 29
rect 9 11 11 16
rect 22 7 24 12
rect 29 7 31 12
rect 36 7 38 12
<< ndiffusion >>
rect 2 24 9 25
rect 2 20 3 24
rect 7 20 9 24
rect 2 19 9 20
rect 4 16 9 19
rect 11 16 22 25
rect 13 12 22 16
rect 24 12 29 25
rect 31 12 36 25
rect 38 18 43 25
rect 38 17 45 18
rect 38 13 40 17
rect 44 13 45 17
rect 38 12 45 13
rect 13 8 20 12
rect 13 4 14 8
rect 18 4 20 8
rect 13 3 20 4
<< pdiffusion >>
rect 33 68 39 69
rect 33 64 34 68
rect 38 64 39 68
rect 33 58 39 64
rect 4 53 9 58
rect 2 52 9 53
rect 2 48 3 52
rect 7 48 9 52
rect 2 45 9 48
rect 2 41 3 45
rect 7 41 9 45
rect 2 40 9 41
rect 11 57 19 58
rect 11 53 13 57
rect 17 53 19 57
rect 11 45 19 53
rect 21 57 29 58
rect 21 53 23 57
rect 27 53 29 57
rect 21 50 29 53
rect 21 46 23 50
rect 27 46 29 50
rect 21 45 29 46
rect 31 57 39 58
rect 31 45 41 57
rect 11 40 17 45
rect 36 44 41 45
rect 43 56 50 57
rect 43 52 45 56
rect 49 52 50 56
rect 43 49 50 52
rect 43 45 45 49
rect 49 45 50 49
rect 43 44 50 45
<< metal1 >>
rect -2 68 58 72
rect -2 64 34 68
rect 38 64 48 68
rect 52 64 58 68
rect 2 52 7 59
rect 12 57 18 64
rect 12 53 13 57
rect 17 53 18 57
rect 23 57 50 58
rect 27 56 50 57
rect 27 54 45 56
rect 2 48 3 52
rect 23 50 27 53
rect 44 52 45 54
rect 49 52 50 56
rect 7 48 15 50
rect 2 46 15 48
rect 18 46 23 49
rect 2 45 7 46
rect 2 41 3 45
rect 18 45 27 46
rect 18 42 22 45
rect 33 42 39 50
rect 44 49 50 52
rect 44 45 45 49
rect 49 45 50 49
rect 2 40 7 41
rect 2 25 6 40
rect 10 38 22 42
rect 25 41 47 42
rect 25 38 30 41
rect 10 34 14 38
rect 29 37 30 38
rect 34 38 47 41
rect 34 37 35 38
rect 17 30 20 34
rect 24 30 30 34
rect 10 25 14 30
rect 2 24 7 25
rect 2 20 3 24
rect 10 21 19 25
rect 26 21 30 30
rect 41 30 42 34
rect 46 30 47 34
rect 41 27 47 30
rect 34 21 47 27
rect 2 19 7 20
rect 2 13 6 19
rect 15 17 19 21
rect 15 13 40 17
rect 44 13 45 17
rect -2 4 4 8
rect 8 4 14 8
rect 18 4 58 8
rect -2 0 58 4
<< ntransistor >>
rect 9 16 11 25
rect 22 12 24 25
rect 29 12 31 25
rect 36 12 38 25
<< ptransistor >>
rect 9 40 11 58
rect 19 45 21 58
rect 29 45 31 58
rect 41 44 43 57
<< polycontact >>
rect 30 37 34 41
rect 10 30 14 34
rect 20 30 24 34
rect 42 30 46 34
<< ndcontact >>
rect 3 20 7 24
rect 40 13 44 17
rect 14 4 18 8
<< pdcontact >>
rect 34 64 38 68
rect 3 48 7 52
rect 3 41 7 45
rect 13 53 17 57
rect 23 53 27 57
rect 23 46 27 50
rect 45 52 49 56
rect 45 45 49 49
<< psubstratepcontact >>
rect 4 4 8 8
<< nsubstratencontact >>
rect 48 64 52 68
<< psubstratepdiff >>
rect 3 8 9 9
rect 3 4 4 8
rect 8 4 9 8
rect 3 3 9 4
<< nsubstratendiff >>
rect 47 68 53 69
rect 47 64 48 68
rect 52 64 53 68
rect 47 63 53 64
<< labels >>
rlabel polycontact 12 32 12 32 6 zn
rlabel metal1 4 36 4 36 6 z
rlabel metal1 20 32 20 32 6 a
rlabel polycontact 12 31 12 31 6 zn
rlabel metal1 12 48 12 48 6 z
rlabel metal1 25 51 25 51 6 zn
rlabel metal1 28 4 28 4 6 vss
rlabel metal1 28 24 28 24 6 a
rlabel metal1 36 24 36 24 6 c
rlabel metal1 28 40 28 40 6 b
rlabel metal1 36 44 36 44 6 b
rlabel metal1 28 68 28 68 6 vdd
rlabel metal1 30 15 30 15 6 zn
rlabel metal1 44 28 44 28 6 c
rlabel polycontact 44 32 44 32 6 c
rlabel metal1 44 40 44 40 6 b
rlabel metal1 47 51 47 51 6 zn
<< end >>
