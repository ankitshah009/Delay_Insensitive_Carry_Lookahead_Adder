magic
tech scmos
timestamp 1179385485
<< checkpaint >>
rect -22 -22 62 94
<< ab >>
rect 0 0 40 72
<< pwell >>
rect -4 -4 44 32
<< nwell >>
rect -4 32 44 76
<< polysilicon >>
rect 9 66 11 70
rect 19 66 21 70
rect 29 65 31 70
rect 9 35 11 38
rect 19 35 21 38
rect 29 35 31 38
rect 9 34 22 35
rect 9 30 17 34
rect 21 30 22 34
rect 9 29 22 30
rect 26 34 32 35
rect 26 30 27 34
rect 31 30 32 34
rect 26 29 32 30
rect 9 26 11 29
rect 19 26 21 29
rect 29 26 31 29
rect 9 7 11 12
rect 19 7 21 12
rect 29 6 31 11
<< ndiffusion >>
rect 2 24 9 26
rect 2 20 3 24
rect 7 20 9 24
rect 2 17 9 20
rect 2 13 3 17
rect 7 13 9 17
rect 2 12 9 13
rect 11 18 19 26
rect 11 14 13 18
rect 17 14 19 18
rect 11 12 19 14
rect 21 17 29 26
rect 21 13 23 17
rect 27 13 29 17
rect 21 12 29 13
rect 23 11 29 12
rect 31 25 38 26
rect 31 21 33 25
rect 37 21 38 25
rect 31 18 38 21
rect 31 14 33 18
rect 37 14 38 18
rect 31 13 38 14
rect 31 11 36 13
<< pdiffusion >>
rect 2 65 9 66
rect 2 61 3 65
rect 7 61 9 65
rect 2 58 9 61
rect 2 54 3 58
rect 7 54 9 58
rect 2 38 9 54
rect 11 58 19 66
rect 11 54 13 58
rect 17 54 19 58
rect 11 51 19 54
rect 11 47 13 51
rect 17 47 19 51
rect 11 38 19 47
rect 21 65 27 66
rect 21 64 29 65
rect 21 60 23 64
rect 27 60 29 64
rect 21 57 29 60
rect 21 53 23 57
rect 27 53 29 57
rect 21 38 29 53
rect 31 58 36 65
rect 31 57 38 58
rect 31 53 33 57
rect 37 53 38 57
rect 31 50 38 53
rect 31 46 33 50
rect 37 46 38 50
rect 31 45 38 46
rect 31 38 36 45
<< metal1 >>
rect -2 65 42 72
rect -2 64 3 65
rect 2 61 3 64
rect 7 64 42 65
rect 7 61 8 64
rect 2 58 8 61
rect 2 54 3 58
rect 7 54 8 58
rect 13 58 17 59
rect 13 51 17 54
rect 23 57 27 60
rect 23 52 27 53
rect 33 57 38 58
rect 37 53 38 57
rect 2 47 13 50
rect 2 46 17 47
rect 33 50 38 53
rect 37 46 38 50
rect 2 33 6 46
rect 33 45 38 46
rect 17 38 31 42
rect 17 34 21 35
rect 2 29 14 33
rect 3 24 7 25
rect 3 17 7 20
rect 10 19 14 29
rect 17 26 21 30
rect 26 34 31 38
rect 26 30 27 34
rect 26 29 31 30
rect 34 26 38 45
rect 17 25 38 26
rect 17 22 33 25
rect 37 22 38 25
rect 10 18 17 19
rect 33 18 37 21
rect 10 14 13 18
rect 10 13 17 14
rect 23 17 27 18
rect 33 13 37 14
rect 3 8 7 13
rect 23 8 27 13
rect -2 0 42 8
<< ntransistor >>
rect 9 12 11 26
rect 19 12 21 26
rect 29 11 31 26
<< ptransistor >>
rect 9 38 11 66
rect 19 38 21 66
rect 29 38 31 65
<< polycontact >>
rect 17 30 21 34
rect 27 30 31 34
<< ndcontact >>
rect 3 20 7 24
rect 3 13 7 17
rect 13 14 17 18
rect 23 13 27 17
rect 33 21 37 25
rect 33 14 37 18
<< pdcontact >>
rect 3 61 7 65
rect 3 54 7 58
rect 13 54 17 58
rect 13 47 17 51
rect 23 60 27 64
rect 23 53 27 57
rect 33 53 37 57
rect 33 46 37 50
<< labels >>
rlabel polysilicon 15 32 15 32 6 an
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 20 12 20 6 z
rlabel metal1 12 48 12 48 6 z
rlabel metal1 20 4 20 4 6 vss
rlabel metal1 19 28 19 28 6 an
rlabel metal1 28 36 28 36 6 a
rlabel metal1 20 40 20 40 6 a
rlabel metal1 20 68 20 68 6 vdd
rlabel metal1 35 19 35 19 6 an
rlabel metal1 36 40 36 40 6 an
<< end >>
