magic
tech scmos
timestamp 1179386055
<< checkpaint >>
rect -22 -22 46 94
<< ab >>
rect 0 0 24 72
<< pwell >>
rect -4 -4 28 32
<< nwell >>
rect -4 32 28 76
<< polysilicon >>
rect 13 56 15 61
rect 13 35 15 41
rect 9 34 15 35
rect 9 30 10 34
rect 14 30 15 34
rect 9 29 15 30
rect 9 25 11 29
rect 9 13 11 18
<< ndiffusion >>
rect 2 24 9 25
rect 2 20 3 24
rect 7 20 9 24
rect 2 18 9 20
rect 11 18 19 25
rect 13 14 14 18
rect 18 14 19 18
rect 13 13 19 14
<< pdiffusion >>
rect 5 58 11 59
rect 5 54 6 58
rect 10 56 11 58
rect 10 54 13 56
rect 5 41 13 54
rect 15 51 20 56
rect 15 50 22 51
rect 15 46 17 50
rect 21 46 22 50
rect 15 45 22 46
rect 15 41 20 45
<< metal1 >>
rect -2 68 26 72
rect -2 64 4 68
rect 8 64 16 68
rect 20 64 26 68
rect 5 58 11 64
rect 5 54 6 58
rect 10 54 11 58
rect 2 46 17 50
rect 21 46 22 50
rect 2 25 6 46
rect 10 34 22 35
rect 14 30 22 34
rect 10 29 22 30
rect 2 24 7 25
rect 2 20 3 24
rect 18 21 22 29
rect 2 19 7 20
rect 13 14 14 18
rect 18 14 19 18
rect 13 8 19 14
rect -2 4 4 8
rect 8 4 16 8
rect 20 4 26 8
rect -2 0 26 4
<< ntransistor >>
rect 9 18 11 25
<< ptransistor >>
rect 13 41 15 56
<< polycontact >>
rect 10 30 14 34
<< ndcontact >>
rect 3 20 7 24
rect 14 14 18 18
<< pdcontact >>
rect 6 54 10 58
rect 17 46 21 50
<< psubstratepcontact >>
rect 4 4 8 8
rect 16 4 20 8
<< nsubstratencontact >>
rect 4 64 8 68
rect 16 64 20 68
<< psubstratepdiff >>
rect 3 8 21 9
rect 3 4 4 8
rect 8 4 16 8
rect 20 4 21 8
rect 3 3 21 4
<< nsubstratendiff >>
rect 3 68 21 69
rect 3 64 4 68
rect 8 64 16 68
rect 20 64 21 68
rect 3 63 21 64
<< labels >>
rlabel metal1 4 32 4 32 6 z
rlabel metal1 12 4 12 4 6 vss
rlabel polycontact 12 32 12 32 6 a
rlabel metal1 12 48 12 48 6 z
rlabel metal1 12 68 12 68 6 vdd
rlabel metal1 20 28 20 28 6 a
<< end >>
