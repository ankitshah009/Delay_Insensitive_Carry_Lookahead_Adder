magic
tech scmos
timestamp 1179387023
<< checkpaint >>
rect -22 -22 86 94
<< ab >>
rect 0 0 64 72
<< pwell >>
rect -4 -4 68 32
<< nwell >>
rect -4 32 68 76
<< polysilicon >>
rect 10 66 12 70
rect 22 66 24 70
rect 29 66 31 70
rect 39 66 41 70
rect 46 66 48 70
rect 10 35 12 38
rect 22 35 24 38
rect 29 35 31 38
rect 39 35 41 38
rect 9 34 15 35
rect 9 30 10 34
rect 14 30 15 34
rect 9 29 15 30
rect 19 34 25 35
rect 19 30 20 34
rect 24 30 25 34
rect 19 29 25 30
rect 29 34 41 35
rect 29 30 34 34
rect 38 30 41 34
rect 29 29 41 30
rect 46 35 48 38
rect 46 34 55 35
rect 46 30 50 34
rect 54 30 55 34
rect 46 29 55 30
rect 9 26 11 29
rect 30 26 32 29
rect 46 26 48 29
rect 20 20 22 25
rect 9 5 11 8
rect 20 5 22 8
rect 9 3 22 5
rect 30 2 32 6
rect 46 2 48 6
<< ndiffusion >>
rect 4 19 9 26
rect 2 18 9 19
rect 2 14 3 18
rect 7 14 9 18
rect 2 13 9 14
rect 4 8 9 13
rect 11 25 18 26
rect 11 21 13 25
rect 17 21 18 25
rect 11 20 18 21
rect 25 20 30 26
rect 11 8 20 20
rect 22 18 30 20
rect 22 14 24 18
rect 28 14 30 18
rect 22 8 30 14
rect 25 6 30 8
rect 32 11 46 26
rect 32 7 37 11
rect 41 7 46 11
rect 32 6 46 7
rect 48 19 53 26
rect 48 18 55 19
rect 48 14 50 18
rect 54 14 55 18
rect 48 13 55 14
rect 48 6 53 13
<< pdiffusion >>
rect 5 59 10 66
rect 2 58 10 59
rect 2 54 3 58
rect 7 54 10 58
rect 2 51 10 54
rect 2 47 3 51
rect 7 47 10 51
rect 2 46 10 47
rect 5 38 10 46
rect 12 65 22 66
rect 12 61 15 65
rect 19 61 22 65
rect 12 38 22 61
rect 24 38 29 66
rect 31 58 39 66
rect 31 54 33 58
rect 37 54 39 58
rect 31 51 39 54
rect 31 47 33 51
rect 37 47 39 51
rect 31 38 39 47
rect 41 38 46 66
rect 48 65 57 66
rect 48 61 51 65
rect 55 61 57 65
rect 48 58 57 61
rect 48 54 51 58
rect 55 54 57 58
rect 48 38 57 54
<< metal1 >>
rect -2 65 66 72
rect -2 64 15 65
rect 14 61 15 64
rect 19 64 51 65
rect 19 61 20 64
rect 50 61 51 64
rect 55 64 66 65
rect 55 61 56 64
rect 50 58 56 61
rect 2 54 3 58
rect 7 54 33 58
rect 37 54 38 58
rect 50 54 51 58
rect 55 54 56 58
rect 2 51 7 54
rect 2 47 3 51
rect 33 51 38 54
rect 2 46 7 47
rect 2 25 6 46
rect 17 43 23 50
rect 37 47 38 51
rect 33 46 38 47
rect 10 38 23 43
rect 42 42 46 51
rect 10 34 14 38
rect 33 37 46 42
rect 33 34 39 37
rect 19 30 20 34
rect 24 30 27 34
rect 33 30 34 34
rect 38 30 39 34
rect 50 34 55 43
rect 54 30 55 34
rect 10 29 14 30
rect 23 26 27 30
rect 50 26 55 30
rect 2 21 13 25
rect 17 21 18 25
rect 23 22 55 26
rect 2 14 3 18
rect 7 14 24 18
rect 28 14 50 18
rect 54 14 55 18
rect 36 8 37 11
rect -2 7 37 8
rect 41 8 42 11
rect 41 7 66 8
rect -2 0 66 7
<< ntransistor >>
rect 9 8 11 26
rect 20 8 22 20
rect 30 6 32 26
rect 46 6 48 26
<< ptransistor >>
rect 10 38 12 66
rect 22 38 24 66
rect 29 38 31 66
rect 39 38 41 66
rect 46 38 48 66
<< polycontact >>
rect 10 30 14 34
rect 20 30 24 34
rect 34 30 38 34
rect 50 30 54 34
<< ndcontact >>
rect 3 14 7 18
rect 13 21 17 25
rect 24 14 28 18
rect 37 7 41 11
rect 50 14 54 18
<< pdcontact >>
rect 3 54 7 58
rect 3 47 7 51
rect 15 61 19 65
rect 33 54 37 58
rect 33 47 37 51
rect 51 61 55 65
rect 51 54 55 58
<< labels >>
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 36 12 36 6 b
rlabel metal1 12 56 12 56 6 z
rlabel metal1 28 24 28 24 6 a1
rlabel metal1 20 44 20 44 6 b
rlabel metal1 20 56 20 56 6 z
rlabel metal1 28 56 28 56 6 z
rlabel metal1 32 4 32 4 6 vss
rlabel metal1 36 24 36 24 6 a1
rlabel metal1 44 24 44 24 6 a1
rlabel metal1 36 36 36 36 6 a2
rlabel metal1 44 44 44 44 6 a2
rlabel metal1 32 68 32 68 6 vdd
rlabel metal1 28 16 28 16 6 n1
rlabel polycontact 52 32 52 32 6 a1
<< end >>
