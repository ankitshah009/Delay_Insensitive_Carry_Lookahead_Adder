magic
tech scmos
timestamp 1185094765
<< checkpaint >>
rect -22 -22 62 122
<< ab >>
rect 0 0 40 100
<< pwell >>
rect -4 -4 44 48
<< nwell >>
rect -4 48 44 104
<< polysilicon >>
rect 15 78 17 83
rect 23 78 25 83
rect 15 43 17 56
rect 23 53 25 56
rect 23 52 29 53
rect 23 48 24 52
rect 28 48 29 52
rect 23 47 29 48
rect 13 42 21 43
rect 13 38 16 42
rect 20 38 21 42
rect 13 37 21 38
rect 13 23 15 37
rect 25 23 27 47
rect 13 12 15 17
rect 25 12 27 17
<< ndiffusion >>
rect 5 22 13 23
rect 5 18 6 22
rect 10 18 13 22
rect 5 17 13 18
rect 15 22 25 23
rect 15 18 18 22
rect 22 18 25 22
rect 15 17 25 18
rect 27 22 35 23
rect 27 18 30 22
rect 34 18 35 22
rect 27 17 35 18
<< pdiffusion >>
rect 10 70 15 78
rect 7 69 15 70
rect 7 65 8 69
rect 12 65 15 69
rect 7 61 15 65
rect 7 57 8 61
rect 12 57 15 61
rect 7 56 15 57
rect 17 56 23 78
rect 25 72 34 78
rect 25 68 28 72
rect 32 68 34 72
rect 25 62 34 68
rect 25 58 28 62
rect 32 58 34 62
rect 25 56 34 58
<< metal1 >>
rect -2 96 42 100
rect -2 92 8 96
rect 12 92 18 96
rect 22 92 42 96
rect -2 88 42 92
rect 28 72 32 88
rect 8 69 12 70
rect 8 61 12 65
rect 8 33 12 57
rect 18 53 22 63
rect 28 62 32 68
rect 28 57 32 58
rect 18 52 32 53
rect 18 48 24 52
rect 28 48 32 52
rect 18 47 32 48
rect 16 42 32 43
rect 20 38 32 42
rect 16 37 32 38
rect 8 27 22 33
rect 28 27 32 37
rect 6 22 10 23
rect 6 12 10 18
rect 18 22 22 27
rect 18 17 22 18
rect 30 22 34 23
rect 30 12 34 18
rect -2 8 42 12
rect -2 4 8 8
rect 12 4 18 8
rect 22 4 42 8
rect -2 0 42 4
<< ntransistor >>
rect 13 17 15 23
rect 25 17 27 23
<< ptransistor >>
rect 15 56 17 78
rect 23 56 25 78
<< polycontact >>
rect 24 48 28 52
rect 16 38 20 42
<< ndcontact >>
rect 6 18 10 22
rect 18 18 22 22
rect 30 18 34 22
<< pdcontact >>
rect 8 65 12 69
rect 8 57 12 61
rect 28 68 32 72
rect 28 58 32 62
<< psubstratepcontact >>
rect 8 4 12 8
rect 18 4 22 8
<< nsubstratencontact >>
rect 8 92 12 96
rect 18 92 22 96
<< psubstratepdiff >>
rect 7 8 23 9
rect 7 4 8 8
rect 12 4 18 8
rect 22 4 23 8
rect 7 3 23 4
<< nsubstratendiff >>
rect 7 96 23 97
rect 7 92 8 96
rect 12 92 18 96
rect 22 92 23 96
rect 7 91 23 92
<< labels >>
rlabel metal1 10 45 10 45 6 z
rlabel psubstratepcontact 20 6 20 6 6 vss
rlabel metal1 20 25 20 25 6 z
rlabel metal1 20 40 20 40 6 b
rlabel metal1 20 55 20 55 6 a
rlabel nsubstratencontact 20 94 20 94 6 vdd
rlabel metal1 30 35 30 35 6 b
rlabel metal1 30 50 30 50 6 a
<< end >>
