.subckt nr2a_x1 a b vdd vss z
*   SPICE3 file   created from nr2a_x1.ext -      technology: scmos
m00 w1     b      z      vdd p w=39u  l=2.3636u ad=117p     pd=45u      as=237p     ps=94u
m01 vdd    an     w1     vdd p w=39u  l=2.3636u ad=277.475p pd=65.2131u as=117p     ps=45u
m02 an     a      vdd    vdd p w=22u  l=2.3636u ad=152p     pd=60u      as=156.525p ps=36.7869u
m03 z      b      vss    vss n w=11u  l=2.3636u ad=55p      pd=21u      as=93p      ps=34u
m04 vss    an     z      vss n w=11u  l=2.3636u ad=93p      pd=34u      as=55p      ps=21u
m05 an     a      vss    vss n w=11u  l=2.3636u ad=73p      pd=38u      as=93p      ps=34u
C0  vss    b      0.062f
C1  w1     vdd    0.011f
C2  a      an     0.214f
C3  z      an     0.053f
C4  vdd    b      0.012f
C5  vss    a      0.014f
C6  vss    z      0.134f
C7  a      w1     0.035f
C8  vss    an     0.043f
C9  a      vdd    0.103f
C10 a      b      0.106f
C11 z      vdd    0.029f
C12 z      b      0.193f
C13 vdd    an     0.024f
C14 an     b      0.209f
C15 a      z      0.103f
C17 a      vss    0.026f
C18 z      vss    0.014f
C20 an     vss    0.040f
C21 b      vss    0.037f
.ends
