magic
tech scmos
timestamp 1185094644
<< checkpaint >>
rect -22 -22 82 122
<< ab >>
rect 0 0 60 100
<< pwell >>
rect -4 -4 64 48
<< nwell >>
rect -4 48 64 104
<< polysilicon >>
rect 11 94 13 98
rect 23 94 25 98
rect 35 94 37 98
rect 47 94 49 98
rect 11 43 13 55
rect 23 52 25 55
rect 35 52 37 55
rect 23 49 27 52
rect 35 51 43 52
rect 35 49 38 51
rect 25 43 27 49
rect 37 47 38 49
rect 42 47 43 51
rect 37 46 43 47
rect 11 42 21 43
rect 11 41 16 42
rect 15 38 16 41
rect 20 38 21 42
rect 15 37 21 38
rect 25 42 33 43
rect 25 38 28 42
rect 32 38 33 42
rect 25 37 33 38
rect 17 34 19 37
rect 25 34 27 37
rect 37 34 39 46
rect 47 43 49 55
rect 47 42 53 43
rect 47 40 48 42
rect 45 38 48 40
rect 52 38 53 42
rect 45 37 53 38
rect 45 34 47 37
rect 17 12 19 17
rect 25 12 27 17
rect 37 12 39 17
rect 45 12 47 17
<< ndiffusion >>
rect 9 17 17 34
rect 19 17 25 34
rect 27 22 37 34
rect 27 18 30 22
rect 34 18 37 22
rect 27 17 37 18
rect 39 17 45 34
rect 47 22 56 34
rect 47 18 50 22
rect 54 18 56 22
rect 47 17 56 18
rect 9 12 15 17
rect 9 8 10 12
rect 14 8 15 12
rect 9 7 15 8
<< pdiffusion >>
rect 6 83 11 94
rect 3 82 11 83
rect 3 78 4 82
rect 8 78 11 82
rect 3 77 11 78
rect 6 55 11 77
rect 13 72 23 94
rect 13 68 16 72
rect 20 68 23 72
rect 13 55 23 68
rect 25 82 35 94
rect 25 78 28 82
rect 32 78 35 82
rect 25 72 35 78
rect 25 68 28 72
rect 32 68 35 72
rect 25 55 35 68
rect 37 92 47 94
rect 37 88 40 92
rect 44 88 47 92
rect 37 82 47 88
rect 37 78 40 82
rect 44 78 47 82
rect 37 55 47 78
rect 49 83 54 94
rect 49 82 57 83
rect 49 78 52 82
rect 56 78 57 82
rect 49 74 57 78
rect 49 70 52 74
rect 56 70 57 74
rect 49 69 57 70
rect 49 55 54 69
<< metal1 >>
rect -2 92 62 100
rect -2 88 40 92
rect 44 88 62 92
rect 40 82 44 88
rect 3 78 4 82
rect 8 78 28 82
rect 32 78 33 82
rect 8 72 23 73
rect 8 68 16 72
rect 20 68 23 72
rect 27 72 33 78
rect 40 77 44 78
rect 52 82 56 83
rect 52 74 56 78
rect 27 68 28 72
rect 32 70 52 72
rect 32 68 56 70
rect 8 22 12 68
rect 17 58 32 63
rect 18 43 22 53
rect 16 42 22 43
rect 20 38 22 42
rect 16 37 22 38
rect 28 42 32 58
rect 28 37 32 38
rect 38 58 53 63
rect 38 51 42 58
rect 38 37 42 47
rect 48 42 52 53
rect 18 32 22 37
rect 48 32 52 38
rect 18 27 33 32
rect 37 27 52 32
rect 50 22 54 23
rect 8 18 30 22
rect 34 18 35 22
rect 8 17 35 18
rect 50 12 54 18
rect -2 8 10 12
rect 14 8 62 12
rect -2 4 38 8
rect 42 4 48 8
rect 52 4 62 8
rect -2 0 62 4
<< ntransistor >>
rect 17 17 19 34
rect 25 17 27 34
rect 37 17 39 34
rect 45 17 47 34
<< ptransistor >>
rect 11 55 13 94
rect 23 55 25 94
rect 35 55 37 94
rect 47 55 49 94
<< polycontact >>
rect 38 47 42 51
rect 16 38 20 42
rect 28 38 32 42
rect 48 38 52 42
<< ndcontact >>
rect 30 18 34 22
rect 50 18 54 22
rect 10 8 14 12
<< pdcontact >>
rect 4 78 8 82
rect 16 68 20 72
rect 28 78 32 82
rect 28 68 32 72
rect 40 88 44 92
rect 40 78 44 82
rect 52 78 56 82
rect 52 70 56 74
<< psubstratepcontact >>
rect 38 4 42 8
rect 48 4 52 8
<< psubstratepdiff >>
rect 37 8 53 9
rect 37 4 38 8
rect 42 4 48 8
rect 52 4 53 8
rect 37 3 53 4
<< labels >>
rlabel metal1 20 20 20 20 6 z
rlabel metal1 20 40 20 40 6 b1
rlabel metal1 10 45 10 45 6 z
rlabel metal1 20 60 20 60 6 b2
rlabel metal1 20 70 20 70 6 z
rlabel metal1 30 6 30 6 6 vss
rlabel metal1 30 20 30 20 6 z
rlabel metal1 30 30 30 30 6 b1
rlabel metal1 30 50 30 50 6 b2
rlabel metal1 30 75 30 75 6 n3
rlabel metal1 18 80 18 80 6 n3
rlabel metal1 30 94 30 94 6 vdd
rlabel metal1 40 30 40 30 6 a1
rlabel polycontact 40 50 40 50 6 a2
rlabel polycontact 50 40 50 40 6 a1
rlabel metal1 50 60 50 60 6 a2
rlabel metal1 54 75 54 75 6 n3
<< end >>
