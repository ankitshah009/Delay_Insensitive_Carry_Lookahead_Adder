magic
tech scmos
timestamp 1179385114
<< checkpaint >>
rect -22 -22 78 94
<< ab >>
rect 0 0 56 72
<< pwell >>
rect -4 -4 60 32
<< nwell >>
rect -4 32 60 76
<< polysilicon >>
rect 9 60 11 65
rect 19 60 21 65
rect 29 60 31 65
rect 41 59 47 60
rect 41 55 42 59
rect 46 55 47 59
rect 41 54 47 55
rect 41 51 43 54
rect 9 27 11 49
rect 19 43 21 49
rect 15 42 21 43
rect 15 38 16 42
rect 20 38 21 42
rect 15 37 21 38
rect 8 26 14 27
rect 8 22 9 26
rect 13 22 14 26
rect 8 21 14 22
rect 12 18 14 21
rect 19 18 21 37
rect 29 27 31 49
rect 25 26 31 27
rect 41 26 43 39
rect 25 22 26 26
rect 30 22 31 26
rect 25 21 31 22
rect 26 18 28 21
rect 41 17 43 20
rect 41 16 47 17
rect 41 12 42 16
rect 46 12 47 16
rect 41 11 47 12
rect 12 2 14 7
rect 19 2 21 7
rect 26 2 28 7
<< ndiffusion >>
rect 33 20 41 26
rect 43 25 50 26
rect 43 21 45 25
rect 49 21 50 25
rect 43 20 50 21
rect 33 18 39 20
rect 5 17 12 18
rect 5 13 6 17
rect 10 13 12 17
rect 5 12 12 13
rect 7 7 12 12
rect 14 7 19 18
rect 21 7 26 18
rect 28 8 39 18
rect 28 7 33 8
rect 30 4 33 7
rect 37 4 39 8
rect 30 3 39 4
<< pdiffusion >>
rect 33 68 39 69
rect 33 64 34 68
rect 38 64 39 68
rect 33 60 39 64
rect 4 55 9 60
rect 2 54 9 55
rect 2 50 3 54
rect 7 50 9 54
rect 2 49 9 50
rect 11 59 19 60
rect 11 55 13 59
rect 17 55 19 59
rect 11 49 19 55
rect 21 56 29 60
rect 21 52 23 56
rect 27 52 29 56
rect 21 49 29 52
rect 31 51 39 60
rect 31 49 41 51
rect 33 39 41 49
rect 43 45 48 51
rect 43 44 50 45
rect 43 40 45 44
rect 49 40 50 44
rect 43 39 50 40
<< metal1 >>
rect -2 68 58 72
rect -2 64 34 68
rect 38 64 44 68
rect 48 64 58 68
rect 12 59 18 64
rect 12 55 13 59
rect 17 55 18 59
rect 23 56 42 59
rect 3 54 7 55
rect 27 55 42 56
rect 46 55 47 59
rect 23 51 27 52
rect 7 50 27 51
rect 3 47 27 50
rect 34 45 46 51
rect 42 44 49 45
rect 2 27 6 43
rect 10 42 30 43
rect 10 38 16 42
rect 20 38 30 42
rect 10 37 30 38
rect 42 40 45 44
rect 42 39 49 40
rect 18 29 22 37
rect 34 27 38 35
rect 2 26 14 27
rect 2 22 9 26
rect 13 22 14 26
rect 2 21 14 22
rect 26 26 38 27
rect 30 22 38 26
rect 26 21 38 22
rect 42 25 46 39
rect 42 21 45 25
rect 49 21 50 25
rect 5 13 6 17
rect 10 16 47 17
rect 10 13 42 16
rect 41 12 42 13
rect 46 12 47 16
rect -2 4 33 8
rect 37 4 44 8
rect 48 4 58 8
rect -2 0 58 4
<< ntransistor >>
rect 41 20 43 26
rect 12 7 14 18
rect 19 7 21 18
rect 26 7 28 18
<< ptransistor >>
rect 9 49 11 60
rect 19 49 21 60
rect 29 49 31 60
rect 41 39 43 51
<< polycontact >>
rect 42 55 46 59
rect 16 38 20 42
rect 9 22 13 26
rect 26 22 30 26
rect 42 12 46 16
<< ndcontact >>
rect 45 21 49 25
rect 6 13 10 17
rect 33 4 37 8
<< pdcontact >>
rect 34 64 38 68
rect 3 50 7 54
rect 13 55 17 59
rect 23 52 27 56
rect 45 40 49 44
<< psubstratepcontact >>
rect 44 4 48 8
<< nsubstratencontact >>
rect 44 64 48 68
<< psubstratepdiff >>
rect 43 8 49 9
rect 43 4 44 8
rect 48 4 49 8
rect 43 3 49 4
<< nsubstratendiff >>
rect 43 68 49 69
rect 43 64 44 68
rect 48 64 49 68
rect 43 63 49 64
<< labels >>
rlabel polycontact 44 14 44 14 6 zn
rlabel polycontact 44 57 44 57 6 zn
rlabel metal1 4 32 4 32 6 c
rlabel polycontact 12 24 12 24 6 c
rlabel metal1 20 36 20 36 6 b
rlabel metal1 12 40 12 40 6 b
rlabel metal1 15 49 15 49 6 zn
rlabel pdcontact 25 53 25 53 6 zn
rlabel metal1 28 4 28 4 6 vss
rlabel polycontact 28 24 28 24 6 a
rlabel metal1 36 28 36 28 6 a
rlabel metal1 28 40 28 40 6 b
rlabel metal1 36 48 36 48 6 z
rlabel metal1 28 68 28 68 6 vdd
rlabel polycontact 44 14 44 14 6 zn
rlabel metal1 26 15 26 15 6 zn
rlabel metal1 44 36 44 36 6 z
rlabel metal1 35 57 35 57 6 zn
<< end >>
