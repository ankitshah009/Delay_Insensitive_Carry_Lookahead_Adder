magic
tech scmos
timestamp 1179386505
<< checkpaint >>
rect -22 -25 78 105
<< ab >>
rect 0 0 56 80
<< pwell >>
rect -4 -7 60 36
<< nwell >>
rect -4 36 60 87
<< polysilicon >>
rect 9 63 11 69
rect 19 63 21 69
rect 31 61 33 65
rect 41 61 43 65
rect 9 39 11 44
rect 19 41 21 44
rect 31 41 33 44
rect 19 40 33 41
rect 9 38 15 39
rect 9 34 10 38
rect 14 34 15 38
rect 9 33 15 34
rect 19 36 26 40
rect 30 39 33 40
rect 41 39 43 44
rect 30 36 31 39
rect 19 35 31 36
rect 41 38 47 39
rect 41 35 42 38
rect 12 30 14 33
rect 19 30 21 35
rect 29 30 31 35
rect 36 34 42 35
rect 46 34 47 38
rect 36 33 47 34
rect 36 30 38 33
rect 12 8 14 13
rect 19 8 21 13
rect 29 12 31 17
rect 36 12 38 17
<< ndiffusion >>
rect 3 13 12 30
rect 14 13 19 30
rect 21 22 29 30
rect 21 18 23 22
rect 27 18 29 22
rect 21 17 29 18
rect 31 17 36 30
rect 38 22 46 30
rect 38 18 40 22
rect 44 18 46 22
rect 38 17 46 18
rect 21 13 26 17
rect 3 12 10 13
rect 3 8 5 12
rect 9 8 10 12
rect 3 7 10 8
<< pdiffusion >>
rect 2 62 9 63
rect 2 58 3 62
rect 7 58 9 62
rect 2 55 9 58
rect 2 51 3 55
rect 7 51 9 55
rect 2 44 9 51
rect 11 56 19 63
rect 11 52 13 56
rect 17 52 19 56
rect 11 49 19 52
rect 11 45 13 49
rect 17 45 19 49
rect 11 44 19 45
rect 21 62 29 63
rect 21 58 24 62
rect 28 61 29 62
rect 28 58 31 61
rect 21 44 31 58
rect 33 60 41 61
rect 33 56 35 60
rect 39 56 41 60
rect 33 53 41 56
rect 33 49 35 53
rect 39 49 41 53
rect 33 44 41 49
rect 43 60 50 61
rect 43 56 45 60
rect 49 56 50 60
rect 43 53 50 56
rect 43 49 45 53
rect 49 49 50 53
rect 43 44 50 49
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect -2 68 58 78
rect 2 62 8 68
rect 2 58 3 62
rect 7 58 8 62
rect 23 62 29 68
rect 23 58 24 62
rect 28 58 29 62
rect 34 60 40 63
rect 2 55 8 58
rect 2 51 3 55
rect 7 51 8 55
rect 13 56 17 58
rect 34 56 35 60
rect 39 56 40 60
rect 34 54 40 56
rect 17 53 40 54
rect 17 52 35 53
rect 13 50 35 52
rect 13 49 17 50
rect 34 49 35 50
rect 39 49 40 53
rect 44 60 50 68
rect 44 56 45 60
rect 49 56 50 60
rect 44 53 50 56
rect 44 49 45 53
rect 49 49 50 53
rect 2 45 13 47
rect 2 43 17 45
rect 2 22 6 43
rect 25 42 39 46
rect 25 40 31 42
rect 10 38 18 39
rect 14 34 18 38
rect 25 36 26 40
rect 30 36 31 40
rect 25 34 31 36
rect 41 34 42 38
rect 46 34 47 38
rect 10 33 18 34
rect 14 30 18 33
rect 41 30 47 34
rect 14 26 47 30
rect 2 18 23 22
rect 27 18 31 22
rect 39 18 40 22
rect 44 18 45 22
rect 39 12 45 18
rect -2 8 5 12
rect 9 8 58 12
rect -2 2 58 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
<< ntransistor >>
rect 12 13 14 30
rect 19 13 21 30
rect 29 17 31 30
rect 36 17 38 30
<< ptransistor >>
rect 9 44 11 63
rect 19 44 21 63
rect 31 44 33 61
rect 41 44 43 61
<< polycontact >>
rect 10 34 14 38
rect 26 36 30 40
rect 42 34 46 38
<< ndcontact >>
rect 23 18 27 22
rect 40 18 44 22
rect 5 8 9 12
<< pdcontact >>
rect 3 58 7 62
rect 3 51 7 55
rect 13 52 17 56
rect 13 45 17 49
rect 24 58 28 62
rect 35 56 39 60
rect 35 49 39 53
rect 45 56 49 60
rect 45 49 49 53
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
<< psubstratepdiff >>
rect 0 2 56 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 56 2
rect 0 -3 56 -2
<< nsubstratendiff >>
rect 0 82 56 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 56 82
rect 0 77 56 78
<< labels >>
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 20 12 20 6 z
rlabel polycontact 12 36 12 36 6 a
rlabel metal1 28 6 28 6 6 vss
rlabel metal1 20 20 20 20 6 z
rlabel metal1 20 28 20 28 6 a
rlabel metal1 28 28 28 28 6 a
rlabel metal1 28 20 28 20 6 z
rlabel metal1 28 40 28 40 6 b
rlabel metal1 28 52 28 52 6 z
rlabel metal1 20 52 20 52 6 z
rlabel metal1 28 74 28 74 6 vdd
rlabel metal1 36 28 36 28 6 a
rlabel metal1 44 32 44 32 6 a
rlabel metal1 36 44 36 44 6 b
rlabel metal1 36 56 36 56 6 z
<< end >>
