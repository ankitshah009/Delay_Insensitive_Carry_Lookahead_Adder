.subckt xor2v0x05 a b vdd vss z
*   SPICE3 file   created from xor2v0x05.ext -      technology: scmos
m00 vdd    b      bn     vdd p w=21u  l=2.3636u ad=145.765p pd=40.7647u as=124p     ps=56u
m01 an     a      vdd    vdd p w=13u  l=2.3636u ad=52p      pd=21u      as=90.2353p ps=25.2353u
m02 z      bn     an     vdd p w=13u  l=2.3636u ad=55.0588p pd=22.1765u as=52p      ps=21u
m03 bn     an     z      vdd p w=21u  l=2.3636u ad=124p     pd=56u      as=88.9412p ps=35.8235u
m04 vss    b      bn     vss n w=7u   l=2.3636u ad=55.3913p pd=24.3478u as=49p      ps=28u
m05 an     a      vss    vss n w=7u   l=2.3636u ad=28p      pd=15u      as=55.3913p ps=24.3478u
m06 z      b      an     vss n w=7u   l=2.3636u ad=28.875p  pd=14.875u  as=28p      ps=15u
m07 w1     bn     z      vss n w=9u   l=2.3636u ad=22.5p    pd=14u      as=37.125p  ps=19.125u
m08 vss    an     w1     vss n w=9u   l=2.3636u ad=71.2174p pd=31.3043u as=22.5p    ps=14u
C0  bn     vdd    0.314f
C1  vss    z      0.148f
C2  vss    an     0.088f
C3  z      a      0.013f
C4  a      an     0.075f
C5  vss    b      0.016f
C6  z      bn     0.164f
C7  a      b      0.071f
C8  z      vdd    0.032f
C9  an     bn     0.165f
C10 an     vdd    0.028f
C11 bn     b      0.114f
C12 w1     z      0.011f
C13 b      vdd    0.113f
C14 vss    a      0.069f
C15 z      an     0.287f
C16 vss    bn     0.040f
C17 z      b      0.004f
C18 a      bn     0.142f
C19 a      vdd    0.017f
C20 an     b      0.026f
C22 z      vss    0.013f
C23 a      vss    0.024f
C24 an     vss    0.032f
C25 bn     vss    0.034f
C26 b      vss    0.052f
.ends
