magic
tech scmos
timestamp 1179385456
<< checkpaint >>
rect -22 -22 126 94
<< ab >>
rect 0 0 104 72
<< pwell >>
rect -4 -4 108 32
<< nwell >>
rect -4 32 108 76
<< polysilicon >>
rect 9 66 11 70
rect 19 66 21 70
rect 29 66 31 70
rect 39 66 41 70
rect 49 66 51 70
rect 59 61 61 66
rect 69 57 71 61
rect 79 57 81 61
rect 89 57 91 61
rect 9 35 11 38
rect 19 35 21 38
rect 29 35 31 38
rect 39 35 41 38
rect 9 34 41 35
rect 9 33 36 34
rect 29 30 36 33
rect 40 30 41 34
rect 29 29 41 30
rect 29 26 31 29
rect 39 26 41 29
rect 49 35 51 38
rect 59 35 61 38
rect 49 34 61 35
rect 49 30 53 34
rect 57 30 61 34
rect 49 29 61 30
rect 49 26 51 29
rect 59 26 61 29
rect 69 35 71 38
rect 79 35 81 38
rect 89 35 91 38
rect 69 34 91 35
rect 69 30 82 34
rect 86 30 91 34
rect 69 29 91 30
rect 69 26 71 29
rect 79 26 81 29
rect 29 2 31 6
rect 39 2 41 6
rect 49 2 51 6
rect 59 2 61 6
rect 69 5 71 10
rect 79 5 81 10
<< ndiffusion >>
rect 21 18 29 26
rect 21 14 23 18
rect 27 14 29 18
rect 21 11 29 14
rect 21 7 23 11
rect 27 7 29 11
rect 21 6 29 7
rect 31 25 39 26
rect 31 21 33 25
rect 37 21 39 25
rect 31 18 39 21
rect 31 14 33 18
rect 37 14 39 18
rect 31 6 39 14
rect 41 18 49 26
rect 41 14 43 18
rect 47 14 49 18
rect 41 11 49 14
rect 41 7 43 11
rect 47 7 49 11
rect 41 6 49 7
rect 51 25 59 26
rect 51 21 53 25
rect 57 21 59 25
rect 51 18 59 21
rect 51 14 53 18
rect 57 14 59 18
rect 51 6 59 14
rect 61 24 69 26
rect 61 20 63 24
rect 67 20 69 24
rect 61 16 69 20
rect 61 12 63 16
rect 67 12 69 16
rect 61 10 69 12
rect 71 25 79 26
rect 71 21 73 25
rect 77 21 79 25
rect 71 17 79 21
rect 71 13 73 17
rect 77 13 79 17
rect 71 10 79 13
rect 81 23 88 26
rect 81 19 83 23
rect 87 19 88 23
rect 81 15 88 19
rect 81 11 83 15
rect 87 11 88 15
rect 81 10 88 11
rect 61 6 67 10
<< pdiffusion >>
rect 2 65 9 66
rect 2 61 3 65
rect 7 61 9 65
rect 2 58 9 61
rect 2 54 3 58
rect 7 54 9 58
rect 2 51 9 54
rect 2 47 3 51
rect 7 47 9 51
rect 2 38 9 47
rect 11 50 19 66
rect 11 46 13 50
rect 17 46 19 50
rect 11 43 19 46
rect 11 39 13 43
rect 17 39 19 43
rect 11 38 19 39
rect 21 65 29 66
rect 21 61 23 65
rect 27 61 29 65
rect 21 57 29 61
rect 21 53 23 57
rect 27 53 29 57
rect 21 38 29 53
rect 31 50 39 66
rect 31 46 33 50
rect 37 46 39 50
rect 31 43 39 46
rect 31 39 33 43
rect 37 39 39 43
rect 31 38 39 39
rect 41 65 49 66
rect 41 61 43 65
rect 47 61 49 65
rect 41 57 49 61
rect 41 53 43 57
rect 47 53 49 57
rect 41 38 49 53
rect 51 61 56 66
rect 51 50 59 61
rect 51 46 53 50
rect 57 46 59 50
rect 51 43 59 46
rect 51 39 53 43
rect 57 39 59 43
rect 51 38 59 39
rect 61 57 67 61
rect 61 56 69 57
rect 61 52 63 56
rect 67 52 69 56
rect 61 49 69 52
rect 61 45 63 49
rect 67 45 69 49
rect 61 38 69 45
rect 71 50 79 57
rect 71 46 73 50
rect 77 46 79 50
rect 71 43 79 46
rect 71 39 73 43
rect 77 39 79 43
rect 71 38 79 39
rect 81 56 89 57
rect 81 52 83 56
rect 87 52 89 56
rect 81 49 89 52
rect 81 45 83 49
rect 87 45 89 49
rect 81 38 89 45
rect 91 51 96 57
rect 91 50 98 51
rect 91 46 93 50
rect 97 46 98 50
rect 91 43 98 46
rect 91 39 93 43
rect 97 39 98 43
rect 91 38 98 39
<< metal1 >>
rect -2 68 106 72
rect -2 65 73 68
rect -2 64 3 65
rect 7 64 23 65
rect 3 58 7 61
rect 3 51 7 54
rect 27 64 43 65
rect 23 57 27 61
rect 23 52 27 53
rect 47 64 73 65
rect 77 64 92 68
rect 96 64 106 68
rect 43 57 47 61
rect 43 52 47 53
rect 62 56 68 64
rect 62 52 63 56
rect 67 52 68 56
rect 3 46 7 47
rect 13 50 17 51
rect 13 43 17 46
rect 9 39 13 42
rect 33 50 38 51
rect 37 46 38 50
rect 33 43 38 46
rect 17 39 33 42
rect 37 42 38 43
rect 53 50 57 51
rect 53 43 57 46
rect 62 49 68 52
rect 82 56 88 64
rect 82 52 83 56
rect 87 52 88 56
rect 62 45 63 49
rect 67 45 68 49
rect 73 50 77 51
rect 37 39 53 42
rect 9 38 57 39
rect 73 43 77 46
rect 82 49 88 52
rect 82 45 83 49
rect 87 45 88 49
rect 93 50 97 51
rect 93 43 97 46
rect 77 39 93 42
rect 73 38 97 39
rect 26 26 30 38
rect 73 34 77 38
rect 35 30 36 34
rect 40 30 53 34
rect 57 30 77 34
rect 81 30 82 34
rect 86 30 95 34
rect 26 25 57 26
rect 73 25 77 30
rect 26 22 33 25
rect 37 22 53 25
rect 37 21 38 22
rect 33 18 38 21
rect 53 18 57 21
rect 22 14 23 18
rect 27 14 28 18
rect 22 11 28 14
rect 37 14 38 18
rect 33 13 38 14
rect 42 14 43 18
rect 47 14 48 18
rect 22 8 23 11
rect -2 4 4 8
rect 8 4 12 8
rect 16 7 23 8
rect 27 8 28 11
rect 42 11 48 14
rect 53 13 57 14
rect 63 24 67 25
rect 63 16 67 20
rect 42 8 43 11
rect 27 7 43 8
rect 47 8 48 11
rect 73 17 77 21
rect 73 12 77 13
rect 83 23 87 24
rect 90 21 95 30
rect 83 15 87 19
rect 63 8 67 12
rect 83 8 87 11
rect 47 7 93 8
rect 16 4 93 7
rect 97 4 106 8
rect -2 0 106 4
<< ntransistor >>
rect 29 6 31 26
rect 39 6 41 26
rect 49 6 51 26
rect 59 6 61 26
rect 69 10 71 26
rect 79 10 81 26
<< ptransistor >>
rect 9 38 11 66
rect 19 38 21 66
rect 29 38 31 66
rect 39 38 41 66
rect 49 38 51 66
rect 59 38 61 61
rect 69 38 71 57
rect 79 38 81 57
rect 89 38 91 57
<< polycontact >>
rect 36 30 40 34
rect 53 30 57 34
rect 82 30 86 34
<< ndcontact >>
rect 23 14 27 18
rect 23 7 27 11
rect 33 21 37 25
rect 33 14 37 18
rect 43 14 47 18
rect 43 7 47 11
rect 53 21 57 25
rect 53 14 57 18
rect 63 20 67 24
rect 63 12 67 16
rect 73 21 77 25
rect 73 13 77 17
rect 83 19 87 23
rect 83 11 87 15
<< pdcontact >>
rect 3 61 7 65
rect 3 54 7 58
rect 3 47 7 51
rect 13 46 17 50
rect 13 39 17 43
rect 23 61 27 65
rect 23 53 27 57
rect 33 46 37 50
rect 33 39 37 43
rect 43 61 47 65
rect 43 53 47 57
rect 53 46 57 50
rect 53 39 57 43
rect 63 52 67 56
rect 63 45 67 49
rect 73 46 77 50
rect 73 39 77 43
rect 83 52 87 56
rect 83 45 87 49
rect 93 46 97 50
rect 93 39 97 43
<< psubstratepcontact >>
rect 4 4 8 8
rect 12 4 16 8
rect 93 4 97 8
<< nsubstratencontact >>
rect 73 64 77 68
rect 92 64 96 68
<< psubstratepdiff >>
rect 3 8 17 24
rect 3 4 4 8
rect 8 4 12 8
rect 16 4 17 8
rect 3 3 17 4
rect 92 8 98 24
rect 92 4 93 8
rect 97 4 98 8
rect 92 3 98 4
<< nsubstratendiff >>
rect 72 68 97 69
rect 72 64 73 68
rect 77 64 92 68
rect 96 64 97 68
rect 72 63 97 64
<< labels >>
rlabel polysilicon 35 32 35 32 6 an
rlabel polycontact 55 32 55 32 6 an
rlabel metal1 12 40 12 40 6 z
rlabel metal1 36 20 36 20 6 z
rlabel metal1 20 40 20 40 6 z
rlabel metal1 28 36 28 36 6 z
rlabel metal1 36 44 36 44 6 z
rlabel metal1 52 4 52 4 6 vss
rlabel metal1 44 24 44 24 6 z
rlabel metal1 52 24 52 24 6 z
rlabel metal1 44 40 44 40 6 z
rlabel metal1 52 40 52 40 6 z
rlabel metal1 52 68 52 68 6 vdd
rlabel polycontact 56 32 56 32 6 an
rlabel metal1 75 31 75 31 6 an
rlabel metal1 92 28 92 28 6 a
rlabel polycontact 84 32 84 32 6 a
rlabel metal1 95 44 95 44 6 an
<< end >>
