.subckt nd2v5x6 a b vdd vss z
*   SPICE3 file   created from nd2v5x6.ext -      technology: scmos
m00 z      b      vdd    vdd p w=27u  l=2.3636u ad=108p     pd=35u      as=135p     ps=46u
m01 vdd    a      z      vdd p w=27u  l=2.3636u ad=135p     pd=46u      as=108p     ps=35u
m02 z      a      vdd    vdd p w=27u  l=2.3636u ad=108p     pd=35u      as=135p     ps=46u
m03 vdd    b      z      vdd p w=27u  l=2.3636u ad=135p     pd=46u      as=108p     ps=35u
m04 z      b      vdd    vdd p w=27u  l=2.3636u ad=108p     pd=35u      as=135p     ps=46u
m05 vdd    a      z      vdd p w=27u  l=2.3636u ad=135p     pd=46u      as=108p     ps=35u
m06 w1     b      z      vss n w=11u  l=2.3636u ad=27.5p    pd=16u      as=48.9608p ps=19.8431u
m07 vss    a      w1     vss n w=11u  l=2.3636u ad=82.6078p pd=26.7451u as=27.5p    ps=16u
m08 w2     a      vss    vss n w=20u  l=2.3636u ad=50p      pd=25u      as=150.196p ps=48.6275u
m09 z      b      w2     vss n w=20u  l=2.3636u ad=89.0196p pd=36.0784u as=50p      ps=25u
m10 w3     b      z      vss n w=20u  l=2.3636u ad=50p      pd=25u      as=89.0196p ps=36.0784u
m11 vss    a      w3     vss n w=20u  l=2.3636u ad=150.196p pd=48.6275u as=50p      ps=25u
C0  w2     b      0.007f
C1  vss    a      0.051f
C2  w1     b      0.005f
C3  z      a      0.396f
C4  vdd    b      0.056f
C5  w2     vss    0.005f
C6  w2     z      0.010f
C7  w1     z      0.006f
C8  w3     b      0.007f
C9  vss    vdd    0.004f
C10 vss    b      0.117f
C11 z      vdd    0.683f
C12 z      b      0.456f
C13 vdd    a      0.102f
C14 w3     vss    0.005f
C15 a      b      0.491f
C16 vss    z      0.310f
C18 z      vss    0.009f
C20 a      vss    0.048f
C21 b      vss    0.049f
.ends
