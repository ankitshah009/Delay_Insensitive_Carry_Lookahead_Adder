magic
tech scmos
timestamp 1185039033
<< checkpaint >>
rect -22 -24 72 124
<< ab >>
rect 0 0 50 100
<< pwell >>
rect -2 -4 52 49
<< nwell >>
rect -2 49 52 104
<< polysilicon >>
rect 19 95 21 98
rect 27 95 29 98
rect 35 95 37 98
rect 19 53 21 55
rect 17 52 23 53
rect 17 49 18 52
rect 11 48 18 49
rect 22 48 23 52
rect 11 47 23 48
rect 11 25 13 47
rect 27 43 29 55
rect 35 53 37 55
rect 35 51 39 53
rect 27 42 33 43
rect 27 39 28 42
rect 23 38 28 39
rect 32 38 33 42
rect 23 37 33 38
rect 23 25 25 37
rect 37 33 39 51
rect 37 32 43 33
rect 37 29 38 32
rect 35 28 38 29
rect 42 28 43 32
rect 35 27 43 28
rect 35 25 37 27
rect 11 12 13 15
rect 23 12 25 15
rect 35 12 37 15
<< ndiffusion >>
rect 3 22 11 25
rect 3 18 4 22
rect 8 18 11 22
rect 3 15 11 18
rect 13 15 23 25
rect 25 22 35 25
rect 25 18 28 22
rect 32 18 35 22
rect 25 15 35 18
rect 37 15 45 25
rect 15 12 21 15
rect 39 12 45 15
rect 15 8 16 12
rect 20 8 21 12
rect 15 7 21 8
rect 39 8 40 12
rect 44 8 45 12
rect 39 7 45 8
<< pdiffusion >>
rect 15 85 19 95
rect 7 82 19 85
rect 7 78 8 82
rect 12 78 19 82
rect 7 72 19 78
rect 7 68 8 72
rect 12 68 19 72
rect 7 62 19 68
rect 7 58 8 62
rect 12 58 19 62
rect 7 55 19 58
rect 21 55 27 95
rect 29 55 35 95
rect 37 92 45 95
rect 37 88 40 92
rect 44 88 45 92
rect 37 55 45 88
<< metal1 >>
rect -2 92 52 101
rect -2 88 40 92
rect 44 88 52 92
rect -2 87 52 88
rect 7 82 13 83
rect 7 78 8 82
rect 12 78 13 82
rect 7 72 13 78
rect 7 68 8 72
rect 12 68 13 72
rect 7 62 13 68
rect 7 58 8 62
rect 12 58 13 62
rect 7 23 13 58
rect 17 52 23 82
rect 17 48 18 52
rect 22 48 23 52
rect 17 28 23 48
rect 27 42 33 82
rect 27 38 28 42
rect 32 38 33 42
rect 27 28 33 38
rect 37 32 43 82
rect 37 28 38 32
rect 42 28 43 32
rect 3 22 33 23
rect 3 18 4 22
rect 8 18 28 22
rect 32 18 33 22
rect 37 18 43 28
rect 3 17 33 18
rect -2 12 52 13
rect -2 8 16 12
rect 20 8 40 12
rect 44 8 52 12
rect -2 -1 52 8
<< ntransistor >>
rect 11 15 13 25
rect 23 15 25 25
rect 35 15 37 25
<< ptransistor >>
rect 19 55 21 95
rect 27 55 29 95
rect 35 55 37 95
<< polycontact >>
rect 18 48 22 52
rect 28 38 32 42
rect 38 28 42 32
<< ndcontact >>
rect 4 18 8 22
rect 28 18 32 22
rect 16 8 20 12
rect 40 8 44 12
<< pdcontact >>
rect 8 78 12 82
rect 8 68 12 72
rect 8 58 12 62
rect 40 88 44 92
<< labels >>
rlabel metal1 10 50 10 50 6 nq
rlabel metal1 10 50 10 50 6 nq
rlabel metal1 20 55 20 55 6 i1
rlabel metal1 20 55 20 55 6 i1
rlabel metal1 25 6 25 6 6 vss
rlabel metal1 25 6 25 6 6 vss
rlabel metal1 30 55 30 55 6 i0
rlabel metal1 30 55 30 55 6 i0
rlabel metal1 25 94 25 94 6 vdd
rlabel metal1 25 94 25 94 6 vdd
rlabel metal1 40 50 40 50 6 i2
rlabel metal1 40 50 40 50 6 i2
<< end >>
