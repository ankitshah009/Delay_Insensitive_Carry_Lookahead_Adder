.subckt xnr2v0x3 a b vdd vss z
*   SPICE3 file   created from xnr2v0x3.ext -      technology: scmos
m00 w1     an     z      vdd p w=28u  l=2.3636u ad=70p      pd=33u      as=122.8p   ps=42.8u
m01 vdd    bn     w1     vdd p w=28u  l=2.3636u ad=148p     pd=42.5714u as=70p      ps=33u
m02 w2     bn     vdd    vdd p w=28u  l=2.3636u ad=70p      pd=33u      as=148p     ps=42.5714u
m03 z      an     w2     vdd p w=28u  l=2.3636u ad=122.8p   pd=42.8u    as=70p      ps=33u
m04 w3     an     z      vdd p w=28u  l=2.3636u ad=70p      pd=33u      as=122.8p   ps=42.8u
m05 vdd    bn     w3     vdd p w=28u  l=2.3636u ad=148p     pd=42.5714u as=70p      ps=33u
m06 an     a      vdd    vdd p w=28u  l=2.3636u ad=112p     pd=36u      as=148p     ps=42.5714u
m07 z      b      an     vdd p w=28u  l=2.3636u ad=122.8p   pd=42.8u    as=112p     ps=36u
m08 an     b      z      vdd p w=28u  l=2.3636u ad=112p     pd=36u      as=122.8p   ps=42.8u
m09 vdd    a      an     vdd p w=28u  l=2.3636u ad=148p     pd=42.5714u as=112p     ps=36u
m10 bn     b      vdd    vdd p w=28u  l=2.3636u ad=112p     pd=36u      as=148p     ps=42.5714u
m11 vdd    b      bn     vdd p w=28u  l=2.3636u ad=148p     pd=42.5714u as=112p     ps=36u
m12 z      bn     an     vss n w=14u  l=2.3636u ad=56p      pd=22u      as=73p      ps=32u
m13 bn     an     z      vss n w=14u  l=2.3636u ad=56p      pd=22u      as=56p      ps=22u
m14 z      an     bn     vss n w=14u  l=2.3636u ad=56p      pd=22u      as=56p      ps=22u
m15 an     bn     z      vss n w=14u  l=2.3636u ad=73p      pd=32u      as=56p      ps=22u
m16 vss    a      an     vss n w=14u  l=2.3636u ad=96.5p    pd=36.5u    as=73p      ps=32u
m17 vss    a      an     vss n w=14u  l=2.3636u ad=96.5p    pd=36.5u    as=73p      ps=32u
m18 bn     b      vss    vss n w=14u  l=2.3636u ad=56p      pd=22u      as=96.5p    ps=36.5u
m19 vss    b      bn     vss n w=14u  l=2.3636u ad=96.5p    pd=36.5u    as=56p      ps=22u
C0  w2     bn     0.019f
C1  vss    vdd    0.008f
C2  z      b      0.009f
C3  w2     vdd    0.005f
C4  b      a      0.175f
C5  z      bn     1.132f
C6  b      an     0.205f
C7  a      bn     0.177f
C8  z      vdd    0.540f
C9  vss    z      0.085f
C10 bn     an     0.803f
C11 a      vdd    0.020f
C12 vss    a      0.060f
C13 w2     z      0.010f
C14 an     vdd    0.077f
C15 w3     bn     0.010f
C16 vss    an     0.640f
C17 z      a      0.077f
C18 w3     vdd    0.005f
C19 w1     vdd    0.005f
C20 b      bn     0.209f
C21 z      an     0.426f
C22 a      an     0.277f
C23 b      vdd    0.056f
C24 w3     z      0.018f
C25 vss    b      0.054f
C26 bn     vdd    0.312f
C27 w1     z      0.007f
C28 vss    bn     0.239f
C30 z      vss    0.013f
C31 b      vss    0.059f
C32 a      vss    0.042f
C33 bn     vss    0.047f
C34 an     vss    0.069f
.ends
