magic
tech scmos
timestamp 1185039168
<< checkpaint >>
rect -22 -24 142 124
<< ab >>
rect 0 0 120 100
<< pwell >>
rect -2 -4 122 49
<< nwell >>
rect -2 49 122 104
<< polysilicon >>
rect 23 95 25 98
rect 35 95 37 98
rect 47 95 49 98
rect 59 95 61 98
rect 11 75 13 78
rect 95 95 97 98
rect 107 95 109 98
rect 71 75 73 78
rect 11 53 13 55
rect 23 53 25 55
rect 11 52 25 53
rect 11 51 18 52
rect 17 48 18 51
rect 22 51 25 52
rect 35 53 37 55
rect 35 52 43 53
rect 35 51 38 52
rect 22 48 23 51
rect 17 47 23 48
rect 37 48 38 51
rect 42 48 43 52
rect 37 47 43 48
rect 3 42 9 43
rect 3 38 4 42
rect 8 41 9 42
rect 47 41 49 55
rect 59 43 61 55
rect 71 53 73 55
rect 67 52 73 53
rect 67 48 68 52
rect 72 48 73 52
rect 67 47 73 48
rect 95 43 97 55
rect 107 43 109 55
rect 8 39 49 41
rect 8 38 9 39
rect 3 37 9 38
rect 17 32 23 33
rect 17 29 18 32
rect 11 28 18 29
rect 22 29 23 32
rect 37 32 43 33
rect 37 29 38 32
rect 22 28 25 29
rect 11 27 25 28
rect 11 25 13 27
rect 23 25 25 27
rect 35 28 38 29
rect 42 28 43 32
rect 35 27 43 28
rect 35 25 37 27
rect 47 25 49 39
rect 57 42 63 43
rect 57 38 58 42
rect 62 41 63 42
rect 77 42 83 43
rect 77 41 78 42
rect 62 39 78 41
rect 62 38 63 39
rect 57 37 63 38
rect 77 38 78 39
rect 82 38 83 42
rect 77 37 83 38
rect 87 42 109 43
rect 87 38 88 42
rect 92 38 109 42
rect 87 37 109 38
rect 67 32 73 33
rect 67 29 68 32
rect 59 28 68 29
rect 72 28 73 32
rect 59 27 73 28
rect 59 25 61 27
rect 71 25 73 27
rect 95 25 97 37
rect 107 25 109 37
rect 11 12 13 15
rect 71 12 73 15
rect 23 2 25 5
rect 35 2 37 5
rect 47 2 49 5
rect 59 2 61 5
rect 95 2 97 5
rect 107 2 109 5
<< ndiffusion >>
rect 75 32 83 33
rect 75 28 78 32
rect 82 28 83 32
rect 75 27 83 28
rect 75 25 81 27
rect 3 22 11 25
rect 3 18 4 22
rect 8 18 11 22
rect 3 15 11 18
rect 13 15 23 25
rect 15 12 23 15
rect 15 8 16 12
rect 20 8 23 12
rect 15 5 23 8
rect 25 5 35 25
rect 37 22 47 25
rect 37 18 40 22
rect 44 18 47 22
rect 37 5 47 18
rect 49 5 59 25
rect 61 15 71 25
rect 73 15 81 25
rect 91 21 95 25
rect 61 12 69 15
rect 87 12 95 21
rect 61 8 64 12
rect 68 8 69 12
rect 61 5 69 8
rect 87 8 88 12
rect 92 8 95 12
rect 87 5 95 8
rect 97 22 107 25
rect 97 18 100 22
rect 104 18 107 22
rect 97 5 107 18
rect 109 22 117 25
rect 109 18 112 22
rect 116 18 117 22
rect 109 12 117 18
rect 109 8 112 12
rect 116 8 117 12
rect 109 5 117 8
<< pdiffusion >>
rect 15 92 23 95
rect 15 88 16 92
rect 20 88 23 92
rect 15 75 23 88
rect 3 72 11 75
rect 3 68 4 72
rect 8 68 11 72
rect 3 62 11 68
rect 3 58 4 62
rect 8 58 11 62
rect 3 55 11 58
rect 13 55 23 75
rect 25 82 35 95
rect 25 78 28 82
rect 32 78 35 82
rect 25 72 35 78
rect 25 68 28 72
rect 32 68 35 72
rect 25 55 35 68
rect 37 72 47 95
rect 37 68 40 72
rect 44 68 47 72
rect 37 55 47 68
rect 49 82 59 95
rect 49 78 52 82
rect 56 78 59 82
rect 49 72 59 78
rect 49 68 52 72
rect 56 68 59 72
rect 49 62 59 68
rect 49 58 52 62
rect 56 58 59 62
rect 49 55 59 58
rect 61 92 69 95
rect 61 88 64 92
rect 68 88 69 92
rect 61 75 69 88
rect 87 92 95 95
rect 87 88 88 92
rect 92 88 95 92
rect 87 82 95 88
rect 87 78 88 82
rect 92 78 95 82
rect 61 55 71 75
rect 73 61 81 75
rect 87 72 95 78
rect 87 68 88 72
rect 92 68 95 72
rect 87 67 95 68
rect 73 60 83 61
rect 73 56 78 60
rect 82 56 83 60
rect 73 55 83 56
rect 91 55 95 67
rect 97 82 107 95
rect 97 78 100 82
rect 104 78 107 82
rect 97 72 107 78
rect 97 68 100 72
rect 104 68 107 72
rect 97 62 107 68
rect 97 58 100 62
rect 104 58 107 62
rect 97 55 107 58
rect 109 92 117 95
rect 109 88 112 92
rect 116 88 117 92
rect 109 82 117 88
rect 109 78 112 82
rect 116 78 117 82
rect 109 72 117 78
rect 109 68 112 72
rect 116 68 117 72
rect 109 62 117 68
rect 109 58 112 62
rect 116 58 117 62
rect 109 55 117 58
<< metal1 >>
rect -2 96 122 101
rect -2 92 4 96
rect 8 92 76 96
rect 80 92 122 96
rect -2 88 16 92
rect 20 88 64 92
rect 68 88 88 92
rect 92 88 112 92
rect 116 88 122 92
rect -2 87 122 88
rect 27 82 33 83
rect 51 82 57 83
rect 87 82 93 87
rect 99 82 105 83
rect 3 72 9 73
rect 3 68 4 72
rect 8 68 9 72
rect 3 67 9 68
rect 4 63 8 67
rect 3 62 9 63
rect 3 58 4 62
rect 8 58 9 62
rect 3 57 9 58
rect 4 43 8 57
rect 17 52 23 82
rect 27 78 28 82
rect 32 78 52 82
rect 56 78 57 82
rect 27 77 33 78
rect 51 77 57 78
rect 28 73 32 77
rect 52 73 56 77
rect 27 72 33 73
rect 27 68 28 72
rect 32 68 33 72
rect 27 67 33 68
rect 39 72 45 73
rect 39 68 40 72
rect 44 68 45 72
rect 39 67 45 68
rect 51 72 57 73
rect 51 68 52 72
rect 56 68 57 72
rect 51 67 57 68
rect 40 62 44 67
rect 52 63 56 67
rect 17 48 18 52
rect 22 48 23 52
rect 3 42 9 43
rect 3 38 4 42
rect 8 38 9 42
rect 3 37 9 38
rect 4 23 8 37
rect 17 32 23 48
rect 17 28 18 32
rect 22 28 23 32
rect 3 22 9 23
rect 3 18 4 22
rect 8 18 9 22
rect 17 18 23 28
rect 28 58 44 62
rect 51 62 57 63
rect 51 58 52 62
rect 56 58 57 62
rect 28 22 32 58
rect 51 57 57 58
rect 37 52 43 53
rect 67 52 73 82
rect 87 78 88 82
rect 92 78 93 82
rect 87 72 93 78
rect 87 68 88 72
rect 92 68 93 72
rect 87 67 93 68
rect 97 78 100 82
rect 104 78 105 82
rect 97 77 105 78
rect 111 82 117 87
rect 111 78 112 82
rect 116 78 117 82
rect 97 73 103 77
rect 97 72 105 73
rect 97 68 100 72
rect 104 68 105 72
rect 97 67 105 68
rect 111 72 117 78
rect 111 68 112 72
rect 116 68 117 72
rect 97 63 103 67
rect 97 62 105 63
rect 77 60 83 61
rect 77 56 78 60
rect 82 56 83 60
rect 77 55 83 56
rect 97 58 100 62
rect 104 58 105 62
rect 97 57 105 58
rect 111 62 117 68
rect 111 58 112 62
rect 116 58 117 62
rect 111 57 117 58
rect 37 48 38 52
rect 42 48 68 52
rect 72 48 73 52
rect 37 47 43 48
rect 57 42 63 43
rect 48 38 58 42
rect 62 38 63 42
rect 37 32 43 33
rect 48 32 52 38
rect 57 37 63 38
rect 37 28 38 32
rect 42 28 52 32
rect 67 32 73 48
rect 78 43 82 55
rect 77 42 83 43
rect 77 38 78 42
rect 82 38 83 42
rect 77 37 83 38
rect 87 42 93 43
rect 87 38 88 42
rect 92 38 93 42
rect 87 37 93 38
rect 78 33 82 37
rect 67 28 68 32
rect 72 28 73 32
rect 37 27 43 28
rect 67 27 73 28
rect 77 32 83 33
rect 77 28 78 32
rect 82 28 83 32
rect 77 27 83 28
rect 39 22 45 23
rect 88 22 92 37
rect 28 18 40 22
rect 44 18 92 22
rect 97 23 103 57
rect 97 22 105 23
rect 97 18 100 22
rect 104 18 105 22
rect 3 17 9 18
rect 39 17 45 18
rect 99 17 105 18
rect 111 22 117 23
rect 111 18 112 22
rect 116 18 117 22
rect 111 13 117 18
rect -2 12 122 13
rect -2 8 16 12
rect 20 8 64 12
rect 68 8 88 12
rect 92 8 112 12
rect 116 8 122 12
rect -2 -1 122 8
<< ntransistor >>
rect 11 15 13 25
rect 23 5 25 25
rect 35 5 37 25
rect 47 5 49 25
rect 59 5 61 25
rect 71 15 73 25
rect 95 5 97 25
rect 107 5 109 25
<< ptransistor >>
rect 11 55 13 75
rect 23 55 25 95
rect 35 55 37 95
rect 47 55 49 95
rect 59 55 61 95
rect 71 55 73 75
rect 95 55 97 95
rect 107 55 109 95
<< polycontact >>
rect 18 48 22 52
rect 38 48 42 52
rect 4 38 8 42
rect 68 48 72 52
rect 18 28 22 32
rect 38 28 42 32
rect 58 38 62 42
rect 78 38 82 42
rect 88 38 92 42
rect 68 28 72 32
<< ndcontact >>
rect 78 28 82 32
rect 4 18 8 22
rect 16 8 20 12
rect 40 18 44 22
rect 64 8 68 12
rect 88 8 92 12
rect 100 18 104 22
rect 112 18 116 22
rect 112 8 116 12
<< pdcontact >>
rect 16 88 20 92
rect 4 68 8 72
rect 4 58 8 62
rect 28 78 32 82
rect 28 68 32 72
rect 40 68 44 72
rect 52 78 56 82
rect 52 68 56 72
rect 52 58 56 62
rect 64 88 68 92
rect 88 88 92 92
rect 88 78 92 82
rect 88 68 92 72
rect 78 56 82 60
rect 100 78 104 82
rect 100 68 104 72
rect 100 58 104 62
rect 112 88 116 92
rect 112 78 116 82
rect 112 68 116 72
rect 112 58 116 62
<< nsubstratencontact >>
rect 4 92 8 96
rect 76 92 80 96
<< nsubstratendiff >>
rect 3 96 9 97
rect 3 92 4 96
rect 8 92 9 96
rect 75 96 81 97
rect 3 85 9 92
rect 75 92 76 96
rect 80 92 81 96
rect 75 85 81 92
<< labels >>
rlabel polycontact 20 50 20 50 6 i0
rlabel polycontact 20 50 20 50 6 i0
rlabel metal1 60 6 60 6 6 vss
rlabel metal1 60 6 60 6 6 vss
rlabel metal1 70 55 70 55 6 i1
rlabel metal1 70 55 70 55 6 i1
rlabel metal1 60 94 60 94 6 vdd
rlabel metal1 60 94 60 94 6 vdd
rlabel metal1 100 50 100 50 6 q
rlabel metal1 100 50 100 50 6 q
<< end >>
