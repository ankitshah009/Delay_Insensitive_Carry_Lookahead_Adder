.subckt tie_x0 vdd vss
*   SPICE3 file   created from tie_x0.ext -      technology: scmos
.ends
