magic
tech scmos
timestamp 1179386545
<< checkpaint >>
rect -22 -22 86 94
<< ab >>
rect 0 0 64 72
<< pwell >>
rect -4 -4 68 32
<< nwell >>
rect -4 32 68 76
<< polysilicon >>
rect 11 66 13 70
rect 21 66 23 70
rect 37 66 39 70
rect 49 66 51 70
rect 11 49 13 52
rect 21 49 23 52
rect 11 48 23 49
rect 11 47 18 48
rect 17 44 18 47
rect 22 44 23 48
rect 17 43 23 44
rect 9 34 15 35
rect 9 30 10 34
rect 14 30 15 34
rect 9 29 15 30
rect 12 26 14 29
rect 19 26 21 43
rect 37 35 39 38
rect 33 34 39 35
rect 33 31 34 34
rect 26 30 34 31
rect 38 30 39 34
rect 49 35 51 38
rect 49 34 55 35
rect 26 29 39 30
rect 26 26 28 29
rect 36 26 38 29
rect 43 26 45 31
rect 49 30 50 34
rect 54 30 55 34
rect 49 29 55 30
rect 50 26 52 29
rect 12 7 14 12
rect 19 4 21 12
rect 26 8 28 12
rect 36 8 38 12
rect 43 4 45 12
rect 50 7 52 12
rect 19 2 45 4
<< ndiffusion >>
rect 2 17 12 26
rect 2 13 3 17
rect 7 13 12 17
rect 2 12 12 13
rect 14 12 19 26
rect 21 12 26 26
rect 28 18 36 26
rect 28 14 30 18
rect 34 14 36 18
rect 28 12 36 14
rect 38 12 43 26
rect 45 12 50 26
rect 52 17 60 26
rect 52 13 54 17
rect 58 13 60 17
rect 52 12 60 13
<< pdiffusion >>
rect 3 65 11 66
rect 3 61 5 65
rect 9 61 11 65
rect 3 52 11 61
rect 13 58 21 66
rect 13 54 15 58
rect 19 54 21 58
rect 13 52 21 54
rect 23 65 37 66
rect 23 61 28 65
rect 32 61 37 65
rect 23 52 37 61
rect 25 38 37 52
rect 39 58 49 66
rect 39 54 42 58
rect 46 54 49 58
rect 39 50 49 54
rect 39 46 42 50
rect 46 46 49 50
rect 39 38 49 46
rect 51 65 59 66
rect 51 61 53 65
rect 57 61 59 65
rect 51 58 59 61
rect 51 54 53 58
rect 57 54 59 58
rect 51 38 59 54
<< metal1 >>
rect -2 65 66 72
rect -2 64 5 65
rect 4 61 5 64
rect 9 64 28 65
rect 9 61 10 64
rect 27 61 28 64
rect 32 64 53 65
rect 32 61 33 64
rect 52 61 53 64
rect 57 64 66 65
rect 57 61 58 64
rect 52 58 58 61
rect 2 54 15 58
rect 19 54 42 58
rect 46 54 47 58
rect 52 54 53 58
rect 57 54 58 58
rect 2 25 6 54
rect 41 50 47 54
rect 17 48 23 50
rect 17 44 18 48
rect 22 44 23 48
rect 41 46 42 50
rect 46 46 47 50
rect 17 42 23 44
rect 17 38 31 42
rect 38 38 47 42
rect 10 34 16 35
rect 14 30 26 34
rect 33 30 34 34
rect 38 30 42 38
rect 49 30 50 34
rect 54 30 55 34
rect 10 29 26 30
rect 22 26 26 29
rect 49 26 55 30
rect 2 21 15 25
rect 22 22 55 26
rect 11 18 15 21
rect 3 17 7 18
rect 11 14 30 18
rect 34 14 35 18
rect 54 17 58 18
rect 3 8 7 13
rect 54 8 58 13
rect -2 0 66 8
<< ntransistor >>
rect 12 12 14 26
rect 19 12 21 26
rect 26 12 28 26
rect 36 12 38 26
rect 43 12 45 26
rect 50 12 52 26
<< ptransistor >>
rect 11 52 13 66
rect 21 52 23 66
rect 37 38 39 66
rect 49 38 51 66
<< polycontact >>
rect 18 44 22 48
rect 10 30 14 34
rect 34 30 38 34
rect 50 30 54 34
<< ndcontact >>
rect 3 13 7 17
rect 30 14 34 18
rect 54 13 58 17
<< pdcontact >>
rect 5 61 9 65
rect 15 54 19 58
rect 28 61 32 65
rect 42 54 46 58
rect 42 46 46 50
rect 53 61 57 65
rect 53 54 57 58
<< labels >>
rlabel metal1 4 36 4 36 6 z
rlabel metal1 20 16 20 16 6 z
rlabel metal1 20 32 20 32 6 a
rlabel metal1 20 44 20 44 6 b
rlabel metal1 20 56 20 56 6 z
rlabel metal1 12 56 12 56 6 z
rlabel metal1 32 4 32 4 6 vss
rlabel metal1 28 16 28 16 6 z
rlabel metal1 28 24 28 24 6 a
rlabel metal1 36 24 36 24 6 a
rlabel metal1 28 40 28 40 6 b
rlabel metal1 36 56 36 56 6 z
rlabel metal1 28 56 28 56 6 z
rlabel metal1 32 68 32 68 6 vdd
rlabel metal1 44 24 44 24 6 a
rlabel metal1 44 40 44 40 6 c
rlabel metal1 44 52 44 52 6 z
rlabel metal1 52 28 52 28 6 a
<< end >>
