.subckt tie_x0 vdd vss
*   SPICE3 file   created from tie_x0.ext -      technology: scmos
m00 w1     vdd    w2     vdd p w=26u  l=2.3636u ad=130p     pd=36u      as=182p     ps=66u
m01 w3     vdd    w1     vdd p w=26u  l=2.3636u ad=182p     pd=66u      as=130p     ps=36u
m02 w4     vdd    w5     vdd p w=26u  l=2.3636u ad=130p     pd=36u      as=182p     ps=66u
m03 w6     vdd    w4     vdd p w=26u  l=2.3636u ad=182p     pd=66u      as=130p     ps=36u
m04 w7     vss    w8     vss n w=18u  l=2.3636u ad=90p      pd=28u      as=126p     ps=50u
m05 w9     vss    w7     vss n w=18u  l=2.3636u ad=126p     pd=50u      as=90p      ps=28u
m06 w10    vss    w11    vss n w=18u  l=2.3636u ad=90p      pd=28u      as=126p     ps=50u
m07 w12    vss    w10    vss n w=18u  l=2.3636u ad=126p     pd=50u      as=90p      ps=28u
C0  vss    vdd    0.193f
.ends
