.subckt vfeed7 vdd vss
*   SPICE3 file   created from vfeed7.ext -      technology: scmos
.ends
