magic
tech scmos
timestamp 1179386717
<< checkpaint >>
rect -22 -22 70 94
<< ab >>
rect 0 0 48 72
<< pwell >>
rect -4 -4 52 32
<< nwell >>
rect -4 32 52 76
<< polysilicon >>
rect 12 59 14 64
rect 19 59 21 64
rect 33 56 35 61
rect 12 38 14 44
rect 9 37 15 38
rect 9 33 10 37
rect 14 33 15 37
rect 9 32 15 33
rect 11 18 13 32
rect 19 27 21 44
rect 33 38 35 44
rect 25 37 35 38
rect 25 33 26 37
rect 30 33 35 37
rect 25 32 35 33
rect 17 26 23 27
rect 33 26 35 32
rect 17 22 18 26
rect 22 22 23 26
rect 17 21 23 22
rect 21 18 23 21
rect 33 15 35 20
rect 11 5 13 10
rect 21 5 23 10
<< ndiffusion >>
rect 25 20 33 26
rect 35 25 42 26
rect 35 21 37 25
rect 41 21 42 25
rect 35 20 42 21
rect 25 18 31 20
rect 3 10 11 18
rect 13 17 21 18
rect 13 13 15 17
rect 19 13 21 17
rect 13 10 21 13
rect 23 16 31 18
rect 23 12 26 16
rect 30 12 31 16
rect 23 10 31 12
rect 3 8 9 10
rect 3 4 4 8
rect 8 4 9 8
rect 3 3 9 4
<< pdiffusion >>
rect 5 58 12 59
rect 5 54 6 58
rect 10 54 12 58
rect 5 53 12 54
rect 7 44 12 53
rect 14 44 19 59
rect 21 58 31 59
rect 21 54 26 58
rect 30 56 31 58
rect 30 54 33 56
rect 21 51 33 54
rect 21 47 27 51
rect 31 47 33 51
rect 21 44 33 47
rect 35 50 40 56
rect 35 49 42 50
rect 35 45 37 49
rect 41 45 42 49
rect 35 44 42 45
<< metal1 >>
rect -2 68 50 72
rect -2 64 28 68
rect 32 64 36 68
rect 40 64 50 68
rect 2 58 14 59
rect 2 54 6 58
rect 10 54 14 58
rect 2 53 14 54
rect 26 58 32 64
rect 30 54 32 58
rect 2 18 6 53
rect 26 51 32 54
rect 18 43 22 51
rect 26 47 27 51
rect 31 47 32 51
rect 37 49 41 50
rect 10 39 22 43
rect 10 37 14 39
rect 26 37 30 43
rect 10 29 14 33
rect 18 33 26 35
rect 18 29 30 33
rect 37 26 41 45
rect 17 22 18 26
rect 22 25 41 26
rect 22 22 37 25
rect 37 20 41 21
rect 2 17 23 18
rect 2 13 15 17
rect 19 13 23 17
rect 26 16 30 17
rect 26 8 30 12
rect -2 4 4 8
rect 8 4 36 8
rect 40 4 50 8
rect -2 0 50 4
<< ntransistor >>
rect 33 20 35 26
rect 11 10 13 18
rect 21 10 23 18
<< ptransistor >>
rect 12 44 14 59
rect 19 44 21 59
rect 33 44 35 56
<< polycontact >>
rect 10 33 14 37
rect 26 33 30 37
rect 18 22 22 26
<< ndcontact >>
rect 37 21 41 25
rect 15 13 19 17
rect 26 12 30 16
rect 4 4 8 8
<< pdcontact >>
rect 6 54 10 58
rect 26 54 30 58
rect 27 47 31 51
rect 37 45 41 49
<< psubstratepcontact >>
rect 36 4 40 8
<< nsubstratencontact >>
rect 28 64 32 68
rect 36 64 40 68
<< psubstratepdiff >>
rect 35 8 41 13
rect 35 4 36 8
rect 40 4 41 8
rect 35 3 41 4
<< nsubstratendiff >>
rect 27 68 41 69
rect 27 64 28 68
rect 32 64 36 68
rect 40 64 41 68
rect 27 63 41 64
<< labels >>
rlabel polycontact 20 24 20 24 6 an
rlabel metal1 4 36 4 36 6 z
rlabel metal1 20 16 20 16 6 z
rlabel metal1 12 16 12 16 6 z
rlabel metal1 20 32 20 32 6 a
rlabel polycontact 12 36 12 36 6 b
rlabel metal1 20 48 20 48 6 b
rlabel metal1 12 56 12 56 6 z
rlabel metal1 24 4 24 4 6 vss
rlabel polycontact 28 36 28 36 6 a
rlabel metal1 24 68 24 68 6 vdd
rlabel metal1 29 24 29 24 6 an
rlabel metal1 39 35 39 35 6 an
<< end >>
