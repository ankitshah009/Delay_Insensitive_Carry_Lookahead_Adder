magic
tech scmos
timestamp 1185094796
<< checkpaint >>
rect -22 -22 92 122
<< ab >>
rect 0 0 70 100
<< pwell >>
rect -4 -4 74 48
<< nwell >>
rect -4 48 74 104
<< polysilicon >>
rect 21 93 23 98
rect 45 93 47 98
rect 53 93 55 98
rect 33 75 35 80
rect 21 42 23 55
rect 33 52 35 55
rect 33 51 41 52
rect 33 47 36 51
rect 40 47 41 51
rect 33 46 41 47
rect 11 41 31 42
rect 11 40 26 41
rect 11 36 13 40
rect 25 37 26 40
rect 30 37 31 41
rect 25 36 31 37
rect 35 33 37 46
rect 45 43 47 55
rect 53 52 55 55
rect 53 51 63 52
rect 53 50 58 51
rect 57 47 58 50
rect 62 47 63 51
rect 57 46 63 47
rect 45 42 53 43
rect 45 38 48 42
rect 52 38 53 42
rect 45 37 53 38
rect 47 33 49 37
rect 57 33 59 46
rect 11 11 13 17
rect 35 11 37 16
rect 47 11 49 16
rect 57 11 59 16
<< ndiffusion >>
rect 3 32 11 36
rect 3 28 4 32
rect 8 28 11 32
rect 3 22 11 28
rect 3 18 4 22
rect 8 18 11 22
rect 3 17 11 18
rect 13 35 21 36
rect 13 31 16 35
rect 20 31 21 35
rect 13 27 21 31
rect 13 23 16 27
rect 20 23 21 27
rect 13 22 21 23
rect 27 32 35 33
rect 27 28 28 32
rect 32 28 35 32
rect 27 24 35 28
rect 13 17 18 22
rect 27 20 28 24
rect 32 20 35 24
rect 27 19 35 20
rect 30 16 35 19
rect 37 22 47 33
rect 37 18 40 22
rect 44 18 47 22
rect 37 16 47 18
rect 49 16 57 33
rect 59 32 67 33
rect 59 28 62 32
rect 66 28 67 32
rect 59 24 67 28
rect 59 20 62 24
rect 66 20 67 24
rect 59 19 67 20
rect 59 16 64 19
rect 51 9 55 16
rect 51 8 57 9
rect 51 4 52 8
rect 56 4 57 8
rect 51 3 57 4
<< pdiffusion >>
rect 16 71 21 93
rect 13 70 21 71
rect 13 66 14 70
rect 18 66 21 70
rect 13 62 21 66
rect 13 58 14 62
rect 18 58 21 62
rect 13 57 21 58
rect 16 55 21 57
rect 23 92 31 93
rect 23 88 26 92
rect 30 88 31 92
rect 23 82 31 88
rect 23 78 26 82
rect 30 78 31 82
rect 23 75 31 78
rect 40 75 45 93
rect 23 72 33 75
rect 23 68 26 72
rect 30 68 33 72
rect 23 55 33 68
rect 35 72 45 75
rect 35 68 38 72
rect 42 68 45 72
rect 35 64 45 68
rect 35 60 38 64
rect 42 60 45 64
rect 35 55 45 60
rect 47 55 53 93
rect 55 92 63 93
rect 55 88 58 92
rect 62 88 63 92
rect 55 82 63 88
rect 55 78 58 82
rect 62 78 63 82
rect 55 55 63 78
<< metal1 >>
rect -2 96 72 100
rect -2 92 4 96
rect 8 92 72 96
rect -2 88 26 92
rect 30 88 58 92
rect 62 88 72 92
rect 26 82 30 88
rect 26 72 30 78
rect 58 82 62 88
rect 58 77 62 78
rect 14 70 18 71
rect 26 67 30 68
rect 38 72 42 73
rect 47 68 62 73
rect 14 63 18 66
rect 38 64 42 68
rect 8 62 22 63
rect 8 58 14 62
rect 18 58 22 62
rect 8 57 22 58
rect 18 36 22 57
rect 28 60 38 62
rect 28 58 42 60
rect 28 42 32 58
rect 36 51 42 53
rect 40 47 42 51
rect 36 46 42 47
rect 26 41 32 42
rect 30 37 32 41
rect 26 36 32 37
rect 16 35 22 36
rect 4 32 8 33
rect 4 22 8 28
rect 20 31 22 35
rect 16 27 22 31
rect 20 23 22 27
rect 16 22 22 23
rect 28 32 32 36
rect 28 24 32 28
rect 38 32 42 46
rect 48 42 52 63
rect 58 51 62 68
rect 58 46 62 47
rect 52 38 63 42
rect 48 37 63 38
rect 62 32 66 33
rect 38 27 53 32
rect 62 24 66 28
rect 28 19 32 20
rect 39 18 40 22
rect 44 20 62 22
rect 44 18 66 20
rect 4 12 8 18
rect -2 8 72 12
rect -2 4 8 8
rect 12 4 18 8
rect 22 4 52 8
rect 56 4 72 8
rect -2 0 72 4
<< ntransistor >>
rect 11 17 13 36
rect 35 16 37 33
rect 47 16 49 33
rect 57 16 59 33
<< ptransistor >>
rect 21 55 23 93
rect 33 55 35 75
rect 45 55 47 93
rect 53 55 55 93
<< polycontact >>
rect 36 47 40 51
rect 26 37 30 41
rect 58 47 62 51
rect 48 38 52 42
<< ndcontact >>
rect 4 28 8 32
rect 4 18 8 22
rect 16 31 20 35
rect 16 23 20 27
rect 28 28 32 32
rect 28 20 32 24
rect 40 18 44 22
rect 62 28 66 32
rect 62 20 66 24
rect 52 4 56 8
<< pdcontact >>
rect 14 66 18 70
rect 14 58 18 62
rect 26 88 30 92
rect 26 78 30 82
rect 26 68 30 72
rect 38 68 42 72
rect 38 60 42 64
rect 58 88 62 92
rect 58 78 62 82
<< psubstratepcontact >>
rect 8 4 12 8
rect 18 4 22 8
<< nsubstratencontact >>
rect 4 92 8 96
<< psubstratepdiff >>
rect 7 8 23 9
rect 7 4 8 8
rect 12 4 18 8
rect 22 4 23 8
rect 7 3 23 4
<< nsubstratendiff >>
rect 3 96 9 97
rect 3 92 4 96
rect 8 92 9 96
rect 3 91 9 92
<< labels >>
rlabel polycontact 28 39 28 39 6 zn
rlabel metal1 20 45 20 45 6 z
rlabel metal1 10 60 10 60 6 z
rlabel metal1 35 6 35 6 6 vss
rlabel polycontact 29 39 29 39 6 zn
rlabel metal1 30 40 30 40 6 zn
rlabel metal1 35 94 35 94 6 vdd
rlabel metal1 50 30 50 30 6 b
rlabel metal1 40 40 40 40 6 b
rlabel metal1 50 50 50 50 6 a2
rlabel metal1 40 65 40 65 6 zn
rlabel metal1 50 70 50 70 6 a1
rlabel metal1 64 25 64 25 6 n2
rlabel metal1 52 20 52 20 6 n2
rlabel metal1 60 40 60 40 6 a2
rlabel metal1 60 60 60 60 6 a1
<< end >>
