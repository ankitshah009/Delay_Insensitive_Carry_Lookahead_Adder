magic
tech scmos
timestamp 1179386124
<< checkpaint >>
rect -22 -25 166 105
<< ab >>
rect 0 0 144 80
<< pwell >>
rect -4 -7 148 36
<< nwell >>
rect -4 36 148 87
<< polysilicon >>
rect 89 72 135 74
rect 19 66 21 71
rect 29 66 31 71
rect 89 69 91 72
rect 39 67 61 69
rect 9 60 11 65
rect 39 64 41 67
rect 49 64 51 67
rect 59 64 61 67
rect 69 67 91 69
rect 69 64 71 67
rect 79 64 81 67
rect 89 64 91 67
rect 99 64 101 68
rect 113 64 115 68
rect 123 64 125 68
rect 133 66 135 72
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 9 38 31 39
rect 39 38 41 42
rect 49 38 51 42
rect 59 39 61 42
rect 55 38 61 39
rect 69 38 71 42
rect 79 38 81 42
rect 89 38 91 42
rect 99 39 101 42
rect 113 39 115 42
rect 123 39 125 42
rect 133 39 135 42
rect 99 38 125 39
rect 9 34 10 38
rect 14 34 18 38
rect 22 34 31 38
rect 55 34 56 38
rect 60 34 61 38
rect 99 34 106 38
rect 110 34 114 38
rect 118 34 125 38
rect 9 33 31 34
rect 9 30 11 33
rect 19 30 21 33
rect 29 30 31 33
rect 39 30 41 34
rect 49 30 51 34
rect 55 32 91 34
rect 9 15 11 19
rect 19 14 21 19
rect 29 14 31 19
rect 39 9 41 15
rect 69 29 71 32
rect 79 29 81 32
rect 89 29 91 32
rect 99 33 125 34
rect 129 38 135 39
rect 129 34 130 38
rect 134 34 135 38
rect 129 33 135 34
rect 99 29 101 33
rect 111 29 113 33
rect 121 29 123 33
rect 133 29 135 33
rect 69 13 71 18
rect 79 13 81 18
rect 89 13 91 18
rect 99 13 101 18
rect 111 13 113 18
rect 121 13 123 18
rect 49 9 51 12
rect 133 9 135 14
rect 39 7 135 9
<< ndiffusion >>
rect 2 24 9 30
rect 2 20 3 24
rect 7 20 9 24
rect 2 19 9 20
rect 11 29 19 30
rect 11 25 13 29
rect 17 25 19 29
rect 11 19 19 25
rect 21 24 29 30
rect 21 20 23 24
rect 27 20 29 24
rect 21 19 29 20
rect 31 29 39 30
rect 31 25 33 29
rect 37 25 39 29
rect 31 19 39 25
rect 34 15 39 19
rect 41 29 49 30
rect 41 25 43 29
rect 47 25 49 29
rect 41 15 49 25
rect 44 12 49 15
rect 51 22 56 30
rect 62 28 69 29
rect 62 24 63 28
rect 67 24 69 28
rect 62 23 69 24
rect 51 21 58 22
rect 51 17 53 21
rect 57 17 58 21
rect 64 18 69 23
rect 71 23 79 29
rect 71 19 73 23
rect 77 19 79 23
rect 71 18 79 19
rect 81 28 89 29
rect 81 24 83 28
rect 87 24 89 28
rect 81 18 89 24
rect 91 28 99 29
rect 91 24 93 28
rect 97 24 99 28
rect 91 18 99 24
rect 101 18 111 29
rect 113 23 121 29
rect 113 19 115 23
rect 119 19 121 23
rect 113 18 121 19
rect 123 23 133 29
rect 123 19 126 23
rect 130 19 133 23
rect 123 18 133 19
rect 51 16 58 17
rect 51 12 56 16
rect 103 16 109 18
rect 103 12 104 16
rect 108 12 109 16
rect 125 14 133 18
rect 135 28 142 29
rect 135 24 137 28
rect 141 24 142 28
rect 135 23 142 24
rect 135 14 140 23
rect 103 11 109 12
<< pdiffusion >>
rect 14 60 19 66
rect 2 59 9 60
rect 2 55 3 59
rect 7 55 9 59
rect 2 42 9 55
rect 11 54 19 60
rect 11 50 13 54
rect 17 50 19 54
rect 11 47 19 50
rect 11 43 13 47
rect 17 43 19 47
rect 11 42 19 43
rect 21 65 29 66
rect 21 61 23 65
rect 27 61 29 65
rect 21 57 29 61
rect 21 53 23 57
rect 27 53 29 57
rect 21 42 29 53
rect 31 64 36 66
rect 127 64 133 66
rect 31 62 39 64
rect 31 58 33 62
rect 37 58 39 62
rect 31 54 39 58
rect 31 50 33 54
rect 37 50 39 54
rect 31 47 39 50
rect 31 43 33 47
rect 37 43 39 47
rect 31 42 39 43
rect 41 54 49 64
rect 41 50 43 54
rect 47 50 49 54
rect 41 47 49 50
rect 41 43 43 47
rect 47 43 49 47
rect 41 42 49 43
rect 51 63 59 64
rect 51 59 53 63
rect 57 59 59 63
rect 51 42 59 59
rect 61 47 69 64
rect 61 43 63 47
rect 67 43 69 47
rect 61 42 69 43
rect 71 54 79 64
rect 71 50 73 54
rect 77 50 79 54
rect 71 47 79 50
rect 71 43 73 47
rect 77 43 79 47
rect 71 42 79 43
rect 81 47 89 64
rect 81 43 83 47
rect 87 43 89 47
rect 81 42 89 43
rect 91 54 99 64
rect 91 50 93 54
rect 97 50 99 54
rect 91 47 99 50
rect 91 43 93 47
rect 97 43 99 47
rect 91 42 99 43
rect 101 63 113 64
rect 101 59 107 63
rect 111 59 113 63
rect 101 42 113 59
rect 115 47 123 64
rect 115 43 117 47
rect 121 43 123 47
rect 115 42 123 43
rect 125 63 133 64
rect 125 59 127 63
rect 131 59 133 63
rect 125 42 133 59
rect 135 55 140 66
rect 135 54 142 55
rect 135 50 137 54
rect 141 50 142 54
rect 135 47 142 50
rect 135 43 137 47
rect 141 43 142 47
rect 135 42 142 43
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect 118 78 122 82
rect 126 78 130 82
rect 134 78 138 82
rect 142 78 146 82
rect -2 68 146 78
rect 3 59 7 68
rect 23 65 27 68
rect 107 63 111 68
rect 23 57 27 61
rect 3 54 7 55
rect 13 54 17 55
rect 23 52 27 53
rect 33 62 53 63
rect 37 59 53 62
rect 57 59 58 63
rect 63 59 104 63
rect 33 54 37 58
rect 63 55 67 59
rect 100 55 104 59
rect 126 63 132 68
rect 126 59 127 63
rect 131 59 132 63
rect 107 58 111 59
rect 13 47 17 50
rect 2 38 6 47
rect 33 47 37 50
rect 17 43 33 46
rect 13 42 37 43
rect 2 34 10 38
rect 14 34 18 38
rect 22 34 23 38
rect 2 33 6 34
rect 33 31 37 42
rect 13 29 37 31
rect 17 27 33 29
rect 3 24 7 25
rect 13 24 17 25
rect 3 12 7 20
rect 22 20 23 24
rect 27 20 28 24
rect 22 12 28 20
rect 33 21 37 25
rect 42 54 47 55
rect 42 50 43 54
rect 42 47 47 50
rect 42 43 43 47
rect 42 30 47 43
rect 56 51 67 55
rect 73 54 97 55
rect 56 38 60 51
rect 77 51 93 54
rect 56 33 60 34
rect 63 47 67 48
rect 63 30 67 43
rect 73 47 77 50
rect 92 50 93 51
rect 100 54 142 55
rect 100 51 137 54
rect 73 42 77 43
rect 82 47 87 48
rect 82 43 83 47
rect 92 47 97 50
rect 141 50 142 54
rect 137 47 142 50
rect 92 43 93 47
rect 97 43 117 47
rect 121 43 122 47
rect 82 30 87 43
rect 42 29 88 30
rect 42 25 43 29
rect 47 28 88 29
rect 47 26 63 28
rect 42 24 47 25
rect 67 26 83 28
rect 82 24 83 26
rect 87 24 88 28
rect 93 28 97 43
rect 130 38 134 47
rect 141 43 142 47
rect 137 42 142 43
rect 105 34 106 38
rect 110 34 114 38
rect 118 34 119 38
rect 105 26 111 34
rect 130 30 134 34
rect 121 26 134 30
rect 138 29 142 42
rect 137 28 142 29
rect 63 23 67 24
rect 93 23 97 24
rect 141 24 142 28
rect 137 23 142 24
rect 33 17 53 21
rect 57 17 58 21
rect 72 19 73 23
rect 77 21 78 23
rect 93 21 115 23
rect 77 19 115 21
rect 119 19 120 23
rect 125 19 126 23
rect 130 19 131 23
rect 72 17 97 19
rect 103 12 104 16
rect 108 12 109 16
rect 125 12 131 19
rect -2 2 146 12
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 122 2
rect 126 -2 130 2
rect 134 -2 138 2
rect 142 -2 146 2
<< ntransistor >>
rect 9 19 11 30
rect 19 19 21 30
rect 29 19 31 30
rect 39 15 41 30
rect 49 12 51 30
rect 69 18 71 29
rect 79 18 81 29
rect 89 18 91 29
rect 99 18 101 29
rect 111 18 113 29
rect 121 18 123 29
rect 133 14 135 29
<< ptransistor >>
rect 9 42 11 60
rect 19 42 21 66
rect 29 42 31 66
rect 39 42 41 64
rect 49 42 51 64
rect 59 42 61 64
rect 69 42 71 64
rect 79 42 81 64
rect 89 42 91 64
rect 99 42 101 64
rect 113 42 115 64
rect 123 42 125 64
rect 133 42 135 66
<< polycontact >>
rect 10 34 14 38
rect 18 34 22 38
rect 56 34 60 38
rect 106 34 110 38
rect 114 34 118 38
rect 130 34 134 38
<< ndcontact >>
rect 3 20 7 24
rect 13 25 17 29
rect 23 20 27 24
rect 33 25 37 29
rect 43 25 47 29
rect 63 24 67 28
rect 53 17 57 21
rect 73 19 77 23
rect 83 24 87 28
rect 93 24 97 28
rect 115 19 119 23
rect 126 19 130 23
rect 104 12 108 16
rect 137 24 141 28
<< pdcontact >>
rect 3 55 7 59
rect 13 50 17 54
rect 13 43 17 47
rect 23 61 27 65
rect 23 53 27 57
rect 33 58 37 62
rect 33 50 37 54
rect 33 43 37 47
rect 43 50 47 54
rect 43 43 47 47
rect 53 59 57 63
rect 63 43 67 47
rect 73 50 77 54
rect 73 43 77 47
rect 83 43 87 47
rect 93 50 97 54
rect 93 43 97 47
rect 107 59 111 63
rect 117 43 121 47
rect 127 59 131 63
rect 137 50 141 54
rect 137 43 141 47
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
rect 90 -2 94 2
rect 98 -2 102 2
rect 106 -2 110 2
rect 114 -2 118 2
rect 122 -2 126 2
rect 130 -2 134 2
rect 138 -2 142 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
rect 90 78 94 82
rect 98 78 102 82
rect 106 78 110 82
rect 114 78 118 82
rect 122 78 126 82
rect 130 78 134 82
rect 138 78 142 82
<< psubstratepdiff >>
rect 0 2 144 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 122 2
rect 126 -2 130 2
rect 134 -2 138 2
rect 142 -2 144 2
rect 0 -3 144 -2
<< nsubstratendiff >>
rect 0 82 144 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect 118 78 122 82
rect 126 78 130 82
rect 134 78 138 82
rect 142 78 144 82
rect 0 77 144 78
<< labels >>
rlabel polycontact 58 35 58 35 6 sn
rlabel metal1 4 40 4 40 6 a1
rlabel polycontact 12 36 12 36 6 a1
rlabel polycontact 20 36 20 36 6 a1
rlabel metal1 15 48 15 48 6 a1n
rlabel metal1 52 28 52 28 6 z
rlabel metal1 25 29 25 29 6 a1n
rlabel metal1 44 40 44 40 6 z
rlabel metal1 35 40 35 40 6 a1n
rlabel metal1 72 6 72 6 6 vss
rlabel metal1 60 28 60 28 6 z
rlabel metal1 45 19 45 19 6 a1n
rlabel metal1 76 28 76 28 6 z
rlabel metal1 68 28 68 28 6 z
rlabel metal1 84 36 84 36 6 z
rlabel metal1 75 48 75 48 6 a0n
rlabel metal1 58 44 58 44 6 sn
rlabel metal1 45 61 45 61 6 a1n
rlabel metal1 72 74 72 74 6 vdd
rlabel metal1 84 19 84 19 6 a0n
rlabel metal1 108 32 108 32 6 a0
rlabel metal1 95 36 95 36 6 a0n
rlabel metal1 106 21 106 21 6 a0n
rlabel metal1 124 28 124 28 6 s
rlabel polycontact 116 36 116 36 6 a0
rlabel metal1 107 45 107 45 6 a0n
rlabel metal1 132 40 132 40 6 s
rlabel metal1 140 39 140 39 6 sn
<< end >>
