magic
tech scmos
timestamp 1179387107
<< checkpaint >>
rect -22 -25 78 105
<< ab >>
rect 0 0 56 80
<< pwell >>
rect -4 -7 60 36
<< nwell >>
rect -4 36 60 87
<< polysilicon >>
rect 23 70 25 74
rect 30 70 32 74
rect 37 70 39 74
rect 13 61 15 66
rect 13 39 15 50
rect 23 40 25 43
rect 9 38 15 39
rect 9 34 10 38
rect 14 34 15 38
rect 9 33 15 34
rect 19 39 26 40
rect 19 35 21 39
rect 25 35 26 39
rect 19 34 26 35
rect 9 23 11 33
rect 19 23 21 34
rect 30 32 32 43
rect 37 40 39 43
rect 37 39 47 40
rect 37 38 42 39
rect 41 35 42 38
rect 46 35 47 39
rect 41 34 47 35
rect 30 31 37 32
rect 30 27 32 31
rect 36 27 37 31
rect 30 26 37 27
rect 31 23 33 26
rect 41 23 43 34
rect 9 9 11 14
rect 19 9 21 14
rect 31 9 33 14
rect 41 9 43 14
<< ndiffusion >>
rect 2 22 9 23
rect 2 18 3 22
rect 7 18 9 22
rect 2 17 9 18
rect 4 14 9 17
rect 11 21 19 23
rect 11 17 13 21
rect 17 17 19 21
rect 11 14 19 17
rect 21 14 31 23
rect 33 21 41 23
rect 33 17 35 21
rect 39 17 41 21
rect 33 14 41 17
rect 43 19 50 23
rect 43 15 45 19
rect 49 15 50 19
rect 43 14 50 15
rect 23 12 29 14
rect 23 8 24 12
rect 28 8 29 12
rect 23 7 29 8
<< pdiffusion >>
rect 5 62 11 63
rect 5 58 6 62
rect 10 61 11 62
rect 18 61 23 70
rect 10 58 13 61
rect 5 50 13 58
rect 15 55 23 61
rect 15 51 17 55
rect 21 51 23 55
rect 15 50 23 51
rect 18 43 23 50
rect 25 43 30 70
rect 32 43 37 70
rect 39 69 48 70
rect 39 65 42 69
rect 46 65 48 69
rect 39 62 48 65
rect 39 58 42 62
rect 46 58 48 62
rect 39 43 48 58
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect -2 69 58 78
rect -2 68 42 69
rect 5 62 11 68
rect 41 65 42 68
rect 46 68 58 69
rect 46 65 47 68
rect 5 58 6 62
rect 10 58 11 62
rect 2 51 17 55
rect 21 51 22 55
rect 2 49 14 51
rect 2 23 6 49
rect 26 47 30 63
rect 41 62 47 65
rect 41 58 42 62
rect 46 58 47 62
rect 34 49 47 55
rect 18 41 30 47
rect 20 39 26 41
rect 42 39 47 49
rect 10 38 14 39
rect 20 35 21 39
rect 25 35 26 39
rect 10 30 14 34
rect 34 32 38 39
rect 46 35 47 39
rect 42 34 47 35
rect 32 31 38 32
rect 10 26 23 30
rect 36 30 38 31
rect 36 27 47 30
rect 32 26 47 27
rect 34 25 47 26
rect 2 22 7 23
rect 2 18 3 22
rect 2 17 7 18
rect 12 17 13 21
rect 17 17 35 21
rect 39 17 40 21
rect 45 19 49 20
rect 45 12 49 15
rect -2 8 24 12
rect 28 8 58 12
rect -2 2 58 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
<< ntransistor >>
rect 9 14 11 23
rect 19 14 21 23
rect 31 14 33 23
rect 41 14 43 23
<< ptransistor >>
rect 13 50 15 61
rect 23 43 25 70
rect 30 43 32 70
rect 37 43 39 70
<< polycontact >>
rect 10 34 14 38
rect 21 35 25 39
rect 42 35 46 39
rect 32 27 36 31
<< ndcontact >>
rect 3 18 7 22
rect 13 17 17 21
rect 35 17 39 21
rect 45 15 49 19
rect 24 8 28 12
<< pdcontact >>
rect 6 58 10 62
rect 17 51 21 55
rect 42 65 46 69
rect 42 58 46 62
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
<< psubstratepdiff >>
rect 0 2 56 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 56 2
rect 0 -3 56 -2
<< nsubstratendiff >>
rect 0 82 56 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 56 82
rect 0 77 56 78
<< labels >>
rlabel metal1 4 36 4 36 6 z
rlabel polycontact 12 36 12 36 6 b
rlabel metal1 20 28 20 28 6 b
rlabel metal1 20 44 20 44 6 a3
rlabel metal1 12 52 12 52 6 z
rlabel metal1 28 6 28 6 6 vss
rlabel metal1 26 19 26 19 6 n3
rlabel metal1 36 32 36 32 6 a2
rlabel metal1 28 52 28 52 6 a3
rlabel metal1 36 52 36 52 6 a1
rlabel metal1 28 74 28 74 6 vdd
rlabel metal1 44 28 44 28 6 a2
rlabel metal1 44 48 44 48 6 a1
<< end >>
