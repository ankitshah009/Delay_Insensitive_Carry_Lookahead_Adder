magic
tech scmos
timestamp 1179387230
<< checkpaint >>
rect -22 -25 94 105
<< ab >>
rect 0 0 72 80
<< pwell >>
rect -4 -7 76 36
<< nwell >>
rect -4 36 76 87
<< polysilicon >>
rect 9 70 11 74
rect 29 72 55 74
rect 22 64 24 69
rect 29 64 31 72
rect 36 64 38 68
rect 46 61 48 66
rect 53 61 55 72
rect 60 61 62 65
rect 9 39 11 42
rect 22 39 24 42
rect 9 38 15 39
rect 9 34 10 38
rect 14 34 15 38
rect 9 33 15 34
rect 19 38 25 39
rect 19 34 20 38
rect 24 34 25 38
rect 19 33 25 34
rect 9 30 11 33
rect 20 22 22 33
rect 29 31 31 42
rect 36 39 38 42
rect 46 39 48 42
rect 36 37 48 39
rect 53 37 55 42
rect 60 39 62 42
rect 60 38 67 39
rect 44 31 48 37
rect 60 34 62 38
rect 66 34 67 38
rect 60 33 67 34
rect 29 30 39 31
rect 29 26 34 30
rect 38 26 39 30
rect 29 25 39 26
rect 44 30 50 31
rect 44 26 45 30
rect 49 26 50 30
rect 44 25 50 26
rect 30 22 32 25
rect 44 22 46 25
rect 9 11 11 16
rect 20 9 22 14
rect 30 9 32 14
rect 44 9 46 14
<< ndiffusion >>
rect 2 29 9 30
rect 2 25 3 29
rect 7 25 9 29
rect 2 22 9 25
rect 2 18 3 22
rect 7 18 9 22
rect 2 16 9 18
rect 11 22 18 30
rect 11 20 20 22
rect 11 16 14 20
rect 18 16 20 20
rect 13 14 20 16
rect 22 21 30 22
rect 22 17 24 21
rect 28 17 30 21
rect 22 14 30 17
rect 32 14 44 22
rect 46 21 53 22
rect 46 17 48 21
rect 52 17 53 21
rect 46 16 53 17
rect 46 14 51 16
rect 34 12 42 14
rect 34 8 36 12
rect 40 8 42 12
rect 34 7 42 8
<< pdiffusion >>
rect 4 55 9 70
rect 2 54 9 55
rect 2 50 3 54
rect 7 50 9 54
rect 2 47 9 50
rect 2 43 3 47
rect 7 43 9 47
rect 2 42 9 43
rect 11 69 20 70
rect 11 65 15 69
rect 19 65 20 69
rect 11 64 20 65
rect 11 62 22 64
rect 11 58 15 62
rect 19 58 22 62
rect 11 42 22 58
rect 24 42 29 64
rect 31 42 36 64
rect 38 61 43 64
rect 38 60 46 61
rect 38 56 40 60
rect 44 56 46 60
rect 38 53 46 56
rect 38 49 40 53
rect 44 49 46 53
rect 38 42 46 49
rect 48 42 53 61
rect 55 42 60 61
rect 62 60 70 61
rect 62 56 64 60
rect 68 56 70 60
rect 62 53 70 56
rect 62 49 64 53
rect 68 49 70 53
rect 62 42 70 49
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect -2 69 74 78
rect -2 68 15 69
rect 14 65 15 68
rect 19 68 74 69
rect 19 65 20 68
rect 14 62 20 65
rect 14 58 15 62
rect 19 58 20 62
rect 63 60 69 68
rect 39 56 40 60
rect 44 56 45 60
rect 2 54 14 55
rect 2 50 3 54
rect 7 50 14 54
rect 39 53 45 56
rect 2 49 14 50
rect 18 49 40 53
rect 44 49 45 53
rect 63 56 64 60
rect 68 56 69 60
rect 63 53 69 56
rect 63 49 64 53
rect 68 49 69 53
rect 2 47 7 49
rect 2 43 3 47
rect 18 46 22 49
rect 2 42 7 43
rect 10 42 22 46
rect 26 42 63 46
rect 2 30 6 42
rect 10 38 14 42
rect 26 39 30 42
rect 2 29 7 30
rect 2 25 3 29
rect 10 29 14 34
rect 20 38 30 39
rect 57 38 63 42
rect 24 34 30 38
rect 20 33 30 34
rect 34 34 47 38
rect 57 34 62 38
rect 66 34 67 38
rect 34 30 38 34
rect 10 25 27 29
rect 44 26 45 30
rect 49 26 63 30
rect 34 25 38 26
rect 2 22 7 25
rect 2 18 3 22
rect 23 21 27 25
rect 2 17 7 18
rect 13 16 14 20
rect 18 16 19 20
rect 23 17 24 21
rect 28 17 48 21
rect 52 17 53 21
rect 57 18 63 26
rect 13 12 19 16
rect -2 8 36 12
rect 40 8 74 12
rect -2 2 74 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
<< ntransistor >>
rect 9 16 11 30
rect 20 14 22 22
rect 30 14 32 22
rect 44 14 46 22
<< ptransistor >>
rect 9 42 11 70
rect 22 42 24 64
rect 29 42 31 64
rect 36 42 38 64
rect 46 42 48 61
rect 53 42 55 61
rect 60 42 62 61
<< polycontact >>
rect 10 34 14 38
rect 20 34 24 38
rect 62 34 66 38
rect 34 26 38 30
rect 45 26 49 30
<< ndcontact >>
rect 3 25 7 29
rect 3 18 7 22
rect 14 16 18 20
rect 24 17 28 21
rect 48 17 52 21
rect 36 8 40 12
<< pdcontact >>
rect 3 50 7 54
rect 3 43 7 47
rect 15 65 19 69
rect 15 58 19 62
rect 40 56 44 60
rect 40 49 44 53
rect 64 56 68 60
rect 64 49 68 53
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
<< psubstratepdiff >>
rect 0 2 72 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 72 2
rect 0 -3 72 -2
<< nsubstratendiff >>
rect 0 82 72 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 72 82
rect 0 77 72 78
<< labels >>
rlabel polycontact 12 36 12 36 6 zn
rlabel metal1 4 36 4 36 6 z
rlabel polycontact 12 35 12 35 6 zn
rlabel metal1 12 52 12 52 6 z
rlabel metal1 36 6 36 6 6 vss
rlabel polycontact 36 28 36 28 6 b
rlabel metal1 28 36 28 36 6 a
rlabel metal1 36 44 36 44 6 a
rlabel metal1 36 74 36 74 6 vdd
rlabel metal1 38 19 38 19 6 zn
rlabel metal1 52 28 52 28 6 c
rlabel metal1 44 36 44 36 6 b
rlabel metal1 44 44 44 44 6 a
rlabel metal1 52 44 52 44 6 a
rlabel metal1 42 54 42 54 6 zn
rlabel metal1 31 51 31 51 6 zn
rlabel metal1 60 24 60 24 6 c
rlabel metal1 60 40 60 40 6 a
<< end >>
