magic
tech scmos
timestamp 1179387670
<< checkpaint >>
rect -22 -22 262 94
<< ab >>
rect 0 0 240 72
<< pwell >>
rect -4 -4 244 32
<< nwell >>
rect -4 32 244 76
<< polysilicon >>
rect 9 65 11 70
rect 19 65 21 70
rect 29 65 31 70
rect 39 65 41 70
rect 49 65 51 70
rect 59 65 61 70
rect 79 68 91 70
rect 79 65 81 68
rect 89 65 91 68
rect 119 65 121 70
rect 129 65 131 70
rect 139 65 141 70
rect 149 65 151 70
rect 159 65 161 70
rect 169 65 171 70
rect 179 65 181 70
rect 189 65 191 70
rect 199 65 201 70
rect 209 65 211 70
rect 219 65 221 70
rect 99 52 101 57
rect 109 52 111 57
rect 9 35 11 38
rect 19 35 21 38
rect 29 35 31 38
rect 39 35 41 38
rect 49 35 51 38
rect 59 35 61 38
rect 9 34 61 35
rect 79 34 81 38
rect 89 35 91 38
rect 99 35 101 38
rect 109 35 111 38
rect 119 35 121 38
rect 129 35 131 38
rect 139 35 141 38
rect 149 35 151 38
rect 85 34 91 35
rect 9 30 10 34
rect 14 30 61 34
rect 9 29 61 30
rect 9 26 11 29
rect 19 26 21 29
rect 29 26 31 29
rect 59 26 61 29
rect 69 26 71 31
rect 85 30 86 34
rect 90 30 91 34
rect 79 26 81 30
rect 85 29 91 30
rect 95 34 115 35
rect 95 30 96 34
rect 100 30 110 34
rect 114 30 115 34
rect 95 29 115 30
rect 119 34 131 35
rect 119 30 123 34
rect 127 30 131 34
rect 119 29 131 30
rect 135 34 151 35
rect 135 30 136 34
rect 140 33 151 34
rect 140 30 141 33
rect 135 29 141 30
rect 159 31 161 38
rect 169 35 171 38
rect 169 34 175 35
rect 169 31 170 34
rect 159 30 170 31
rect 174 30 175 34
rect 159 29 175 30
rect 89 26 91 29
rect 96 26 98 29
rect 112 26 114 29
rect 119 26 121 29
rect 129 26 131 29
rect 136 26 138 29
rect 152 28 161 29
rect 9 3 11 8
rect 19 3 21 8
rect 29 3 31 8
rect 59 5 61 8
rect 69 5 71 8
rect 79 5 81 8
rect 152 24 153 28
rect 157 24 161 28
rect 172 26 174 29
rect 179 26 181 38
rect 189 35 191 38
rect 199 35 201 38
rect 209 35 211 38
rect 219 35 221 38
rect 189 34 231 35
rect 189 30 226 34
rect 230 30 231 34
rect 189 29 231 30
rect 189 26 191 29
rect 199 26 201 29
rect 209 26 211 29
rect 152 23 161 24
rect 59 3 81 5
rect 89 2 91 6
rect 96 2 98 6
rect 112 2 114 6
rect 119 2 121 6
rect 129 3 131 8
rect 136 4 138 8
rect 172 8 174 12
rect 179 4 181 12
rect 136 2 181 4
rect 189 3 191 8
rect 199 3 201 8
rect 209 3 211 8
<< ndiffusion >>
rect 2 21 9 26
rect 2 17 3 21
rect 7 17 9 21
rect 2 13 9 17
rect 2 9 3 13
rect 7 9 9 13
rect 2 8 9 9
rect 11 25 19 26
rect 11 21 13 25
rect 17 21 19 25
rect 11 18 19 21
rect 11 14 13 18
rect 17 14 19 18
rect 11 8 19 14
rect 21 13 29 26
rect 21 9 23 13
rect 27 9 29 13
rect 21 8 29 9
rect 31 25 38 26
rect 31 21 33 25
rect 37 21 38 25
rect 52 25 59 26
rect 31 18 38 21
rect 31 14 33 18
rect 37 14 38 18
rect 31 13 38 14
rect 31 8 36 13
rect 52 21 53 25
rect 57 21 59 25
rect 52 18 59 21
rect 52 14 53 18
rect 57 14 59 18
rect 52 13 59 14
rect 54 8 59 13
rect 61 18 69 26
rect 61 14 63 18
rect 67 14 69 18
rect 61 8 69 14
rect 71 25 79 26
rect 71 21 73 25
rect 77 21 79 25
rect 71 8 79 21
rect 81 18 89 26
rect 81 14 83 18
rect 87 14 89 18
rect 81 8 89 14
rect 84 6 89 8
rect 91 6 96 26
rect 98 11 112 26
rect 98 7 103 11
rect 107 7 112 11
rect 98 6 112 7
rect 114 6 119 26
rect 121 18 129 26
rect 121 14 123 18
rect 127 14 129 18
rect 121 8 129 14
rect 131 8 136 26
rect 138 11 147 26
rect 165 25 172 26
rect 165 21 166 25
rect 170 21 172 25
rect 165 20 172 21
rect 138 8 141 11
rect 121 6 126 8
rect 140 7 141 8
rect 145 7 147 11
rect 140 6 147 7
rect 167 12 172 20
rect 174 12 179 26
rect 181 24 189 26
rect 181 20 183 24
rect 187 20 189 24
rect 181 17 189 20
rect 181 13 183 17
rect 187 13 189 17
rect 181 12 189 13
rect 184 8 189 12
rect 191 25 199 26
rect 191 21 193 25
rect 197 21 199 25
rect 191 18 199 21
rect 191 14 193 18
rect 197 14 199 18
rect 191 8 199 14
rect 201 21 209 26
rect 201 17 203 21
rect 207 17 209 21
rect 201 13 209 17
rect 201 9 203 13
rect 207 9 209 13
rect 201 8 209 9
rect 211 25 218 26
rect 211 21 213 25
rect 217 21 218 25
rect 211 18 218 21
rect 211 14 213 18
rect 217 14 218 18
rect 211 13 218 14
rect 211 8 216 13
<< pdiffusion >>
rect 2 64 9 65
rect 2 60 3 64
rect 7 60 9 64
rect 2 57 9 60
rect 2 53 3 57
rect 7 53 9 57
rect 2 38 9 53
rect 11 50 19 65
rect 11 46 13 50
rect 17 46 19 50
rect 11 43 19 46
rect 11 39 13 43
rect 17 39 19 43
rect 11 38 19 39
rect 21 64 29 65
rect 21 60 23 64
rect 27 60 29 64
rect 21 57 29 60
rect 21 53 23 57
rect 27 53 29 57
rect 21 38 29 53
rect 31 50 39 65
rect 31 46 33 50
rect 37 46 39 50
rect 31 43 39 46
rect 31 39 33 43
rect 37 39 39 43
rect 31 38 39 39
rect 41 64 49 65
rect 41 60 43 64
rect 47 60 49 64
rect 41 57 49 60
rect 41 53 43 57
rect 47 53 49 57
rect 41 38 49 53
rect 51 50 59 65
rect 51 46 53 50
rect 57 46 59 50
rect 51 43 59 46
rect 51 39 53 43
rect 57 39 59 43
rect 51 38 59 39
rect 61 64 68 65
rect 61 60 63 64
rect 67 60 68 64
rect 61 57 68 60
rect 74 58 79 65
rect 61 53 63 57
rect 67 53 68 57
rect 61 38 68 53
rect 72 57 79 58
rect 72 53 73 57
rect 77 53 79 57
rect 72 50 79 53
rect 72 46 73 50
rect 77 46 79 50
rect 72 45 79 46
rect 74 38 79 45
rect 81 50 89 65
rect 81 46 83 50
rect 87 46 89 50
rect 81 43 89 46
rect 81 39 83 43
rect 87 39 89 43
rect 81 38 89 39
rect 91 52 96 65
rect 114 52 119 65
rect 91 51 99 52
rect 91 47 93 51
rect 97 47 99 51
rect 91 38 99 47
rect 101 43 109 52
rect 101 39 103 43
rect 107 39 109 43
rect 101 38 109 39
rect 111 51 119 52
rect 111 47 113 51
rect 117 47 119 51
rect 111 38 119 47
rect 121 43 129 65
rect 121 39 123 43
rect 127 39 129 43
rect 121 38 129 39
rect 131 58 139 65
rect 131 54 133 58
rect 137 54 139 58
rect 131 38 139 54
rect 141 43 149 65
rect 141 39 143 43
rect 147 39 149 43
rect 141 38 149 39
rect 151 58 159 65
rect 151 54 153 58
rect 157 54 159 58
rect 151 38 159 54
rect 161 50 169 65
rect 161 46 163 50
rect 167 46 169 50
rect 161 38 169 46
rect 171 57 179 65
rect 171 53 173 57
rect 177 53 179 57
rect 171 50 179 53
rect 171 46 173 50
rect 177 46 179 50
rect 171 43 179 46
rect 171 39 173 43
rect 177 39 179 43
rect 171 38 179 39
rect 181 50 189 65
rect 181 46 183 50
rect 187 46 189 50
rect 181 43 189 46
rect 181 39 183 43
rect 187 39 189 43
rect 181 38 189 39
rect 191 64 199 65
rect 191 60 193 64
rect 197 60 199 64
rect 191 57 199 60
rect 191 53 193 57
rect 197 53 199 57
rect 191 38 199 53
rect 201 50 209 65
rect 201 46 203 50
rect 207 46 209 50
rect 201 43 209 46
rect 201 39 203 43
rect 207 39 209 43
rect 201 38 209 39
rect 211 64 219 65
rect 211 60 213 64
rect 217 60 219 64
rect 211 57 219 60
rect 211 53 213 57
rect 217 53 219 57
rect 211 38 219 53
rect 221 51 226 65
rect 221 50 228 51
rect 221 46 223 50
rect 227 46 228 50
rect 221 43 228 46
rect 221 39 223 43
rect 227 39 228 43
rect 221 38 228 39
<< metal1 >>
rect -2 68 242 72
rect -2 64 103 68
rect 107 64 232 68
rect 236 64 242 68
rect 3 57 7 60
rect 3 52 7 53
rect 23 57 27 60
rect 23 52 27 53
rect 43 57 47 60
rect 43 52 47 53
rect 63 57 67 60
rect 63 52 67 53
rect 73 57 133 58
rect 77 54 133 57
rect 137 54 153 58
rect 157 57 177 58
rect 157 54 173 57
rect 77 53 78 54
rect 13 50 17 51
rect 13 43 17 46
rect 2 34 6 43
rect 33 50 37 51
rect 33 43 37 46
rect 17 39 33 42
rect 53 50 57 51
rect 53 43 57 46
rect 73 50 78 53
rect 92 51 98 54
rect 77 46 78 50
rect 73 45 78 46
rect 83 50 87 51
rect 92 47 93 51
rect 97 47 98 51
rect 112 51 118 54
rect 112 47 113 51
rect 117 47 118 51
rect 173 50 177 53
rect 193 57 197 60
rect 193 52 197 53
rect 213 57 217 60
rect 213 52 217 53
rect 37 39 53 42
rect 83 43 87 46
rect 134 46 163 50
rect 167 46 168 50
rect 57 39 83 42
rect 103 43 107 44
rect 134 43 138 46
rect 173 43 177 46
rect 87 39 100 42
rect 13 38 100 39
rect 2 30 10 34
rect 14 30 15 34
rect 2 29 15 30
rect 33 25 37 38
rect 86 34 90 35
rect 86 26 90 30
rect 96 34 100 38
rect 96 29 100 30
rect 103 26 107 39
rect 110 39 123 43
rect 127 39 138 43
rect 142 39 143 43
rect 147 39 149 43
rect 110 34 114 39
rect 134 34 138 39
rect 110 29 114 30
rect 122 30 123 34
rect 127 30 128 34
rect 134 30 136 34
rect 140 30 141 34
rect 122 26 128 30
rect 145 28 149 39
rect 162 39 173 42
rect 162 38 177 39
rect 183 50 187 51
rect 183 43 187 46
rect 203 50 207 51
rect 203 43 207 46
rect 223 50 228 51
rect 227 46 228 50
rect 223 43 228 46
rect 187 39 203 43
rect 207 39 223 43
rect 227 39 228 43
rect 145 26 153 28
rect 3 21 7 22
rect 3 13 7 17
rect 12 21 13 25
rect 17 21 33 25
rect 12 18 17 21
rect 12 14 13 18
rect 33 18 37 21
rect 12 13 17 14
rect 23 13 27 14
rect 33 13 37 14
rect 53 25 153 26
rect 57 22 73 25
rect 72 21 73 22
rect 77 24 153 25
rect 157 24 158 28
rect 77 22 149 24
rect 77 21 78 22
rect 53 18 57 21
rect 162 18 166 38
rect 183 34 187 39
rect 169 30 170 34
rect 174 30 187 34
rect 193 25 197 39
rect 170 21 171 25
rect 183 24 187 25
rect 62 14 63 18
rect 67 14 83 18
rect 87 14 123 18
rect 127 14 166 18
rect 183 17 187 20
rect 53 13 57 14
rect 213 25 217 39
rect 226 34 238 35
rect 230 30 238 34
rect 226 29 238 30
rect 193 18 197 21
rect 193 13 197 14
rect 203 21 207 22
rect 203 13 207 17
rect 234 21 238 29
rect 213 18 217 21
rect 213 13 217 14
rect 3 8 7 9
rect 23 8 27 9
rect 102 8 103 11
rect -2 4 43 8
rect 47 7 103 8
rect 107 8 108 11
rect 140 8 141 11
rect 107 7 141 8
rect 145 8 146 11
rect 155 8 156 11
rect 145 7 156 8
rect 160 8 161 11
rect 183 8 187 13
rect 203 8 207 9
rect 160 7 232 8
rect 47 4 232 7
rect 236 4 242 8
rect -2 0 242 4
<< ntransistor >>
rect 9 8 11 26
rect 19 8 21 26
rect 29 8 31 26
rect 59 8 61 26
rect 69 8 71 26
rect 79 8 81 26
rect 89 6 91 26
rect 96 6 98 26
rect 112 6 114 26
rect 119 6 121 26
rect 129 8 131 26
rect 136 8 138 26
rect 172 12 174 26
rect 179 12 181 26
rect 189 8 191 26
rect 199 8 201 26
rect 209 8 211 26
<< ptransistor >>
rect 9 38 11 65
rect 19 38 21 65
rect 29 38 31 65
rect 39 38 41 65
rect 49 38 51 65
rect 59 38 61 65
rect 79 38 81 65
rect 89 38 91 65
rect 99 38 101 52
rect 109 38 111 52
rect 119 38 121 65
rect 129 38 131 65
rect 139 38 141 65
rect 149 38 151 65
rect 159 38 161 65
rect 169 38 171 65
rect 179 38 181 65
rect 189 38 191 65
rect 199 38 201 65
rect 209 38 211 65
rect 219 38 221 65
<< polycontact >>
rect 10 30 14 34
rect 86 30 90 34
rect 96 30 100 34
rect 110 30 114 34
rect 123 30 127 34
rect 136 30 140 34
rect 170 30 174 34
rect 153 24 157 28
rect 226 30 230 34
<< ndcontact >>
rect 3 17 7 21
rect 3 9 7 13
rect 13 21 17 25
rect 13 14 17 18
rect 23 9 27 13
rect 33 21 37 25
rect 33 14 37 18
rect 53 21 57 25
rect 53 14 57 18
rect 63 14 67 18
rect 73 21 77 25
rect 83 14 87 18
rect 103 7 107 11
rect 123 14 127 18
rect 166 21 170 25
rect 141 7 145 11
rect 183 20 187 24
rect 183 13 187 17
rect 193 21 197 25
rect 193 14 197 18
rect 203 17 207 21
rect 203 9 207 13
rect 213 21 217 25
rect 213 14 217 18
<< pdcontact >>
rect 3 60 7 64
rect 3 53 7 57
rect 13 46 17 50
rect 13 39 17 43
rect 23 60 27 64
rect 23 53 27 57
rect 33 46 37 50
rect 33 39 37 43
rect 43 60 47 64
rect 43 53 47 57
rect 53 46 57 50
rect 53 39 57 43
rect 63 60 67 64
rect 63 53 67 57
rect 73 53 77 57
rect 73 46 77 50
rect 83 46 87 50
rect 83 39 87 43
rect 93 47 97 51
rect 103 39 107 43
rect 113 47 117 51
rect 123 39 127 43
rect 133 54 137 58
rect 143 39 147 43
rect 153 54 157 58
rect 163 46 167 50
rect 173 53 177 57
rect 173 46 177 50
rect 173 39 177 43
rect 183 46 187 50
rect 183 39 187 43
rect 193 60 197 64
rect 193 53 197 57
rect 203 46 207 50
rect 203 39 207 43
rect 213 60 217 64
rect 213 53 217 57
rect 223 46 227 50
rect 223 39 227 43
<< psubstratepcontact >>
rect 43 4 47 8
rect 156 7 160 11
rect 232 4 236 8
<< nsubstratencontact >>
rect 103 64 107 68
rect 232 64 236 68
<< psubstratepdiff >>
rect 42 8 48 24
rect 42 4 43 8
rect 47 4 48 8
rect 42 3 48 4
rect 155 11 161 20
rect 155 7 156 11
rect 160 7 161 11
rect 155 6 161 7
rect 231 8 237 24
rect 231 4 232 8
rect 236 4 237 8
rect 231 3 237 4
<< nsubstratendiff >>
rect 100 68 110 69
rect 100 64 103 68
rect 107 64 110 68
rect 231 68 237 69
rect 100 63 110 64
rect 231 64 232 68
rect 236 64 237 68
rect 231 55 237 64
<< labels >>
rlabel polycontact 88 32 88 32 6 an
rlabel polysilicon 105 32 105 32 6 bn
rlabel polycontact 125 32 125 32 6 an
rlabel polycontact 138 32 138 32 6 bn
rlabel polycontact 156 26 156 26 6 an
rlabel polycontact 172 32 172 32 6 an
rlabel metal1 14 19 14 19 6 bn
rlabel polycontact 12 32 12 32 6 b
rlabel metal1 4 36 4 36 6 b
rlabel metal1 15 44 15 44 6 bn
rlabel metal1 35 32 35 32 6 bn
rlabel metal1 92 16 92 16 6 z
rlabel ndcontact 84 16 84 16 6 z
rlabel metal1 76 16 76 16 6 z
rlabel metal1 68 16 68 16 6 z
rlabel metal1 55 19 55 19 6 an
rlabel metal1 88 28 88 28 6 an
rlabel metal1 85 44 85 44 6 bn
rlabel metal1 55 44 55 44 6 bn
rlabel metal1 76 52 76 52 6 z
rlabel metal1 92 56 92 56 6 z
rlabel metal1 84 56 84 56 6 z
rlabel metal1 120 4 120 4 6 vss
rlabel metal1 100 16 100 16 6 z
rlabel metal1 108 16 108 16 6 z
rlabel metal1 116 16 116 16 6 z
rlabel ndcontact 124 16 124 16 6 z
rlabel metal1 132 16 132 16 6 z
rlabel metal1 140 16 140 16 6 z
rlabel metal1 125 28 125 28 6 an
rlabel metal1 98 35 98 35 6 bn
rlabel pdcontact 124 41 124 41 6 bn
rlabel metal1 112 36 112 36 6 bn
rlabel metal1 105 33 105 33 6 an
rlabel metal1 136 40 136 40 6 bn
rlabel metal1 140 56 140 56 6 z
rlabel metal1 132 56 132 56 6 z
rlabel metal1 124 56 124 56 6 z
rlabel metal1 116 56 116 56 6 z
rlabel metal1 108 56 108 56 6 z
rlabel metal1 100 56 100 56 6 z
rlabel metal1 120 68 120 68 6 vdd
rlabel metal1 156 16 156 16 6 z
rlabel metal1 148 16 148 16 6 z
rlabel metal1 101 24 101 24 6 an
rlabel metal1 164 28 164 28 6 z
rlabel metal1 178 32 178 32 6 an
rlabel metal1 151 26 151 26 6 an
rlabel metal1 172 40 172 40 6 z
rlabel pdcontact 145 41 145 41 6 an
rlabel metal1 151 48 151 48 6 bn
rlabel metal1 172 56 172 56 6 z
rlabel metal1 164 56 164 56 6 z
rlabel pdcontact 156 56 156 56 6 z
rlabel metal1 148 56 148 56 6 z
rlabel polycontact 228 32 228 32 6 a
rlabel metal1 236 28 236 28 6 a
rlabel metal1 205 45 205 45 6 an
rlabel metal1 225 45 225 45 6 an
rlabel pdcontact 205 41 205 41 6 an
rlabel metal1 215 28 215 28 6 an
rlabel metal1 195 28 195 28 6 an
<< end >>
