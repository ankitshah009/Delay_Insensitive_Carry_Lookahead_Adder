magic
tech scmos
timestamp 1179386065
<< checkpaint >>
rect -22 -25 78 105
<< ab >>
rect 0 0 56 80
<< pwell >>
rect -4 -7 60 36
<< nwell >>
rect -4 36 60 87
<< polysilicon >>
rect 9 66 11 71
rect 16 66 18 71
rect 26 66 28 71
rect 33 66 35 71
rect 45 63 51 64
rect 45 59 46 63
rect 50 59 51 63
rect 45 58 51 59
rect 45 55 47 58
rect 9 47 11 50
rect 2 46 11 47
rect 2 42 3 46
rect 7 45 11 46
rect 7 42 8 45
rect 2 41 8 42
rect 16 41 18 50
rect 26 47 28 50
rect 23 46 29 47
rect 23 42 24 46
rect 28 42 29 46
rect 23 41 29 42
rect 6 27 8 41
rect 12 40 18 41
rect 12 36 13 40
rect 17 37 18 40
rect 33 40 35 50
rect 45 46 47 49
rect 45 44 52 46
rect 33 39 46 40
rect 17 36 28 37
rect 12 35 28 36
rect 16 30 22 31
rect 6 25 11 27
rect 9 22 11 25
rect 16 26 17 30
rect 21 26 22 30
rect 16 25 22 26
rect 16 22 18 25
rect 26 22 28 35
rect 33 35 41 39
rect 45 35 46 39
rect 33 34 46 35
rect 33 22 35 34
rect 50 30 52 44
rect 45 28 52 30
rect 45 25 47 28
rect 45 15 47 19
rect 9 10 11 15
rect 16 10 18 15
rect 26 10 28 15
rect 33 10 35 15
<< ndiffusion >>
rect 37 22 45 25
rect 2 20 9 22
rect 2 16 3 20
rect 7 16 9 20
rect 2 15 9 16
rect 11 15 16 22
rect 18 21 26 22
rect 18 17 20 21
rect 24 17 26 21
rect 18 15 26 17
rect 28 15 33 22
rect 35 19 45 22
rect 47 24 54 25
rect 47 20 49 24
rect 53 20 54 24
rect 47 19 54 20
rect 35 15 43 19
rect 37 12 43 15
rect 37 8 38 12
rect 42 8 43 12
rect 37 7 43 8
<< pdiffusion >>
rect 37 72 43 73
rect 37 68 38 72
rect 42 68 43 72
rect 37 66 43 68
rect 2 65 9 66
rect 2 61 3 65
rect 7 61 9 65
rect 2 50 9 61
rect 11 50 16 66
rect 18 55 26 66
rect 18 51 20 55
rect 24 51 26 55
rect 18 50 26 51
rect 28 50 33 66
rect 35 55 43 66
rect 35 50 45 55
rect 37 49 45 50
rect 47 54 54 55
rect 47 50 49 54
rect 53 50 54 54
rect 47 49 54 50
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect -2 72 58 78
rect -2 68 38 72
rect 42 68 58 72
rect 3 65 7 68
rect 45 62 46 63
rect 3 60 7 61
rect 11 59 46 62
rect 50 59 51 63
rect 11 58 51 59
rect 11 55 15 58
rect 2 50 15 55
rect 19 51 20 55
rect 24 54 25 55
rect 49 54 53 55
rect 24 51 38 54
rect 19 50 38 51
rect 2 46 8 50
rect 2 42 3 46
rect 7 42 8 46
rect 23 42 24 46
rect 28 42 30 46
rect 12 38 13 40
rect 2 36 13 38
rect 17 36 18 40
rect 2 34 18 36
rect 2 25 6 34
rect 26 30 30 42
rect 16 26 17 30
rect 21 26 30 30
rect 34 22 38 50
rect 49 40 53 50
rect 41 39 53 40
rect 45 35 53 39
rect 41 34 53 35
rect 17 21 38 22
rect 3 20 7 21
rect 17 17 20 21
rect 24 17 38 21
rect 49 24 53 34
rect 49 19 53 20
rect 3 12 7 16
rect -2 8 38 12
rect 42 8 58 12
rect -2 2 58 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
<< ntransistor >>
rect 9 15 11 22
rect 16 15 18 22
rect 26 15 28 22
rect 33 15 35 22
rect 45 19 47 25
<< ptransistor >>
rect 9 50 11 66
rect 16 50 18 66
rect 26 50 28 66
rect 33 50 35 66
rect 45 49 47 55
<< polycontact >>
rect 46 59 50 63
rect 3 42 7 46
rect 24 42 28 46
rect 13 36 17 40
rect 17 26 21 30
rect 41 35 45 39
<< ndcontact >>
rect 3 16 7 20
rect 20 17 24 21
rect 49 20 53 24
rect 38 8 42 12
<< pdcontact >>
rect 38 68 42 72
rect 3 61 7 65
rect 20 51 24 55
rect 49 50 53 54
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
<< psubstratepdiff >>
rect 0 2 56 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 56 2
rect 0 -3 56 -2
<< nsubstratendiff >>
rect 0 82 56 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 56 82
rect 0 77 56 78
<< labels >>
rlabel polysilicon 39 37 39 37 6 sn
rlabel metal1 4 28 4 28 6 a0
rlabel metal1 4 52 4 52 6 s
rlabel metal1 12 36 12 36 6 a0
rlabel metal1 12 52 12 52 6 s
rlabel metal1 28 6 28 6 6 vss
rlabel polycontact 20 28 20 28 6 a1
rlabel metal1 20 20 20 20 6 z
rlabel metal1 28 20 28 20 6 z
rlabel metal1 28 36 28 36 6 a1
rlabel metal1 28 52 28 52 6 z
rlabel metal1 20 60 20 60 6 s
rlabel metal1 28 60 28 60 6 s
rlabel metal1 28 74 28 74 6 vdd
rlabel metal1 36 32 36 32 6 z
rlabel metal1 36 60 36 60 6 s
rlabel metal1 44 60 44 60 6 s
rlabel metal1 47 37 47 37 6 sn
rlabel metal1 51 37 51 37 6 sn
<< end >>
