magic
tech scmos
timestamp 1179385481
<< checkpaint >>
rect -22 -25 62 105
<< ab >>
rect 0 0 40 80
<< pwell >>
rect -4 -7 44 36
<< nwell >>
rect -4 36 44 87
<< polysilicon >>
rect 19 65 21 70
rect 29 65 31 70
rect 9 61 11 65
rect 9 39 11 43
rect 19 39 21 43
rect 9 38 21 39
rect 9 34 16 38
rect 20 34 21 38
rect 9 33 21 34
rect 9 30 11 33
rect 29 31 31 43
rect 25 30 31 31
rect 25 26 26 30
rect 30 26 31 30
rect 25 25 31 26
rect 29 22 31 25
rect 9 6 11 10
rect 29 6 31 10
<< ndiffusion >>
rect 2 29 9 30
rect 2 25 3 29
rect 7 25 9 29
rect 2 22 9 25
rect 2 18 3 22
rect 7 18 9 22
rect 2 17 9 18
rect 4 10 9 17
rect 11 22 22 30
rect 11 18 16 22
rect 20 18 29 22
rect 11 15 29 18
rect 11 11 16 15
rect 20 11 29 15
rect 11 10 29 11
rect 31 21 38 22
rect 31 17 33 21
rect 37 17 38 21
rect 31 16 38 17
rect 31 10 36 16
<< pdiffusion >>
rect 14 61 19 65
rect 2 60 9 61
rect 2 56 3 60
rect 7 56 9 60
rect 2 53 9 56
rect 2 49 3 53
rect 7 49 9 53
rect 2 43 9 49
rect 11 55 19 61
rect 11 51 13 55
rect 17 51 19 55
rect 11 48 19 51
rect 11 44 13 48
rect 17 44 19 48
rect 11 43 19 44
rect 21 64 29 65
rect 21 60 23 64
rect 27 60 29 64
rect 21 57 29 60
rect 21 53 23 57
rect 27 53 29 57
rect 21 43 29 53
rect 31 56 36 65
rect 31 55 38 56
rect 31 51 33 55
rect 37 51 38 55
rect 31 48 38 51
rect 31 44 33 48
rect 37 44 38 48
rect 31 43 38 44
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect -2 68 42 78
rect 2 60 8 68
rect 2 56 3 60
rect 7 56 8 60
rect 23 64 27 68
rect 23 57 27 60
rect 2 53 8 56
rect 2 49 3 53
rect 7 49 8 53
rect 13 55 17 56
rect 23 52 27 53
rect 33 55 37 56
rect 13 48 17 51
rect 2 44 13 46
rect 33 48 37 51
rect 17 44 23 46
rect 2 42 23 44
rect 2 30 6 42
rect 33 38 37 44
rect 15 34 16 38
rect 20 34 37 38
rect 17 30 30 31
rect 2 29 7 30
rect 2 25 3 29
rect 17 26 26 30
rect 2 22 7 25
rect 2 18 3 22
rect 2 17 7 18
rect 15 18 16 22
rect 20 18 21 22
rect 15 15 21 18
rect 26 17 30 26
rect 33 21 37 34
rect 33 16 37 17
rect 15 12 16 15
rect -2 11 16 12
rect 20 12 21 15
rect 20 11 42 12
rect -2 2 42 11
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
<< ntransistor >>
rect 9 10 11 30
rect 29 10 31 22
<< ptransistor >>
rect 9 43 11 61
rect 19 43 21 65
rect 29 43 31 65
<< polycontact >>
rect 16 34 20 38
rect 26 26 30 30
<< ndcontact >>
rect 3 25 7 29
rect 3 18 7 22
rect 16 18 20 22
rect 16 11 20 15
rect 33 17 37 21
<< pdcontact >>
rect 3 56 7 60
rect 3 49 7 53
rect 13 51 17 55
rect 13 44 17 48
rect 23 60 27 64
rect 23 53 27 57
rect 33 51 37 55
rect 33 44 37 48
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
<< psubstratepdiff >>
rect 0 2 40 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 40 2
rect 0 -3 40 -2
<< nsubstratendiff >>
rect 0 82 40 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 40 82
rect 0 77 40 78
<< labels >>
rlabel ndcontact 4 28 4 28 6 z
rlabel metal1 12 44 12 44 6 z
rlabel metal1 20 6 20 6 6 vss
rlabel metal1 20 28 20 28 6 a
rlabel metal1 28 24 28 24 6 a
rlabel metal1 20 44 20 44 6 z
rlabel metal1 20 74 20 74 6 vdd
rlabel metal1 26 36 26 36 6 an
rlabel metal1 35 36 35 36 6 an
<< end >>
