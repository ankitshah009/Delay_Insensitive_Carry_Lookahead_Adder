magic
tech scmos
timestamp 1179387485
<< checkpaint >>
rect -22 -22 86 94
<< ab >>
rect 0 0 64 72
<< pwell >>
rect -4 -4 68 32
<< nwell >>
rect -4 32 68 76
<< polysilicon >>
rect 11 67 34 69
rect 11 61 13 67
rect 9 58 13 61
rect 22 59 24 63
rect 32 59 34 67
rect 42 65 44 70
rect 49 65 51 70
rect 9 55 11 58
rect 22 44 24 47
rect 9 40 11 43
rect 22 42 27 44
rect 32 42 34 47
rect 42 42 44 47
rect 49 44 51 47
rect 9 39 15 40
rect 9 35 10 39
rect 14 35 15 39
rect 9 34 15 35
rect 13 31 15 34
rect 25 35 27 42
rect 39 40 44 42
rect 48 43 54 44
rect 25 34 31 35
rect 13 29 19 31
rect 25 30 26 34
rect 30 30 31 34
rect 25 29 31 30
rect 17 26 19 29
rect 29 26 31 29
rect 39 26 41 40
rect 48 39 49 43
rect 53 39 54 43
rect 48 38 54 39
rect 49 26 51 38
rect 7 17 13 18
rect 7 13 8 17
rect 12 13 13 17
rect 17 15 19 20
rect 7 12 13 13
rect 29 15 31 20
rect 11 10 13 12
rect 39 10 41 20
rect 49 15 51 20
rect 55 17 61 18
rect 55 13 56 17
rect 60 13 61 17
rect 55 12 61 13
rect 55 10 57 12
rect 11 8 57 10
<< ndiffusion >>
rect 9 25 17 26
rect 9 21 10 25
rect 14 21 17 25
rect 9 20 17 21
rect 19 20 29 26
rect 31 25 39 26
rect 31 21 33 25
rect 37 21 39 25
rect 31 20 39 21
rect 41 25 49 26
rect 41 21 43 25
rect 47 21 49 25
rect 41 20 49 21
rect 51 25 58 26
rect 51 21 53 25
rect 57 21 58 25
rect 51 20 58 21
rect 21 17 27 20
rect 21 13 22 17
rect 26 13 27 17
rect 21 12 27 13
<< pdiffusion >>
rect 53 68 60 69
rect 53 65 54 68
rect 37 59 42 65
rect 15 58 22 59
rect 15 55 16 58
rect 4 49 9 55
rect 2 48 9 49
rect 2 44 3 48
rect 7 44 9 48
rect 2 43 9 44
rect 11 54 16 55
rect 20 54 22 58
rect 11 47 22 54
rect 24 52 32 59
rect 24 48 26 52
rect 30 48 32 52
rect 24 47 32 48
rect 34 58 42 59
rect 34 54 36 58
rect 40 54 42 58
rect 34 47 42 54
rect 44 47 49 65
rect 51 64 54 65
rect 58 64 60 68
rect 51 47 60 64
rect 11 43 20 47
<< metal1 >>
rect -2 68 66 72
rect -2 64 4 68
rect 8 64 54 68
rect 58 64 66 68
rect 15 58 21 64
rect 15 54 16 58
rect 20 54 21 58
rect 35 54 36 58
rect 40 54 62 58
rect 26 52 30 53
rect 2 48 7 49
rect 2 44 3 48
rect 2 43 7 44
rect 17 43 23 50
rect 30 48 38 50
rect 26 46 38 48
rect 2 26 6 43
rect 10 39 23 43
rect 14 38 23 39
rect 34 43 38 46
rect 34 39 49 43
rect 53 39 54 43
rect 10 34 14 35
rect 18 30 26 34
rect 30 30 31 34
rect 2 25 14 26
rect 2 22 10 25
rect 7 21 10 22
rect 18 21 22 30
rect 34 26 38 39
rect 58 34 62 54
rect 33 25 38 26
rect 37 21 38 25
rect 7 20 14 21
rect 33 20 38 21
rect 42 30 62 34
rect 42 25 47 30
rect 42 21 43 25
rect 42 20 47 21
rect 53 25 57 26
rect 7 17 13 20
rect 53 17 57 21
rect 7 13 8 17
rect 12 13 13 17
rect 21 13 22 17
rect 26 13 27 17
rect 53 13 56 17
rect 60 13 61 17
rect 21 8 27 13
rect -2 4 4 8
rect 8 4 66 8
rect -2 0 66 4
<< ntransistor >>
rect 17 20 19 26
rect 29 20 31 26
rect 39 20 41 26
rect 49 20 51 26
<< ptransistor >>
rect 9 43 11 55
rect 22 47 24 59
rect 32 47 34 59
rect 42 47 44 65
rect 49 47 51 65
<< polycontact >>
rect 10 35 14 39
rect 26 30 30 34
rect 49 39 53 43
rect 8 13 12 17
rect 56 13 60 17
<< ndcontact >>
rect 10 21 14 25
rect 33 21 37 25
rect 43 21 47 25
rect 53 21 57 25
rect 22 13 26 17
<< pdcontact >>
rect 3 44 7 48
rect 16 54 20 58
rect 26 48 30 52
rect 36 54 40 58
rect 54 64 58 68
<< psubstratepcontact >>
rect 4 4 8 8
<< nsubstratencontact >>
rect 4 64 8 68
<< psubstratepdiff >>
rect 3 8 9 9
rect 3 4 4 8
rect 8 4 9 8
rect 3 3 9 4
<< nsubstratendiff >>
rect 3 68 9 69
rect 3 64 4 68
rect 8 64 9 68
rect 3 63 9 64
<< labels >>
rlabel polycontact 10 15 10 15 6 bn
rlabel polycontact 58 15 58 15 6 bn
rlabel polycontact 50 42 50 42 6 an
rlabel metal1 10 19 10 19 6 bn
rlabel metal1 12 40 12 40 6 b
rlabel pdcontact 4 46 4 46 6 bn
rlabel polycontact 28 32 28 32 6 a
rlabel metal1 20 24 20 24 6 a
rlabel metal1 20 44 20 44 6 b
rlabel metal1 32 4 32 4 6 vss
rlabel ndcontact 44 24 44 24 6 z
rlabel metal1 36 35 36 35 6 an
rlabel metal1 32 48 32 48 6 an
rlabel metal1 44 56 44 56 6 z
rlabel metal1 32 68 32 68 6 vdd
rlabel metal1 55 19 55 19 6 bn
rlabel metal1 52 32 52 32 6 z
rlabel metal1 44 41 44 41 6 an
rlabel metal1 60 44 60 44 6 z
rlabel metal1 52 56 52 56 6 z
<< end >>
