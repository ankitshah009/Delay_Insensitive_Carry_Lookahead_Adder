magic
tech scmos
timestamp 1179387027
<< checkpaint >>
rect -22 -25 86 105
<< ab >>
rect 0 0 64 80
<< pwell >>
rect -4 -7 68 36
<< nwell >>
rect -4 36 68 87
<< polysilicon >>
rect 10 70 12 74
rect 22 70 24 74
rect 29 70 31 74
rect 39 70 41 74
rect 46 70 48 74
rect 10 39 12 42
rect 22 39 24 42
rect 29 39 31 42
rect 39 39 41 42
rect 9 38 15 39
rect 9 34 10 38
rect 14 34 15 38
rect 9 33 15 34
rect 19 38 25 39
rect 19 34 20 38
rect 24 34 25 38
rect 19 33 25 34
rect 29 38 41 39
rect 29 34 34 38
rect 38 34 41 38
rect 29 33 41 34
rect 46 39 48 42
rect 46 38 55 39
rect 46 34 50 38
rect 54 34 55 38
rect 46 33 55 34
rect 9 30 11 33
rect 30 30 32 33
rect 46 30 48 33
rect 20 24 22 29
rect 9 9 11 12
rect 20 9 22 12
rect 9 7 22 9
rect 30 6 32 10
rect 46 6 48 10
<< ndiffusion >>
rect 4 23 9 30
rect 2 22 9 23
rect 2 18 3 22
rect 7 18 9 22
rect 2 17 9 18
rect 4 12 9 17
rect 11 29 18 30
rect 11 25 13 29
rect 17 25 18 29
rect 11 24 18 25
rect 25 24 30 30
rect 11 12 20 24
rect 22 22 30 24
rect 22 18 24 22
rect 28 18 30 22
rect 22 12 30 18
rect 25 10 30 12
rect 32 15 46 30
rect 32 11 37 15
rect 41 11 46 15
rect 32 10 46 11
rect 48 23 53 30
rect 48 22 55 23
rect 48 18 50 22
rect 54 18 55 22
rect 48 17 55 18
rect 48 10 53 17
<< pdiffusion >>
rect 5 63 10 70
rect 2 62 10 63
rect 2 58 3 62
rect 7 58 10 62
rect 2 55 10 58
rect 2 51 3 55
rect 7 51 10 55
rect 2 50 10 51
rect 5 42 10 50
rect 12 69 22 70
rect 12 65 15 69
rect 19 65 22 69
rect 12 42 22 65
rect 24 42 29 70
rect 31 62 39 70
rect 31 58 33 62
rect 37 58 39 62
rect 31 55 39 58
rect 31 51 33 55
rect 37 51 39 55
rect 31 42 39 51
rect 41 42 46 70
rect 48 69 57 70
rect 48 65 51 69
rect 55 65 57 69
rect 48 62 57 65
rect 48 58 51 62
rect 55 58 57 62
rect 48 42 57 58
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect -2 69 66 78
rect -2 68 15 69
rect 14 65 15 68
rect 19 68 51 69
rect 19 65 20 68
rect 50 65 51 68
rect 55 68 66 69
rect 55 65 56 68
rect 50 62 56 65
rect 2 58 3 62
rect 7 58 33 62
rect 37 58 38 62
rect 50 58 51 62
rect 55 58 56 62
rect 2 55 7 58
rect 2 51 3 55
rect 33 55 38 58
rect 2 50 7 51
rect 2 29 6 50
rect 17 47 23 54
rect 37 51 38 55
rect 33 50 38 51
rect 10 42 23 47
rect 42 46 46 55
rect 10 38 14 42
rect 33 41 46 46
rect 33 38 39 41
rect 19 34 20 38
rect 24 34 27 38
rect 33 34 34 38
rect 38 34 39 38
rect 50 38 55 47
rect 54 34 55 38
rect 10 33 14 34
rect 23 30 27 34
rect 50 30 55 34
rect 2 25 13 29
rect 17 25 18 29
rect 23 26 55 30
rect 2 18 3 22
rect 7 18 24 22
rect 28 18 50 22
rect 54 18 55 22
rect 36 12 37 15
rect -2 11 37 12
rect 41 12 42 15
rect 41 11 66 12
rect -2 2 66 11
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
<< ntransistor >>
rect 9 12 11 30
rect 20 12 22 24
rect 30 10 32 30
rect 46 10 48 30
<< ptransistor >>
rect 10 42 12 70
rect 22 42 24 70
rect 29 42 31 70
rect 39 42 41 70
rect 46 42 48 70
<< polycontact >>
rect 10 34 14 38
rect 20 34 24 38
rect 34 34 38 38
rect 50 34 54 38
<< ndcontact >>
rect 3 18 7 22
rect 13 25 17 29
rect 24 18 28 22
rect 37 11 41 15
rect 50 18 54 22
<< pdcontact >>
rect 3 58 7 62
rect 3 51 7 55
rect 15 65 19 69
rect 33 58 37 62
rect 33 51 37 55
rect 51 65 55 69
rect 51 58 55 62
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
<< psubstratepdiff >>
rect 0 2 64 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 64 2
rect 0 -3 64 -2
<< nsubstratendiff >>
rect 0 82 64 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 64 82
rect 0 77 64 78
<< labels >>
rlabel metal1 4 40 4 40 6 z
rlabel metal1 12 40 12 40 6 b
rlabel metal1 20 48 20 48 6 b
rlabel metal1 12 60 12 60 6 z
rlabel metal1 20 60 20 60 6 z
rlabel metal1 32 6 32 6 6 vss
rlabel metal1 28 28 28 28 6 a1
rlabel metal1 36 28 36 28 6 a1
rlabel metal1 36 40 36 40 6 a2
rlabel metal1 28 60 28 60 6 z
rlabel metal1 32 74 32 74 6 vdd
rlabel metal1 44 28 44 28 6 a1
rlabel metal1 44 48 44 48 6 a2
rlabel metal1 28 20 28 20 6 n1
rlabel polycontact 52 36 52 36 6 a1
<< end >>
