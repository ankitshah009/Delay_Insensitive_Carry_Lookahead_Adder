magic
tech scmos
timestamp 1179386357
<< checkpaint >>
rect -22 -25 70 105
<< ab >>
rect 0 0 48 80
<< pwell >>
rect -4 -7 52 36
<< nwell >>
rect -4 36 52 87
<< polysilicon >>
rect 9 67 11 72
rect 19 67 21 72
rect 9 30 11 50
rect 19 47 21 50
rect 19 46 31 47
rect 19 45 26 46
rect 25 42 26 45
rect 30 42 31 46
rect 25 41 31 42
rect 26 35 28 41
rect 35 38 41 39
rect 35 36 36 38
rect 16 33 28 35
rect 16 30 18 33
rect 26 30 28 33
rect 33 34 36 36
rect 40 34 41 38
rect 33 33 41 34
rect 33 30 35 33
rect 9 8 11 16
rect 16 12 18 16
rect 26 12 28 16
rect 33 8 35 16
rect 9 6 35 8
<< ndiffusion >>
rect 2 28 9 30
rect 2 24 3 28
rect 7 24 9 28
rect 2 21 9 24
rect 2 17 3 21
rect 7 17 9 21
rect 2 16 9 17
rect 11 16 16 30
rect 18 29 26 30
rect 18 25 20 29
rect 24 25 26 29
rect 18 22 26 25
rect 18 18 20 22
rect 24 18 26 22
rect 18 16 26 18
rect 28 16 33 30
rect 35 28 43 30
rect 35 24 37 28
rect 41 24 43 28
rect 35 21 43 24
rect 35 17 37 21
rect 41 17 43 21
rect 35 16 43 17
<< pdiffusion >>
rect 2 66 9 67
rect 2 62 3 66
rect 7 62 9 66
rect 2 59 9 62
rect 2 55 3 59
rect 7 55 9 59
rect 2 50 9 55
rect 11 55 19 67
rect 11 51 13 55
rect 17 51 19 55
rect 11 50 19 51
rect 21 66 29 67
rect 21 62 23 66
rect 27 62 29 66
rect 21 50 29 62
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect -2 68 50 78
rect 3 66 7 68
rect 3 59 7 62
rect 23 66 27 68
rect 23 61 27 62
rect 3 54 7 55
rect 10 51 13 55
rect 17 51 18 55
rect 10 31 14 51
rect 26 49 38 55
rect 26 46 30 49
rect 26 41 30 42
rect 42 39 46 47
rect 34 38 46 39
rect 34 34 36 38
rect 40 34 46 38
rect 34 33 46 34
rect 10 29 24 31
rect 3 28 7 29
rect 10 27 20 29
rect 3 21 7 24
rect 18 25 20 27
rect 18 22 24 25
rect 18 18 20 22
rect 18 17 24 18
rect 36 24 37 28
rect 41 24 42 28
rect 36 21 42 24
rect 36 17 37 21
rect 41 17 42 21
rect 3 12 7 17
rect 36 12 42 17
rect -2 2 50 12
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
<< ntransistor >>
rect 9 16 11 30
rect 16 16 18 30
rect 26 16 28 30
rect 33 16 35 30
<< ptransistor >>
rect 9 50 11 67
rect 19 50 21 67
<< polycontact >>
rect 26 42 30 46
rect 36 34 40 38
<< ndcontact >>
rect 3 24 7 28
rect 3 17 7 21
rect 20 25 24 29
rect 20 18 24 22
rect 37 24 41 28
rect 37 17 41 21
<< pdcontact >>
rect 3 62 7 66
rect 3 55 7 59
rect 13 51 17 55
rect 23 62 27 66
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
<< psubstratepdiff >>
rect 0 2 48 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 48 2
rect 0 -3 48 -2
<< nsubstratendiff >>
rect 0 82 48 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 48 82
rect 0 77 48 78
<< labels >>
rlabel metal1 20 24 20 24 6 z
rlabel metal1 12 44 12 44 6 z
rlabel metal1 24 6 24 6 6 vss
rlabel metal1 28 48 28 48 6 b
rlabel metal1 24 74 24 74 6 vdd
rlabel metal1 36 36 36 36 6 a
rlabel metal1 44 40 44 40 6 a
rlabel metal1 36 52 36 52 6 b
<< end >>
