magic
tech scmos
timestamp 1182409147
<< checkpaint >>
rect -22 -22 118 94
<< ab >>
rect 0 0 96 72
<< pwell >>
rect -4 -4 100 32
<< nwell >>
rect -4 32 100 76
<< polysilicon >>
rect 9 66 11 70
rect 19 66 21 70
rect 29 66 31 70
rect 39 66 41 70
rect 49 66 51 70
rect 59 66 61 70
rect 69 66 71 70
rect 79 66 81 70
rect 9 35 11 38
rect 19 35 21 38
rect 29 35 31 38
rect 39 35 41 38
rect 9 34 15 35
rect 9 30 10 34
rect 14 30 15 34
rect 9 29 15 30
rect 19 34 31 35
rect 19 30 26 34
rect 30 30 31 34
rect 19 29 31 30
rect 35 34 41 35
rect 35 30 36 34
rect 40 31 41 34
rect 49 31 51 38
rect 59 35 61 38
rect 69 35 71 38
rect 79 35 81 38
rect 58 34 71 35
rect 40 30 53 31
rect 35 29 53 30
rect 12 26 14 29
rect 19 26 21 29
rect 29 26 31 29
rect 36 26 38 29
rect 51 26 53 29
rect 58 30 60 34
rect 64 30 71 34
rect 58 29 71 30
rect 75 34 81 35
rect 75 30 76 34
rect 80 30 81 34
rect 75 29 81 30
rect 58 26 60 29
rect 68 26 70 29
rect 75 26 77 29
rect 68 8 70 13
rect 75 8 77 13
rect 12 2 14 6
rect 19 2 21 6
rect 29 2 31 6
rect 36 2 38 6
rect 51 2 53 7
rect 58 2 60 7
<< ndiffusion >>
rect 3 11 12 26
rect 3 7 5 11
rect 9 7 12 11
rect 3 6 12 7
rect 14 6 19 26
rect 21 18 29 26
rect 21 14 23 18
rect 27 14 29 18
rect 21 6 29 14
rect 31 6 36 26
rect 38 11 51 26
rect 38 7 43 11
rect 47 7 51 11
rect 53 7 58 26
rect 60 18 68 26
rect 60 14 62 18
rect 66 14 68 18
rect 60 13 68 14
rect 70 13 75 26
rect 77 25 86 26
rect 77 21 80 25
rect 84 21 86 25
rect 77 18 86 21
rect 77 14 80 18
rect 84 14 86 18
rect 77 13 86 14
rect 60 7 65 13
rect 38 6 49 7
<< pdiffusion >>
rect 2 65 9 66
rect 2 61 3 65
rect 7 61 9 65
rect 2 58 9 61
rect 2 54 3 58
rect 7 54 9 58
rect 2 38 9 54
rect 11 57 19 66
rect 11 53 13 57
rect 17 53 19 57
rect 11 50 19 53
rect 11 46 13 50
rect 17 46 19 50
rect 11 38 19 46
rect 21 65 29 66
rect 21 61 23 65
rect 27 61 29 65
rect 21 58 29 61
rect 21 54 23 58
rect 27 54 29 58
rect 21 38 29 54
rect 31 58 39 66
rect 31 54 33 58
rect 37 54 39 58
rect 31 50 39 54
rect 31 46 33 50
rect 37 46 39 50
rect 31 38 39 46
rect 41 65 49 66
rect 41 61 43 65
rect 47 61 49 65
rect 41 58 49 61
rect 41 54 43 58
rect 47 54 49 58
rect 41 38 49 54
rect 51 50 59 66
rect 51 46 53 50
rect 57 46 59 50
rect 51 43 59 46
rect 51 39 53 43
rect 57 39 59 43
rect 51 38 59 39
rect 61 65 69 66
rect 61 61 63 65
rect 67 61 69 65
rect 61 58 69 61
rect 61 54 63 58
rect 67 54 69 58
rect 61 38 69 54
rect 71 50 79 66
rect 71 46 73 50
rect 77 46 79 50
rect 71 43 79 46
rect 71 39 73 43
rect 77 39 79 43
rect 71 38 79 39
rect 81 65 89 66
rect 81 61 83 65
rect 87 61 89 65
rect 81 58 89 61
rect 81 54 83 58
rect 87 54 89 58
rect 81 38 89 54
<< metal1 >>
rect -2 65 98 72
rect -2 64 3 65
rect 2 61 3 64
rect 7 64 23 65
rect 7 61 8 64
rect 2 58 8 61
rect 22 61 23 64
rect 27 64 43 65
rect 27 61 28 64
rect 22 58 28 61
rect 42 61 43 64
rect 47 64 63 65
rect 47 61 48 64
rect 2 54 3 58
rect 7 54 8 58
rect 13 57 17 58
rect 22 54 23 58
rect 27 54 28 58
rect 33 58 38 59
rect 37 54 38 58
rect 42 58 48 61
rect 42 54 43 58
rect 47 54 48 58
rect 62 61 63 64
rect 67 64 83 65
rect 67 61 68 64
rect 62 58 68 61
rect 62 54 63 58
rect 67 54 68 58
rect 82 61 83 64
rect 87 64 98 65
rect 87 61 88 64
rect 82 58 88 61
rect 82 54 83 58
rect 87 54 88 58
rect 13 50 17 53
rect 33 50 38 54
rect 73 50 79 51
rect 2 46 13 50
rect 17 46 33 50
rect 37 46 53 50
rect 57 46 58 50
rect 2 18 6 46
rect 53 43 58 46
rect 25 38 49 42
rect 57 42 58 43
rect 77 46 79 50
rect 73 43 79 46
rect 57 39 73 42
rect 77 39 79 43
rect 53 38 79 39
rect 10 34 14 35
rect 25 34 31 38
rect 45 34 49 38
rect 25 30 26 34
rect 30 30 31 34
rect 35 30 36 34
rect 40 30 41 34
rect 45 30 60 34
rect 64 30 65 34
rect 71 30 76 34
rect 80 30 87 34
rect 10 26 14 30
rect 35 26 41 30
rect 71 26 75 30
rect 10 22 75 26
rect 79 21 80 25
rect 84 21 85 25
rect 79 18 85 21
rect 2 14 23 18
rect 27 14 62 18
rect 66 14 67 18
rect 79 14 80 18
rect 84 14 85 18
rect 4 8 5 11
rect -2 7 5 8
rect 9 8 10 11
rect 42 8 43 11
rect 9 7 43 8
rect 47 8 48 11
rect 79 8 85 14
rect 47 7 84 8
rect -2 4 84 7
rect 88 4 98 8
rect -2 0 98 4
<< ntransistor >>
rect 12 6 14 26
rect 19 6 21 26
rect 29 6 31 26
rect 36 6 38 26
rect 51 7 53 26
rect 58 7 60 26
rect 68 13 70 26
rect 75 13 77 26
<< ptransistor >>
rect 9 38 11 66
rect 19 38 21 66
rect 29 38 31 66
rect 39 38 41 66
rect 49 38 51 66
rect 59 38 61 66
rect 69 38 71 66
rect 79 38 81 66
<< polycontact >>
rect 10 30 14 34
rect 26 30 30 34
rect 36 30 40 34
rect 60 30 64 34
rect 76 30 80 34
<< ndcontact >>
rect 5 7 9 11
rect 23 14 27 18
rect 43 7 47 11
rect 62 14 66 18
rect 80 21 84 25
rect 80 14 84 18
<< pdcontact >>
rect 3 61 7 65
rect 3 54 7 58
rect 13 53 17 57
rect 13 46 17 50
rect 23 61 27 65
rect 23 54 27 58
rect 33 54 37 58
rect 33 46 37 50
rect 43 61 47 65
rect 43 54 47 58
rect 53 46 57 50
rect 53 39 57 43
rect 63 61 67 65
rect 63 54 67 58
rect 73 46 77 50
rect 73 39 77 43
rect 83 61 87 65
rect 83 54 87 58
<< psubstratepcontact >>
rect 84 4 88 8
<< psubstratepdiff >>
rect 83 8 89 9
rect 83 4 84 8
rect 88 4 89 8
rect 83 3 89 4
<< labels >>
rlabel metal1 12 16 12 16 6 z
rlabel metal1 4 32 4 32 6 z
rlabel polycontact 12 32 12 32 6 a
rlabel metal1 12 48 12 48 6 z
rlabel metal1 28 16 28 16 6 z
rlabel metal1 20 16 20 16 6 z
rlabel metal1 20 24 20 24 6 a
rlabel metal1 28 24 28 24 6 a
rlabel metal1 28 36 28 36 6 b
rlabel metal1 20 48 20 48 6 z
rlabel metal1 28 48 28 48 6 z
rlabel metal1 48 4 48 4 6 vss
rlabel metal1 52 16 52 16 6 z
rlabel metal1 44 16 44 16 6 z
rlabel metal1 36 16 36 16 6 z
rlabel metal1 36 24 36 24 6 a
rlabel metal1 52 24 52 24 6 a
rlabel metal1 44 24 44 24 6 a
rlabel metal1 52 32 52 32 6 b
rlabel metal1 36 40 36 40 6 b
rlabel metal1 44 40 44 40 6 b
rlabel metal1 36 52 36 52 6 z
rlabel metal1 52 48 52 48 6 z
rlabel metal1 44 48 44 48 6 z
rlabel metal1 48 68 48 68 6 vdd
rlabel metal1 60 16 60 16 6 z
rlabel metal1 60 24 60 24 6 a
rlabel metal1 68 24 68 24 6 a
rlabel metal1 76 32 76 32 6 a
rlabel metal1 60 32 60 32 6 b
rlabel metal1 60 40 60 40 6 z
rlabel metal1 68 40 68 40 6 z
rlabel metal1 76 44 76 44 6 z
rlabel metal1 84 32 84 32 6 a
<< end >>
