magic
tech scmos
timestamp 1179386520
<< checkpaint >>
rect -22 -22 78 94
<< ab >>
rect 0 0 56 72
<< pwell >>
rect -4 -4 60 32
<< nwell >>
rect -4 32 60 76
<< polysilicon >>
rect 9 56 11 61
rect 21 56 23 61
rect 31 56 33 61
rect 45 60 47 65
rect 9 28 11 46
rect 21 35 23 46
rect 31 35 33 46
rect 45 45 47 48
rect 41 44 47 45
rect 41 40 42 44
rect 46 40 47 44
rect 41 39 47 40
rect 19 34 25 35
rect 19 30 20 34
rect 24 30 25 34
rect 19 29 25 30
rect 31 34 41 35
rect 31 30 36 34
rect 40 30 41 34
rect 31 29 41 30
rect 9 27 15 28
rect 9 23 10 27
rect 14 25 15 27
rect 14 23 17 25
rect 9 22 17 23
rect 15 19 17 22
rect 22 19 24 29
rect 31 25 33 29
rect 45 26 47 39
rect 29 22 33 25
rect 29 19 31 22
rect 45 15 47 20
rect 15 4 17 9
rect 22 4 24 9
rect 29 4 31 9
<< ndiffusion >>
rect 35 20 45 26
rect 47 25 54 26
rect 47 21 49 25
rect 53 21 54 25
rect 47 20 54 21
rect 35 19 43 20
rect 8 17 15 19
rect 8 13 9 17
rect 13 13 15 17
rect 8 12 15 13
rect 10 9 15 12
rect 17 9 22 19
rect 24 9 29 19
rect 31 16 43 19
rect 31 12 36 16
rect 40 12 43 16
rect 31 9 43 12
<< pdiffusion >>
rect 35 56 45 60
rect 4 52 9 56
rect 2 51 9 52
rect 2 47 3 51
rect 7 47 9 51
rect 2 46 9 47
rect 11 55 21 56
rect 11 51 14 55
rect 18 51 21 55
rect 11 46 21 51
rect 23 51 31 56
rect 23 47 25 51
rect 29 47 31 51
rect 23 46 31 47
rect 33 55 45 56
rect 33 51 35 55
rect 39 51 45 55
rect 33 48 45 51
rect 47 54 52 60
rect 47 53 54 54
rect 47 49 49 53
rect 53 49 54 53
rect 47 48 54 49
rect 33 46 39 48
<< metal1 >>
rect -2 68 58 72
rect -2 64 4 68
rect 8 64 12 68
rect 16 64 58 68
rect 14 55 18 64
rect 2 51 7 52
rect 2 47 3 51
rect 35 55 39 64
rect 14 50 18 51
rect 25 51 29 52
rect 2 42 7 47
rect 35 50 39 51
rect 25 42 29 47
rect 42 44 46 59
rect 2 38 29 42
rect 33 40 42 42
rect 33 38 46 40
rect 49 53 53 54
rect 2 17 6 38
rect 49 34 53 49
rect 19 30 20 34
rect 24 30 31 34
rect 35 30 36 34
rect 40 30 53 34
rect 10 27 14 28
rect 26 27 31 30
rect 14 23 22 25
rect 10 21 22 23
rect 26 21 38 27
rect 49 25 53 30
rect 2 13 9 17
rect 13 13 14 17
rect 18 13 22 21
rect 49 20 53 21
rect 36 16 40 17
rect 36 8 40 12
rect -2 4 48 8
rect 52 4 58 8
rect -2 0 58 4
<< ntransistor >>
rect 45 20 47 26
rect 15 9 17 19
rect 22 9 24 19
rect 29 9 31 19
<< ptransistor >>
rect 9 46 11 56
rect 21 46 23 56
rect 31 46 33 56
rect 45 48 47 60
<< polycontact >>
rect 42 40 46 44
rect 20 30 24 34
rect 36 30 40 34
rect 10 23 14 27
<< ndcontact >>
rect 49 21 53 25
rect 9 13 13 17
rect 36 12 40 16
<< pdcontact >>
rect 3 47 7 51
rect 14 51 18 55
rect 25 47 29 51
rect 35 51 39 55
rect 49 49 53 53
<< psubstratepcontact >>
rect 48 4 52 8
<< nsubstratencontact >>
rect 4 64 8 68
rect 12 64 16 68
<< psubstratepdiff >>
rect 47 8 53 9
rect 47 4 48 8
rect 52 4 53 8
rect 47 3 53 4
<< nsubstratendiff >>
rect 3 68 17 69
rect 3 64 4 68
rect 8 64 12 68
rect 16 64 17 68
rect 3 63 17 64
<< labels >>
rlabel polysilicon 36 32 36 32 6 an
rlabel metal1 4 32 4 32 6 z
rlabel metal1 20 16 20 16 6 c
rlabel polycontact 12 24 12 24 6 c
rlabel metal1 20 40 20 40 6 z
rlabel metal1 12 40 12 40 6 z
rlabel metal1 28 4 28 4 6 vss
rlabel metal1 28 28 28 28 6 b
rlabel metal1 36 24 36 24 6 b
rlabel metal1 36 40 36 40 6 a
rlabel metal1 28 68 28 68 6 vdd
rlabel metal1 44 32 44 32 6 an
rlabel metal1 51 37 51 37 6 an
rlabel metal1 44 52 44 52 6 a
<< end >>
