.subckt noa2ao222_x1 i0 i1 i2 i3 i4 nq vdd vss
*   SPICE3 file   created from noa2ao222_x1.ext -      technology: scmos
m00 vdd    i0     w1     vdd p w=29u  l=2.3636u ad=172p     pd=48u      as=186.188p ps=56.7391u
m01 w1     i1     vdd    vdd p w=29u  l=2.3636u ad=186.188p pd=56.7391u as=172p     ps=48u
m02 nq     i4     w1     vdd p w=40u  l=2.3636u ad=200p     pd=50u      as=256.812p ps=78.2609u
m03 w2     i2     nq     vdd p w=40u  l=2.3636u ad=160p     pd=48u      as=200p     ps=50u
m04 w1     i3     w2     vdd p w=40u  l=2.3636u ad=256.812p pd=78.2609u as=160p     ps=48u
m05 w3     i0     vss    vss n w=18u  l=2.3636u ad=72p      pd=26u      as=148p     ps=49.3333u
m06 nq     i1     w3     vss n w=18u  l=2.3636u ad=90p      pd=28u      as=72p      ps=26u
m07 w4     i4     nq     vss n w=18u  l=2.3636u ad=108p     pd=36u      as=90p      ps=28u
m08 vss    i2     w4     vss n w=18u  l=2.3636u ad=148p     pd=49.3333u as=108p     ps=36u
m09 w4     i3     vss    vss n w=18u  l=2.3636u ad=108p     pd=36u      as=148p     ps=49.3333u
C0  w1     i4     0.086f
C1  i1     i2     0.060f
C2  w3     i1     0.012f
C3  w4     i0     0.006f
C4  vdd    i2     0.012f
C5  i0     i4     0.097f
C6  nq     w1     0.068f
C7  w4     i3     0.050f
C8  vss    i0     0.063f
C9  i3     i4     0.064f
C10 w1     i1     0.036f
C11 w2     vdd    0.019f
C12 vss    i3     0.016f
C13 nq     i0     0.084f
C14 w4     vss    0.225f
C15 vss    i4     0.009f
C16 w2     i2     0.012f
C17 i1     i0     0.398f
C18 nq     i3     0.097f
C19 w1     vdd    0.463f
C20 w4     nq     0.117f
C21 nq     i4     0.350f
C22 i0     vdd    0.023f
C23 i1     i3     0.051f
C24 w1     i2     0.017f
C25 vss    nq     0.091f
C26 i0     i2     0.042f
C27 vdd    i3     0.017f
C28 i1     i4     0.319f
C29 w2     w1     0.016f
C30 vss    i1     0.013f
C31 w3     i0     0.009f
C32 vdd    i4     0.017f
C33 i3     i2     0.322f
C34 nq     i1     0.126f
C35 w4     i2     0.036f
C36 i2     i4     0.094f
C37 nq     vdd    0.041f
C38 w2     i3     0.009f
C39 vss    i2     0.028f
C40 w1     i0     0.064f
C41 i1     vdd    0.050f
C42 w1     i3     0.064f
C43 nq     i2     0.262f
C45 nq     vss    0.015f
C46 i1     vss    0.024f
C47 i0     vss    0.023f
C49 i3     vss    0.023f
C50 i2     vss    0.024f
C51 i4     vss    0.028f
.ends
