.subckt noa2a22_x1 i0 i1 i2 i3 nq vdd vss
*   SPICE3 file   created from noa2a22_x1.ext -      technology: scmos
m00 nq     i0     w1     vdd p w=39u  l=2.3636u ad=195p     pd=49u      as=244.5p   ps=71.5u
m01 w1     i1     nq     vdd p w=39u  l=2.3636u ad=244.5p   pd=71.5u    as=195p     ps=49u
m02 vdd    i3     w1     vdd p w=39u  l=2.3636u ad=195p     pd=49u      as=244.5p   ps=71.5u
m03 w1     i2     vdd    vdd p w=39u  l=2.3636u ad=244.5p   pd=71.5u    as=195p     ps=49u
m04 w2     i0     vss    vss n w=19u  l=2.3636u ad=95p      pd=29u      as=152p     ps=54u
m05 nq     i1     w2     vss n w=19u  l=2.3636u ad=95p      pd=29u      as=95p      ps=29u
m06 w3     i3     nq     vss n w=19u  l=2.3636u ad=95p      pd=29u      as=95p      ps=29u
m07 vss    i2     w3     vss n w=19u  l=2.3636u ad=152p     pd=54u      as=95p      ps=29u
C0  vdd    i2     0.061f
C1  vss    i3     0.029f
C2  nq     w1     0.150f
C3  w2     i1     0.018f
C4  vss    i0     0.040f
C5  w1     i2     0.053f
C6  nq     i3     0.283f
C7  vdd    i1     0.014f
C8  w3     vss    0.019f
C9  w1     i1     0.013f
C10 i2     i3     0.361f
C11 nq     i0     0.087f
C12 i3     i1     0.150f
C13 i2     i0     0.057f
C14 vss    nq     0.043f
C15 i1     i0     0.310f
C16 vss    i2     0.040f
C17 vdd    w1     0.366f
C18 nq     i2     0.106f
C19 vdd    i3     0.074f
C20 vss    i1     0.029f
C21 vdd    i0     0.010f
C22 w1     i3     0.029f
C23 nq     i1     0.280f
C24 w2     vss    0.019f
C25 i2     i1     0.082f
C26 w1     i0     0.024f
C27 vss    vdd    0.003f
C28 i3     i0     0.082f
C29 vdd    nq     0.068f
C30 w3     i3     0.018f
C33 nq     vss    0.015f
C34 i2     vss    0.030f
C35 i3     vss    0.035f
C36 i1     vss    0.035f
C37 i0     vss    0.030f
.ends
