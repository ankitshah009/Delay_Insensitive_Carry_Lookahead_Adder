magic
tech scmos
timestamp 1179385849
<< checkpaint >>
rect -22 -25 62 105
<< ab >>
rect 0 0 40 80
<< pwell >>
rect -4 -7 44 36
<< nwell >>
rect -4 36 44 87
<< polysilicon >>
rect 9 69 11 74
rect 19 69 21 74
rect 29 69 31 74
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 9 38 31 39
rect 9 34 18 38
rect 22 34 26 38
rect 30 34 31 38
rect 9 33 31 34
rect 9 30 11 33
rect 19 30 21 33
rect 9 6 11 10
rect 19 6 21 10
<< ndiffusion >>
rect 2 22 9 30
rect 2 18 3 22
rect 7 18 9 22
rect 2 15 9 18
rect 2 11 3 15
rect 7 11 9 15
rect 2 10 9 11
rect 11 29 19 30
rect 11 25 13 29
rect 17 25 19 29
rect 11 22 19 25
rect 11 18 13 22
rect 17 18 19 22
rect 11 10 19 18
rect 21 29 29 30
rect 21 25 23 29
rect 27 25 29 29
rect 21 22 29 25
rect 21 18 23 22
rect 27 18 29 22
rect 21 17 29 18
rect 21 10 27 17
<< pdiffusion >>
rect 4 55 9 69
rect 2 54 9 55
rect 2 50 3 54
rect 7 50 9 54
rect 2 47 9 50
rect 2 43 3 47
rect 7 43 9 47
rect 2 42 9 43
rect 11 68 19 69
rect 11 64 13 68
rect 17 64 19 68
rect 11 60 19 64
rect 11 56 13 60
rect 17 56 19 60
rect 11 42 19 56
rect 21 54 29 69
rect 21 50 23 54
rect 27 50 29 54
rect 21 47 29 50
rect 21 43 23 47
rect 27 43 29 47
rect 21 42 29 43
rect 31 68 38 69
rect 31 64 33 68
rect 37 64 38 68
rect 31 60 38 64
rect 31 56 33 60
rect 37 56 38 60
rect 31 42 38 56
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect -2 68 42 78
rect 13 60 17 64
rect 13 55 17 56
rect 33 60 37 64
rect 33 55 37 56
rect 2 54 7 55
rect 2 50 3 54
rect 2 47 7 50
rect 2 43 3 47
rect 23 54 27 55
rect 23 47 27 50
rect 7 43 23 46
rect 2 42 27 43
rect 2 30 6 42
rect 34 38 38 47
rect 17 34 18 38
rect 22 34 26 38
rect 30 34 38 38
rect 2 29 17 30
rect 2 26 13 29
rect 13 22 17 25
rect 2 18 3 22
rect 7 18 8 22
rect 2 15 8 18
rect 13 17 17 18
rect 22 25 23 29
rect 27 25 28 29
rect 34 25 38 34
rect 22 22 28 25
rect 22 18 23 22
rect 27 18 28 22
rect 2 12 3 15
rect -2 11 3 12
rect 7 12 8 15
rect 22 12 28 18
rect 7 11 42 12
rect -2 2 42 11
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
<< ntransistor >>
rect 9 10 11 30
rect 19 10 21 30
<< ptransistor >>
rect 9 42 11 69
rect 19 42 21 69
rect 29 42 31 69
<< polycontact >>
rect 18 34 22 38
rect 26 34 30 38
<< ndcontact >>
rect 3 18 7 22
rect 3 11 7 15
rect 13 25 17 29
rect 13 18 17 22
rect 23 25 27 29
rect 23 18 27 22
<< pdcontact >>
rect 3 50 7 54
rect 3 43 7 47
rect 13 64 17 68
rect 13 56 17 60
rect 23 50 27 54
rect 23 43 27 47
rect 33 64 37 68
rect 33 56 37 60
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
<< psubstratepdiff >>
rect 0 2 40 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 40 2
rect 0 -3 40 -2
<< nsubstratendiff >>
rect 0 82 40 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 40 82
rect 0 77 40 78
<< labels >>
rlabel pdcontact 4 44 4 44 6 z
rlabel metal1 12 28 12 28 6 z
rlabel metal1 12 44 12 44 6 z
rlabel metal1 20 6 20 6 6 vss
rlabel polycontact 20 36 20 36 6 a
rlabel metal1 20 44 20 44 6 z
rlabel metal1 20 74 20 74 6 vdd
rlabel metal1 36 36 36 36 6 a
<< end >>
