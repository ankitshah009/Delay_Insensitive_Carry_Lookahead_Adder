magic
tech scmos
timestamp 1180640122
<< checkpaint >>
rect -24 -26 84 126
<< ab >>
rect 0 0 60 100
<< pwell >>
rect -4 -6 64 49
<< nwell >>
rect -4 49 64 106
<< polysilicon >>
rect 17 94 19 98
rect 25 94 27 98
rect 37 94 39 98
rect 45 94 47 98
rect 17 52 19 55
rect 25 52 27 55
rect 15 51 21 52
rect 15 48 16 51
rect 11 47 16 48
rect 20 47 21 51
rect 11 46 21 47
rect 25 51 33 52
rect 25 47 28 51
rect 32 47 33 51
rect 25 46 33 47
rect 11 34 13 46
rect 25 40 27 46
rect 37 43 39 55
rect 45 52 47 55
rect 45 51 53 52
rect 45 49 48 51
rect 47 47 48 49
rect 52 47 53 51
rect 47 46 53 47
rect 37 42 43 43
rect 37 40 38 42
rect 23 37 27 40
rect 35 38 38 40
rect 42 38 43 42
rect 35 37 43 38
rect 23 34 25 37
rect 35 34 37 37
rect 47 34 49 46
rect 11 12 13 17
rect 23 12 25 17
rect 35 12 37 17
rect 47 12 49 17
<< ndiffusion >>
rect 6 23 11 34
rect 3 22 11 23
rect 3 18 4 22
rect 8 18 11 22
rect 3 17 11 18
rect 13 32 23 34
rect 13 28 16 32
rect 20 28 23 32
rect 13 17 23 28
rect 25 22 35 34
rect 25 18 28 22
rect 32 18 35 22
rect 25 17 35 18
rect 37 17 47 34
rect 49 31 54 34
rect 49 30 57 31
rect 49 26 52 30
rect 56 26 57 30
rect 49 22 57 26
rect 49 18 52 22
rect 56 18 57 22
rect 49 17 57 18
rect 39 12 45 17
rect 39 8 40 12
rect 44 8 45 12
rect 39 7 45 8
<< pdiffusion >>
rect 8 92 17 94
rect 8 88 10 92
rect 14 88 17 92
rect 8 82 17 88
rect 8 78 10 82
rect 14 78 17 82
rect 8 55 17 78
rect 19 55 25 94
rect 27 82 37 94
rect 27 78 30 82
rect 34 78 37 82
rect 27 72 37 78
rect 27 68 30 72
rect 34 68 37 72
rect 27 55 37 68
rect 39 55 45 94
rect 47 92 56 94
rect 47 88 50 92
rect 54 88 56 92
rect 47 82 56 88
rect 47 78 50 82
rect 54 78 56 82
rect 47 55 56 78
<< metal1 >>
rect -2 92 62 100
rect -2 88 10 92
rect 14 88 50 92
rect 54 88 62 92
rect 10 82 14 88
rect 10 77 14 78
rect 28 82 34 83
rect 28 78 30 82
rect 28 73 34 78
rect 50 82 54 88
rect 50 77 54 78
rect 8 72 34 73
rect 8 68 30 72
rect 8 67 34 68
rect 38 67 52 73
rect 8 32 12 67
rect 18 58 33 63
rect 18 52 22 58
rect 16 51 22 52
rect 20 47 22 51
rect 16 46 22 47
rect 18 37 22 46
rect 28 51 32 53
rect 28 32 32 47
rect 37 42 42 63
rect 48 51 52 67
rect 48 46 52 47
rect 37 38 38 42
rect 42 38 53 42
rect 8 28 16 32
rect 20 28 23 32
rect 8 27 23 28
rect 28 27 43 32
rect 51 26 52 30
rect 56 26 57 30
rect 51 22 57 26
rect 3 18 4 22
rect 8 18 28 22
rect 32 18 52 22
rect 56 18 57 22
rect -2 8 40 12
rect 44 8 62 12
rect -2 0 62 8
<< ntransistor >>
rect 11 17 13 34
rect 23 17 25 34
rect 35 17 37 34
rect 47 17 49 34
<< ptransistor >>
rect 17 55 19 94
rect 25 55 27 94
rect 37 55 39 94
rect 45 55 47 94
<< polycontact >>
rect 16 47 20 51
rect 28 47 32 51
rect 48 47 52 51
rect 38 38 42 42
<< ndcontact >>
rect 4 18 8 22
rect 16 28 20 32
rect 28 18 32 22
rect 52 26 56 30
rect 52 18 56 22
rect 40 8 44 12
<< pdcontact >>
rect 10 88 14 92
rect 10 78 14 82
rect 30 78 34 82
rect 30 68 34 72
rect 50 88 54 92
rect 50 78 54 82
<< psubstratepcontact >>
rect 8 4 12 8
rect 18 4 22 8
<< psubstratepdiff >>
rect 7 8 23 9
rect 7 4 8 8
rect 12 4 18 8
rect 22 4 23 8
rect 7 3 23 4
<< labels >>
rlabel metal1 20 30 20 30 6 z
rlabel metal1 20 30 20 30 6 z
rlabel metal1 10 50 10 50 6 z
rlabel metal1 10 50 10 50 6 z
rlabel metal1 20 50 20 50 6 b1
rlabel metal1 20 50 20 50 6 b1
rlabel metal1 20 70 20 70 6 z
rlabel metal1 20 70 20 70 6 z
rlabel metal1 30 6 30 6 6 vss
rlabel metal1 30 6 30 6 6 vss
rlabel metal1 30 40 30 40 6 b2
rlabel metal1 30 40 30 40 6 b2
rlabel metal1 30 60 30 60 6 b1
rlabel metal1 30 60 30 60 6 b1
rlabel metal1 30 75 30 75 6 z
rlabel metal1 30 75 30 75 6 z
rlabel metal1 30 94 30 94 6 vdd
rlabel metal1 30 94 30 94 6 vdd
rlabel metal1 40 30 40 30 6 b2
rlabel metal1 40 30 40 30 6 b2
rlabel metal1 40 50 40 50 6 a2
rlabel metal1 40 50 40 50 6 a2
rlabel metal1 40 70 40 70 6 a1
rlabel metal1 40 70 40 70 6 a1
rlabel metal1 54 24 54 24 6 n3
rlabel ndcontact 30 20 30 20 6 n3
rlabel metal1 50 40 50 40 6 a2
rlabel metal1 50 40 50 40 6 a2
rlabel metal1 50 60 50 60 6 a1
rlabel metal1 50 60 50 60 6 a1
<< end >>
