magic
tech scmos
timestamp 1180600658
<< checkpaint >>
rect -22 -22 52 122
<< ab >>
rect 0 0 30 100
<< pwell >>
rect -4 -4 34 48
<< nwell >>
rect -4 48 34 104
<< polysilicon >>
rect 13 85 15 89
rect 13 43 15 55
rect 7 42 15 43
rect 7 38 8 42
rect 12 38 15 42
rect 7 37 15 38
rect 13 34 15 37
rect 13 10 15 14
<< ndiffusion >>
rect 3 14 13 34
rect 15 32 23 34
rect 15 28 18 32
rect 22 28 23 32
rect 15 22 23 28
rect 15 18 18 22
rect 22 18 23 22
rect 15 14 23 18
rect 3 12 11 14
rect 3 8 6 12
rect 10 8 11 12
rect 3 7 11 8
<< pdiffusion >>
rect 3 92 11 93
rect 3 88 6 92
rect 10 88 11 92
rect 3 85 11 88
rect 3 55 13 85
rect 15 82 23 85
rect 15 78 18 82
rect 22 78 23 82
rect 15 72 23 78
rect 15 68 18 72
rect 22 68 23 72
rect 15 62 23 68
rect 15 58 18 62
rect 22 58 23 62
rect 15 55 23 58
<< metal1 >>
rect -2 92 32 100
rect -2 88 6 92
rect 10 88 32 92
rect 8 42 12 83
rect 8 17 12 38
rect 18 82 22 83
rect 18 72 22 78
rect 18 62 22 68
rect 18 32 22 58
rect 18 22 22 28
rect 18 17 22 18
rect -2 8 6 12
rect 10 8 32 12
rect -2 0 32 8
<< ntransistor >>
rect 13 14 15 34
<< ptransistor >>
rect 13 55 15 85
<< polycontact >>
rect 8 38 12 42
<< ndcontact >>
rect 18 28 22 32
rect 18 18 22 22
rect 6 8 10 12
<< pdcontact >>
rect 6 88 10 92
rect 18 78 22 82
rect 18 68 22 72
rect 18 58 22 62
<< labels >>
rlabel metal1 15 6 15 6 6 vss
rlabel metal1 10 50 10 50 6 i
rlabel metal1 15 94 15 94 6 vdd
rlabel metal1 20 50 20 50 6 nq
<< end >>
