magic
tech scmos
timestamp 1179386666
<< checkpaint >>
rect -22 -25 118 105
<< ab >>
rect 0 0 96 80
<< pwell >>
rect -4 -7 100 36
<< nwell >>
rect -4 36 100 87
<< polysilicon >>
rect 9 70 11 74
rect 19 70 21 74
rect 31 70 33 74
rect 41 70 43 74
rect 53 70 55 74
rect 63 70 65 74
rect 75 70 77 74
rect 85 70 87 74
rect 9 39 11 52
rect 19 49 21 52
rect 19 48 27 49
rect 19 44 21 48
rect 25 44 27 48
rect 19 43 27 44
rect 9 38 21 39
rect 9 37 16 38
rect 15 34 16 37
rect 20 34 21 38
rect 15 33 21 34
rect 25 36 27 43
rect 31 47 33 54
rect 41 51 43 54
rect 53 51 55 54
rect 63 51 65 54
rect 41 49 55 51
rect 59 49 65 51
rect 75 49 77 56
rect 85 53 87 56
rect 83 50 87 53
rect 31 46 37 47
rect 31 42 32 46
rect 36 42 37 46
rect 31 41 37 42
rect 25 33 28 36
rect 19 30 21 33
rect 26 30 28 33
rect 33 30 35 41
rect 41 39 43 49
rect 59 45 61 49
rect 54 44 61 45
rect 54 40 55 44
rect 59 42 61 44
rect 73 48 79 49
rect 73 44 74 48
rect 78 44 79 48
rect 73 43 79 44
rect 59 40 60 42
rect 73 41 75 43
rect 54 39 60 40
rect 65 39 75 41
rect 83 39 85 50
rect 41 38 47 39
rect 41 36 42 38
rect 40 34 42 36
rect 46 35 47 38
rect 46 34 52 35
rect 40 33 52 34
rect 40 30 42 33
rect 50 30 52 33
rect 57 30 59 39
rect 65 36 67 39
rect 64 33 67 36
rect 81 38 87 39
rect 81 35 82 38
rect 71 34 82 35
rect 86 34 87 38
rect 71 33 87 34
rect 64 30 66 33
rect 71 30 73 33
rect 19 6 21 11
rect 26 6 28 11
rect 33 6 35 11
rect 40 6 42 11
rect 50 6 52 11
rect 57 6 59 11
rect 64 6 66 11
rect 71 6 73 11
<< ndiffusion >>
rect 10 15 19 30
rect 10 11 12 15
rect 16 11 19 15
rect 21 11 26 30
rect 28 11 33 30
rect 35 11 40 30
rect 42 22 50 30
rect 42 18 44 22
rect 48 18 50 22
rect 42 11 50 18
rect 52 11 57 30
rect 59 11 64 30
rect 66 11 71 30
rect 73 16 81 30
rect 73 12 75 16
rect 79 12 81 16
rect 73 11 81 12
rect 10 9 17 11
<< pdiffusion >>
rect 2 69 9 70
rect 2 65 3 69
rect 7 65 9 69
rect 2 62 9 65
rect 2 58 3 62
rect 7 58 9 62
rect 2 52 9 58
rect 11 62 19 70
rect 11 58 13 62
rect 17 58 19 62
rect 11 52 19 58
rect 21 69 31 70
rect 21 65 24 69
rect 28 65 31 69
rect 21 54 31 65
rect 33 62 41 70
rect 33 58 35 62
rect 39 58 41 62
rect 33 54 41 58
rect 43 69 53 70
rect 43 65 46 69
rect 50 65 53 69
rect 43 54 53 65
rect 55 62 63 70
rect 55 58 57 62
rect 61 58 63 62
rect 55 54 63 58
rect 65 69 75 70
rect 65 65 68 69
rect 72 65 75 69
rect 65 56 75 65
rect 77 62 85 70
rect 77 58 79 62
rect 83 58 85 62
rect 77 56 85 58
rect 87 69 94 70
rect 87 65 89 69
rect 93 65 94 69
rect 87 61 94 65
rect 87 57 89 61
rect 93 57 94 61
rect 87 56 94 57
rect 65 54 73 56
rect 21 52 29 54
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect -2 69 98 78
rect -2 68 3 69
rect 2 65 3 68
rect 7 68 24 69
rect 7 65 8 68
rect 23 65 24 68
rect 28 68 46 69
rect 28 65 29 68
rect 45 65 46 68
rect 50 68 68 69
rect 50 65 51 68
rect 67 65 68 68
rect 72 68 89 69
rect 72 65 73 68
rect 88 65 89 68
rect 93 68 98 69
rect 2 62 8 65
rect 2 58 3 62
rect 7 58 8 62
rect 12 58 13 62
rect 17 58 35 62
rect 39 58 57 62
rect 61 58 79 62
rect 83 58 84 62
rect 88 61 93 65
rect 12 55 16 58
rect 2 50 16 55
rect 88 57 89 61
rect 21 50 78 54
rect 2 22 6 50
rect 21 48 25 50
rect 17 44 21 46
rect 74 48 78 50
rect 17 42 25 44
rect 31 42 32 46
rect 36 44 63 46
rect 36 42 55 44
rect 59 40 63 44
rect 55 39 63 40
rect 15 34 16 38
rect 20 34 27 38
rect 33 34 42 38
rect 46 34 47 38
rect 57 34 63 39
rect 23 30 27 34
rect 74 33 78 44
rect 88 42 93 57
rect 82 38 86 39
rect 23 29 63 30
rect 82 29 86 34
rect 23 26 86 29
rect 57 25 86 26
rect 2 18 44 22
rect 48 18 49 22
rect 82 17 86 25
rect 75 16 79 17
rect 11 12 12 15
rect -2 11 12 12
rect 16 12 17 15
rect 16 11 98 12
rect -2 2 98 11
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
<< ntransistor >>
rect 19 11 21 30
rect 26 11 28 30
rect 33 11 35 30
rect 40 11 42 30
rect 50 11 52 30
rect 57 11 59 30
rect 64 11 66 30
rect 71 11 73 30
<< ptransistor >>
rect 9 52 11 70
rect 19 52 21 70
rect 31 54 33 70
rect 41 54 43 70
rect 53 54 55 70
rect 63 54 65 70
rect 75 56 77 70
rect 85 56 87 70
<< polycontact >>
rect 21 44 25 48
rect 16 34 20 38
rect 32 42 36 46
rect 55 40 59 44
rect 74 44 78 48
rect 42 34 46 38
rect 82 34 86 38
<< ndcontact >>
rect 12 11 16 15
rect 44 18 48 22
rect 75 12 79 16
<< pdcontact >>
rect 3 65 7 69
rect 3 58 7 62
rect 13 58 17 62
rect 24 65 28 69
rect 35 58 39 62
rect 46 65 50 69
rect 57 58 61 62
rect 68 65 72 69
rect 79 58 83 62
rect 89 65 93 69
rect 89 57 93 61
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
rect 90 -2 94 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
rect 90 78 94 82
<< psubstratepdiff >>
rect 0 2 96 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 96 2
rect 0 -3 96 -2
<< nsubstratendiff >>
rect 0 82 96 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 96 82
rect 0 77 96 78
<< labels >>
rlabel metal1 12 20 12 20 6 z
rlabel metal1 4 40 4 40 6 z
rlabel metal1 12 52 12 52 6 z
rlabel metal1 20 20 20 20 6 z
rlabel metal1 28 20 28 20 6 z
rlabel metal1 28 28 28 28 6 a
rlabel metal1 20 36 20 36 6 a
rlabel metal1 20 44 20 44 6 b
rlabel metal1 28 52 28 52 6 b
rlabel metal1 20 60 20 60 6 z
rlabel metal1 28 60 28 60 6 z
rlabel metal1 48 6 48 6 6 vss
rlabel metal1 36 20 36 20 6 z
rlabel metal1 36 28 36 28 6 a
rlabel metal1 44 20 44 20 6 z
rlabel metal1 44 28 44 28 6 a
rlabel metal1 52 28 52 28 6 a
rlabel metal1 36 36 36 36 6 d
rlabel metal1 36 44 36 44 6 c
rlabel polycontact 44 36 44 36 6 d
rlabel metal1 44 44 44 44 6 c
rlabel metal1 52 44 52 44 6 c
rlabel metal1 44 52 44 52 6 b
rlabel metal1 52 52 52 52 6 b
rlabel metal1 36 52 36 52 6 b
rlabel pdcontact 36 60 36 60 6 z
rlabel metal1 44 60 44 60 6 z
rlabel metal1 52 60 52 60 6 z
rlabel metal1 48 74 48 74 6 vdd
rlabel metal1 60 28 60 28 6 a
rlabel metal1 60 40 60 40 6 c
rlabel metal1 76 40 76 40 6 b
rlabel metal1 68 52 68 52 6 b
rlabel metal1 60 52 60 52 6 b
rlabel pdcontact 60 60 60 60 6 z
rlabel metal1 68 60 68 60 6 z
rlabel metal1 76 60 76 60 6 z
rlabel metal1 84 28 84 28 6 a
<< end >>
