magic
tech scmos
timestamp 1179386575
<< checkpaint >>
rect -22 -22 158 94
<< ab >>
rect 0 0 136 72
<< pwell >>
rect -4 -4 140 32
<< nwell >>
rect -4 32 140 76
<< polysilicon >>
rect 9 66 11 70
rect 19 66 21 70
rect 29 66 31 70
rect 39 66 41 70
rect 49 66 51 70
rect 59 66 61 70
rect 69 66 71 70
rect 79 66 81 70
rect 89 66 91 70
rect 99 66 101 70
rect 109 66 111 70
rect 119 57 121 61
rect 9 35 11 44
rect 19 43 21 46
rect 19 42 25 43
rect 19 38 20 42
rect 24 38 25 42
rect 19 37 25 38
rect 9 34 15 35
rect 9 30 10 34
rect 14 32 15 34
rect 14 30 17 32
rect 9 29 17 30
rect 15 26 17 29
rect 22 26 24 37
rect 29 35 31 46
rect 39 35 41 46
rect 49 43 51 46
rect 45 42 51 43
rect 45 38 46 42
rect 50 38 51 42
rect 45 37 51 38
rect 29 34 41 35
rect 29 30 36 34
rect 40 30 41 34
rect 29 29 41 30
rect 29 26 31 29
rect 39 26 41 29
rect 46 26 48 37
rect 59 31 61 46
rect 69 31 71 46
rect 79 43 81 46
rect 79 42 85 43
rect 79 38 80 42
rect 84 38 85 42
rect 79 37 85 38
rect 53 29 77 31
rect 53 26 55 29
rect 62 26 68 29
rect 75 26 77 29
rect 82 26 84 37
rect 89 35 91 46
rect 99 35 101 46
rect 109 42 111 46
rect 105 41 111 42
rect 105 37 106 41
rect 110 37 111 41
rect 105 36 111 37
rect 89 34 101 35
rect 89 30 91 34
rect 95 30 101 34
rect 89 29 101 30
rect 89 26 91 29
rect 99 26 101 29
rect 106 26 108 36
rect 119 35 121 39
rect 119 34 127 35
rect 119 31 122 34
rect 113 30 122 31
rect 126 30 127 34
rect 113 29 127 30
rect 113 26 115 29
rect 62 22 63 26
rect 67 22 68 26
rect 62 21 68 22
rect 15 2 17 6
rect 22 2 24 6
rect 29 2 31 6
rect 39 2 41 6
rect 46 2 48 6
rect 53 2 55 6
rect 75 2 77 6
rect 82 2 84 6
rect 89 2 91 6
rect 99 2 101 6
rect 106 2 108 6
rect 113 2 115 6
<< ndiffusion >>
rect 7 11 15 26
rect 7 7 9 11
rect 13 7 15 11
rect 7 6 15 7
rect 17 6 22 26
rect 24 6 29 26
rect 31 18 39 26
rect 31 14 33 18
rect 37 14 39 18
rect 31 6 39 14
rect 41 6 46 26
rect 48 6 53 26
rect 55 18 60 26
rect 70 18 75 26
rect 55 11 75 18
rect 55 7 57 11
rect 61 7 69 11
rect 73 7 75 11
rect 55 6 75 7
rect 77 6 82 26
rect 84 6 89 26
rect 91 18 99 26
rect 91 14 93 18
rect 97 14 99 18
rect 91 6 99 14
rect 101 6 106 26
rect 108 6 113 26
rect 115 18 123 26
rect 115 14 117 18
rect 121 14 123 18
rect 115 11 123 14
rect 115 7 117 11
rect 121 7 123 11
rect 115 6 123 7
<< pdiffusion >>
rect 2 65 9 66
rect 2 61 3 65
rect 7 61 9 65
rect 2 58 9 61
rect 2 54 3 58
rect 7 54 9 58
rect 2 44 9 54
rect 11 58 19 66
rect 11 54 13 58
rect 17 54 19 58
rect 11 51 19 54
rect 11 47 13 51
rect 17 47 19 51
rect 11 46 19 47
rect 21 65 29 66
rect 21 61 23 65
rect 27 61 29 65
rect 21 58 29 61
rect 21 54 23 58
rect 27 54 29 58
rect 21 46 29 54
rect 31 58 39 66
rect 31 54 33 58
rect 37 54 39 58
rect 31 51 39 54
rect 31 47 33 51
rect 37 47 39 51
rect 31 46 39 47
rect 41 65 49 66
rect 41 61 43 65
rect 47 61 49 65
rect 41 58 49 61
rect 41 54 43 58
rect 47 54 49 58
rect 41 46 49 54
rect 51 58 59 66
rect 51 54 53 58
rect 57 54 59 58
rect 51 51 59 54
rect 51 47 53 51
rect 57 47 59 51
rect 51 46 59 47
rect 61 65 69 66
rect 61 61 63 65
rect 67 61 69 65
rect 61 58 69 61
rect 61 54 63 58
rect 67 54 69 58
rect 61 46 69 54
rect 71 58 79 66
rect 71 54 73 58
rect 77 54 79 58
rect 71 51 79 54
rect 71 47 73 51
rect 77 47 79 51
rect 71 46 79 47
rect 81 65 89 66
rect 81 61 83 65
rect 87 61 89 65
rect 81 58 89 61
rect 81 54 83 58
rect 87 54 89 58
rect 81 46 89 54
rect 91 58 99 66
rect 91 54 93 58
rect 97 54 99 58
rect 91 51 99 54
rect 91 47 93 51
rect 97 47 99 51
rect 91 46 99 47
rect 101 65 109 66
rect 101 61 103 65
rect 107 61 109 65
rect 101 58 109 61
rect 101 54 103 58
rect 107 54 109 58
rect 101 46 109 54
rect 111 57 116 66
rect 111 54 119 57
rect 111 50 113 54
rect 117 50 119 54
rect 111 46 119 50
rect 11 44 16 46
rect 114 39 119 46
rect 121 56 129 57
rect 121 52 124 56
rect 128 52 129 56
rect 121 49 129 52
rect 121 45 124 49
rect 128 45 129 49
rect 121 39 129 45
<< metal1 >>
rect -2 68 138 72
rect -2 65 125 68
rect -2 64 3 65
rect 2 61 3 64
rect 7 64 23 65
rect 7 61 8 64
rect 2 58 8 61
rect 22 61 23 64
rect 27 64 43 65
rect 27 61 28 64
rect 2 54 3 58
rect 7 54 8 58
rect 13 58 17 59
rect 22 58 28 61
rect 42 61 43 64
rect 47 64 63 65
rect 47 61 48 64
rect 22 54 23 58
rect 27 54 28 58
rect 33 58 38 59
rect 37 54 38 58
rect 42 58 48 61
rect 62 61 63 64
rect 67 64 83 65
rect 67 61 68 64
rect 42 54 43 58
rect 47 54 48 58
rect 53 58 57 59
rect 62 58 68 61
rect 82 61 83 64
rect 87 64 103 65
rect 87 61 88 64
rect 62 54 63 58
rect 67 54 68 58
rect 73 58 78 59
rect 77 54 78 58
rect 82 58 88 61
rect 102 61 103 64
rect 107 64 125 65
rect 129 64 138 68
rect 107 61 108 64
rect 82 54 83 58
rect 87 54 88 58
rect 93 58 97 59
rect 102 58 108 61
rect 102 54 103 58
rect 107 54 108 58
rect 113 54 119 59
rect 13 51 17 54
rect 2 47 13 50
rect 33 51 38 54
rect 17 47 33 50
rect 37 50 38 51
rect 53 51 57 54
rect 37 47 53 50
rect 73 51 78 54
rect 57 47 73 50
rect 77 50 78 51
rect 93 51 97 54
rect 77 47 93 50
rect 117 50 119 54
rect 97 47 119 50
rect 2 46 119 47
rect 123 56 129 64
rect 123 52 124 56
rect 128 52 129 56
rect 123 49 129 52
rect 2 18 6 46
rect 123 45 124 49
rect 128 45 129 49
rect 19 38 20 42
rect 24 38 46 42
rect 50 38 80 42
rect 84 41 119 42
rect 84 38 106 41
rect 105 37 106 38
rect 110 38 119 41
rect 110 37 111 38
rect 10 34 14 35
rect 33 30 36 34
rect 40 30 91 34
rect 95 30 96 34
rect 105 30 111 37
rect 121 30 122 34
rect 126 30 127 34
rect 10 26 14 30
rect 121 26 127 30
rect 10 22 63 26
rect 67 22 127 26
rect 2 14 33 18
rect 37 14 93 18
rect 97 14 103 18
rect 116 14 117 18
rect 121 14 122 18
rect 116 11 122 14
rect 8 8 9 11
rect -2 7 9 8
rect 13 8 14 11
rect 56 8 57 11
rect 13 7 57 8
rect 61 8 62 11
rect 68 8 69 11
rect 61 7 69 8
rect 73 8 74 11
rect 116 8 117 11
rect 73 7 117 8
rect 121 8 122 11
rect 121 7 128 8
rect -2 4 128 7
rect 132 4 138 8
rect -2 0 138 4
<< ntransistor >>
rect 15 6 17 26
rect 22 6 24 26
rect 29 6 31 26
rect 39 6 41 26
rect 46 6 48 26
rect 53 6 55 26
rect 75 6 77 26
rect 82 6 84 26
rect 89 6 91 26
rect 99 6 101 26
rect 106 6 108 26
rect 113 6 115 26
<< ptransistor >>
rect 9 44 11 66
rect 19 46 21 66
rect 29 46 31 66
rect 39 46 41 66
rect 49 46 51 66
rect 59 46 61 66
rect 69 46 71 66
rect 79 46 81 66
rect 89 46 91 66
rect 99 46 101 66
rect 109 46 111 66
rect 119 39 121 57
<< polycontact >>
rect 20 38 24 42
rect 10 30 14 34
rect 46 38 50 42
rect 36 30 40 34
rect 80 38 84 42
rect 106 37 110 41
rect 91 30 95 34
rect 122 30 126 34
rect 63 22 67 26
<< ndcontact >>
rect 9 7 13 11
rect 33 14 37 18
rect 57 7 61 11
rect 69 7 73 11
rect 93 14 97 18
rect 117 14 121 18
rect 117 7 121 11
<< pdcontact >>
rect 3 61 7 65
rect 3 54 7 58
rect 13 54 17 58
rect 13 47 17 51
rect 23 61 27 65
rect 23 54 27 58
rect 33 54 37 58
rect 33 47 37 51
rect 43 61 47 65
rect 43 54 47 58
rect 53 54 57 58
rect 53 47 57 51
rect 63 61 67 65
rect 63 54 67 58
rect 73 54 77 58
rect 73 47 77 51
rect 83 61 87 65
rect 83 54 87 58
rect 93 54 97 58
rect 93 47 97 51
rect 103 61 107 65
rect 103 54 107 58
rect 113 50 117 54
rect 124 52 128 56
rect 124 45 128 49
<< psubstratepcontact >>
rect 128 4 132 8
<< nsubstratencontact >>
rect 125 64 129 68
<< psubstratepdiff >>
rect 127 8 133 24
rect 127 4 128 8
rect 132 4 133 8
rect 127 3 133 4
<< nsubstratendiff >>
rect 121 68 133 69
rect 121 64 125 68
rect 129 64 133 68
rect 121 63 133 64
<< labels >>
rlabel metal1 12 16 12 16 6 z
rlabel metal1 4 32 4 32 6 z
rlabel polycontact 12 32 12 32 6 a
rlabel metal1 12 48 12 48 6 z
rlabel metal1 20 16 20 16 6 z
rlabel metal1 28 16 28 16 6 z
rlabel ndcontact 36 16 36 16 6 z
rlabel metal1 28 24 28 24 6 a
rlabel metal1 36 24 36 24 6 a
rlabel metal1 20 24 20 24 6 a
rlabel metal1 36 32 36 32 6 c
rlabel metal1 28 40 28 40 6 b
rlabel metal1 36 40 36 40 6 b
rlabel metal1 28 48 28 48 6 z
rlabel metal1 36 52 36 52 6 z
rlabel metal1 20 48 20 48 6 z
rlabel metal1 44 16 44 16 6 z
rlabel metal1 52 16 52 16 6 z
rlabel metal1 60 16 60 16 6 z
rlabel metal1 52 24 52 24 6 a
rlabel metal1 60 24 60 24 6 a
rlabel metal1 44 24 44 24 6 a
rlabel metal1 44 32 44 32 6 c
rlabel metal1 52 32 52 32 6 c
rlabel metal1 60 32 60 32 6 c
rlabel metal1 52 40 52 40 6 b
rlabel metal1 60 40 60 40 6 b
rlabel metal1 44 40 44 40 6 b
rlabel metal1 52 48 52 48 6 z
rlabel metal1 60 48 60 48 6 z
rlabel metal1 44 48 44 48 6 z
rlabel metal1 68 4 68 4 6 vss
rlabel metal1 68 16 68 16 6 z
rlabel metal1 76 16 76 16 6 z
rlabel metal1 84 16 84 16 6 z
rlabel metal1 76 24 76 24 6 a
rlabel metal1 84 24 84 24 6 a
rlabel metal1 68 24 68 24 6 a
rlabel metal1 68 32 68 32 6 c
rlabel metal1 76 32 76 32 6 c
rlabel metal1 84 32 84 32 6 c
rlabel metal1 76 40 76 40 6 b
rlabel metal1 84 40 84 40 6 b
rlabel metal1 68 40 68 40 6 b
rlabel metal1 76 52 76 52 6 z
rlabel metal1 84 48 84 48 6 z
rlabel metal1 68 48 68 48 6 z
rlabel metal1 68 68 68 68 6 vdd
rlabel metal1 92 16 92 16 6 z
rlabel metal1 100 16 100 16 6 z
rlabel metal1 100 24 100 24 6 a
rlabel metal1 108 24 108 24 6 a
rlabel metal1 92 24 92 24 6 a
rlabel polycontact 92 32 92 32 6 c
rlabel metal1 100 40 100 40 6 b
rlabel metal1 108 36 108 36 6 b
rlabel metal1 92 40 92 40 6 b
rlabel metal1 100 48 100 48 6 z
rlabel metal1 108 48 108 48 6 z
rlabel metal1 92 48 92 48 6 z
rlabel metal1 124 28 124 28 6 a
rlabel metal1 116 24 116 24 6 a
rlabel metal1 116 40 116 40 6 b
rlabel pdcontact 116 52 116 52 6 z
<< end >>
