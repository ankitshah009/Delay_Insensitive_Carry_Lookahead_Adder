magic
tech scmos
timestamp 1179385117
<< checkpaint >>
rect -22 -25 78 105
<< ab >>
rect 0 0 56 80
<< pwell >>
rect -4 -7 60 36
<< nwell >>
rect -4 36 60 87
<< polysilicon >>
rect 9 64 11 69
rect 19 64 21 69
rect 29 64 31 69
rect 41 63 47 64
rect 41 59 42 63
rect 46 59 47 63
rect 41 58 47 59
rect 41 55 43 58
rect 9 31 11 53
rect 19 47 21 53
rect 15 46 21 47
rect 15 42 16 46
rect 20 42 21 46
rect 15 41 21 42
rect 8 30 14 31
rect 8 26 9 30
rect 13 26 14 30
rect 8 25 14 26
rect 12 22 14 25
rect 19 22 21 41
rect 29 31 31 53
rect 25 30 31 31
rect 41 30 43 43
rect 25 26 26 30
rect 30 26 31 30
rect 25 25 31 26
rect 26 22 28 25
rect 41 21 43 24
rect 41 20 47 21
rect 41 16 42 20
rect 46 16 47 20
rect 41 15 47 16
rect 12 6 14 11
rect 19 6 21 11
rect 26 6 28 11
<< ndiffusion >>
rect 33 24 41 30
rect 43 29 50 30
rect 43 25 45 29
rect 49 25 50 29
rect 43 24 50 25
rect 33 22 39 24
rect 5 21 12 22
rect 5 17 6 21
rect 10 17 12 21
rect 5 16 12 17
rect 7 11 12 16
rect 14 11 19 22
rect 21 11 26 22
rect 28 12 39 22
rect 28 11 33 12
rect 30 8 33 11
rect 37 8 39 12
rect 30 7 39 8
<< pdiffusion >>
rect 33 72 39 73
rect 33 68 34 72
rect 38 68 39 72
rect 33 64 39 68
rect 4 59 9 64
rect 2 58 9 59
rect 2 54 3 58
rect 7 54 9 58
rect 2 53 9 54
rect 11 63 19 64
rect 11 59 13 63
rect 17 59 19 63
rect 11 53 19 59
rect 21 60 29 64
rect 21 56 23 60
rect 27 56 29 60
rect 21 53 29 56
rect 31 55 39 64
rect 31 53 41 55
rect 33 43 41 53
rect 43 49 48 55
rect 43 48 50 49
rect 43 44 45 48
rect 49 44 50 48
rect 43 43 50 44
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect -2 72 58 78
rect -2 68 34 72
rect 38 68 58 72
rect 12 63 18 68
rect 12 59 13 63
rect 17 59 18 63
rect 23 60 42 63
rect 3 58 7 59
rect 27 59 42 60
rect 46 59 47 63
rect 23 55 27 56
rect 7 54 27 55
rect 3 51 27 54
rect 34 49 46 55
rect 42 48 49 49
rect 2 31 6 47
rect 10 46 30 47
rect 10 42 16 46
rect 20 42 30 46
rect 10 41 30 42
rect 42 44 45 48
rect 42 43 49 44
rect 18 33 22 41
rect 34 31 38 39
rect 2 30 14 31
rect 2 26 9 30
rect 13 26 14 30
rect 2 25 14 26
rect 26 30 38 31
rect 30 26 38 30
rect 26 25 38 26
rect 42 29 46 43
rect 42 25 45 29
rect 49 25 50 29
rect 5 17 6 21
rect 10 20 47 21
rect 10 17 42 20
rect 41 16 42 17
rect 46 16 47 20
rect -2 8 33 12
rect 37 8 58 12
rect -2 2 58 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
<< ntransistor >>
rect 41 24 43 30
rect 12 11 14 22
rect 19 11 21 22
rect 26 11 28 22
<< ptransistor >>
rect 9 53 11 64
rect 19 53 21 64
rect 29 53 31 64
rect 41 43 43 55
<< polycontact >>
rect 42 59 46 63
rect 16 42 20 46
rect 9 26 13 30
rect 26 26 30 30
rect 42 16 46 20
<< ndcontact >>
rect 45 25 49 29
rect 6 17 10 21
rect 33 8 37 12
<< pdcontact >>
rect 34 68 38 72
rect 3 54 7 58
rect 13 59 17 63
rect 23 56 27 60
rect 45 44 49 48
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
<< psubstratepdiff >>
rect 0 2 56 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 56 2
rect 0 -3 56 -2
<< nsubstratendiff >>
rect 0 82 56 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 56 82
rect 0 77 56 78
<< labels >>
rlabel polycontact 44 18 44 18 6 zn
rlabel polycontact 44 61 44 61 6 zn
rlabel metal1 4 36 4 36 6 c
rlabel polycontact 12 28 12 28 6 c
rlabel metal1 20 40 20 40 6 b
rlabel metal1 12 44 12 44 6 b
rlabel metal1 15 53 15 53 6 zn
rlabel pdcontact 25 57 25 57 6 zn
rlabel metal1 28 6 28 6 6 vss
rlabel polycontact 28 28 28 28 6 a
rlabel metal1 36 32 36 32 6 a
rlabel metal1 28 44 28 44 6 b
rlabel metal1 36 52 36 52 6 z
rlabel metal1 28 74 28 74 6 vdd
rlabel metal1 26 19 26 19 6 zn
rlabel metal1 44 40 44 40 6 z
rlabel metal1 35 61 35 61 6 zn
<< end >>
