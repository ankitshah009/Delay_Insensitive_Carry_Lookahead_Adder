.subckt xor2v2x1 a b vdd vss z
*   SPICE3 file   created from xor2v2x1.ext -      technology: scmos
m00 z      bn     an     vdd p w=28u  l=2.3636u ad=112p     pd=36u      as=132p     ps=57u
m01 bn     an     z      vdd p w=28u  l=2.3636u ad=112p     pd=36u      as=112p     ps=36u
m02 vdd    b      bn     vdd p w=28u  l=2.3636u ad=161p     pd=58u      as=112p     ps=36u
m03 an     a      vdd    vdd p w=14u  l=2.3636u ad=66p      pd=28.5u    as=80.5p    ps=29u
m04 vdd    a      an     vdd p w=14u  l=2.3636u ad=80.5p    pd=29u      as=66p      ps=28.5u
m05 w1     bn     z      vss n w=19u  l=2.3636u ad=47.5p    pd=24u      as=88.5319p ps=38.8085u
m06 vss    an     w1     vss n w=19u  l=2.3636u ad=137.606p pd=54.1212u as=47.5p    ps=24u
m07 bn     b      vss    vss n w=7u   l=2.3636u ad=30.3333p pd=14.6667u as=50.697p  ps=19.9394u
m08 z      a      bn     vss n w=14u  l=2.3636u ad=65.234p  pd=28.5957u as=60.6667p ps=29.3333u
m09 an     b      z      vss n w=14u  l=2.3636u ad=60.6667p pd=29.3333u as=65.234p  ps=28.5957u
m10 vss    a      an     vss n w=7u   l=2.3636u ad=50.697p  pd=19.9394u as=30.3333p ps=14.6667u
C0  vdd    an     0.390f
C1  z      bn     0.550f
C2  a      b      0.184f
C3  a      bn     0.033f
C4  b      an     0.221f
C5  vss    z      0.280f
C6  an     bn     0.586f
C7  vss    a      0.015f
C8  z      a      0.027f
C9  vss    an     0.100f
C10 w1     bn     0.007f
C11 z      an     0.371f
C12 vdd    b      0.027f
C13 vdd    bn     0.060f
C14 a      an     0.174f
C15 vss    w1     0.004f
C16 b      bn     0.040f
C17 w1     z      0.010f
C18 vss    vdd    0.003f
C19 z      vdd    0.047f
C20 vss    b      0.066f
C21 vdd    a      0.049f
C22 vss    bn     0.102f
C23 z      b      0.006f
C25 z      vss    0.016f
C27 a      vss    0.049f
C28 b      vss    0.047f
C29 an     vss    0.026f
C30 bn     vss    0.016f
.ends
