magic
tech scmos
timestamp 1179384953
<< checkpaint >>
rect -22 -25 62 105
<< ab >>
rect 0 0 40 80
<< pwell >>
rect -4 -7 44 36
<< nwell >>
rect -4 36 44 87
<< polysilicon >>
rect 19 62 25 63
rect 9 54 11 59
rect 19 58 20 62
rect 24 58 25 62
rect 19 57 25 58
rect 19 52 21 57
rect 29 52 31 57
rect 9 39 11 42
rect 19 39 21 42
rect 9 38 15 39
rect 9 34 10 38
rect 14 34 15 38
rect 19 36 23 39
rect 9 33 15 34
rect 9 25 11 33
rect 21 22 23 36
rect 29 31 31 42
rect 28 30 34 31
rect 28 26 29 30
rect 33 26 34 30
rect 28 25 34 26
rect 28 22 30 25
rect 9 15 11 19
rect 21 8 23 13
rect 28 8 30 13
<< ndiffusion >>
rect 2 24 9 25
rect 2 20 3 24
rect 7 20 9 24
rect 2 19 9 20
rect 11 22 19 25
rect 11 19 21 22
rect 13 13 21 19
rect 23 13 28 22
rect 30 21 37 22
rect 30 17 32 21
rect 36 17 37 21
rect 30 16 37 17
rect 30 13 35 16
rect 13 12 19 13
rect 13 8 14 12
rect 18 8 19 12
rect 13 7 19 8
<< pdiffusion >>
rect 4 48 9 54
rect 2 47 9 48
rect 2 43 3 47
rect 7 43 9 47
rect 2 42 9 43
rect 11 52 17 54
rect 11 47 19 52
rect 11 43 13 47
rect 17 43 19 47
rect 11 42 19 43
rect 21 47 29 52
rect 21 43 23 47
rect 27 43 29 47
rect 21 42 29 43
rect 31 51 38 52
rect 31 47 33 51
rect 37 47 38 51
rect 31 42 38 47
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect -2 68 42 78
rect 2 48 6 55
rect 2 47 7 48
rect 2 43 3 47
rect 10 47 14 68
rect 17 62 30 63
rect 17 58 20 62
rect 24 58 30 62
rect 17 57 30 58
rect 17 50 23 57
rect 33 51 37 68
rect 10 43 13 47
rect 17 43 18 47
rect 22 43 23 47
rect 27 43 28 47
rect 33 46 37 47
rect 2 42 7 43
rect 2 25 6 42
rect 22 38 28 43
rect 9 34 10 38
rect 14 34 28 38
rect 2 24 7 25
rect 2 20 3 24
rect 7 20 14 23
rect 2 17 14 20
rect 18 21 22 34
rect 34 30 38 39
rect 25 26 29 30
rect 33 26 38 30
rect 25 25 38 26
rect 18 17 32 21
rect 36 17 37 21
rect -2 8 14 12
rect 18 8 42 12
rect -2 2 42 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
<< ntransistor >>
rect 9 19 11 25
rect 21 13 23 22
rect 28 13 30 22
<< ptransistor >>
rect 9 42 11 54
rect 19 42 21 52
rect 29 42 31 52
<< polycontact >>
rect 20 58 24 62
rect 10 34 14 38
rect 29 26 33 30
<< ndcontact >>
rect 3 20 7 24
rect 32 17 36 21
rect 14 8 18 12
<< pdcontact >>
rect 3 43 7 47
rect 13 43 17 47
rect 23 43 27 47
rect 33 47 37 51
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
<< psubstratepdiff >>
rect 0 2 40 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 40 2
rect 0 -3 40 -2
<< nsubstratendiff >>
rect 0 82 40 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 40 82
rect 0 77 40 78
<< labels >>
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 20 12 20 6 z
rlabel metal1 20 6 20 6 6 vss
rlabel metal1 18 36 18 36 6 zn
rlabel metal1 28 28 28 28 6 b
rlabel metal1 25 40 25 40 6 zn
rlabel metal1 20 56 20 56 6 a
rlabel metal1 28 60 28 60 6 a
rlabel metal1 20 74 20 74 6 vdd
rlabel metal1 27 19 27 19 6 zn
rlabel metal1 36 32 36 32 6 b
<< end >>
