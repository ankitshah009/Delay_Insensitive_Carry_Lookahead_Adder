magic
tech scmos
timestamp 1179386374
<< checkpaint >>
rect -22 -25 86 105
<< ab >>
rect 0 0 64 80
<< pwell >>
rect -4 -7 68 36
<< nwell >>
rect -4 36 68 87
<< polysilicon >>
rect 9 65 11 70
rect 19 65 21 70
rect 29 65 31 70
rect 39 65 41 70
rect 9 45 11 48
rect 9 44 15 45
rect 9 40 10 44
rect 14 40 15 44
rect 9 39 15 40
rect 19 39 21 48
rect 29 39 31 48
rect 10 30 12 39
rect 19 38 31 39
rect 19 35 26 38
rect 17 34 26 35
rect 30 34 31 38
rect 39 39 41 48
rect 39 38 48 39
rect 39 35 42 38
rect 17 33 31 34
rect 17 30 19 33
rect 29 30 31 33
rect 36 34 42 35
rect 46 34 48 38
rect 36 33 48 34
rect 36 30 38 33
rect 46 30 48 33
rect 53 38 59 39
rect 53 34 54 38
rect 58 34 59 38
rect 53 33 59 34
rect 53 30 55 33
rect 10 8 12 13
rect 17 8 19 13
rect 29 6 31 10
rect 36 6 38 10
rect 46 6 48 10
rect 53 6 55 10
<< ndiffusion >>
rect 3 29 10 30
rect 3 25 4 29
rect 8 25 10 29
rect 3 22 10 25
rect 3 18 4 22
rect 8 18 10 22
rect 3 17 10 18
rect 5 13 10 17
rect 12 13 17 30
rect 19 15 29 30
rect 19 13 22 15
rect 21 11 22 13
rect 26 11 29 15
rect 21 10 29 11
rect 31 10 36 30
rect 38 22 46 30
rect 38 18 40 22
rect 44 18 46 22
rect 38 10 46 18
rect 48 10 53 30
rect 55 22 62 30
rect 55 18 57 22
rect 61 18 62 22
rect 55 15 62 18
rect 55 11 57 15
rect 61 11 62 15
rect 55 10 62 11
<< pdiffusion >>
rect 2 64 9 65
rect 2 60 3 64
rect 7 60 9 64
rect 2 48 9 60
rect 11 62 19 65
rect 11 58 13 62
rect 17 58 19 62
rect 11 54 19 58
rect 11 50 13 54
rect 17 50 19 54
rect 11 48 19 50
rect 21 64 29 65
rect 21 60 23 64
rect 27 60 29 64
rect 21 48 29 60
rect 31 62 39 65
rect 31 58 33 62
rect 37 58 39 62
rect 31 54 39 58
rect 31 50 33 54
rect 37 50 39 54
rect 31 48 39 50
rect 41 64 49 65
rect 41 60 43 64
rect 47 60 49 64
rect 41 56 49 60
rect 41 52 43 56
rect 47 52 49 56
rect 41 48 49 52
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect -2 68 66 78
rect 3 64 7 68
rect 23 64 27 68
rect 3 59 7 60
rect 13 62 17 63
rect 43 64 47 68
rect 23 59 27 60
rect 33 62 38 63
rect 13 54 17 58
rect 37 58 38 62
rect 33 54 38 58
rect 2 50 13 54
rect 17 50 33 54
rect 37 50 38 54
rect 43 56 47 60
rect 43 51 47 52
rect 2 30 6 50
rect 10 44 21 45
rect 14 40 21 44
rect 10 39 21 40
rect 17 30 21 39
rect 25 42 55 46
rect 25 38 31 42
rect 51 38 55 42
rect 25 34 26 38
rect 30 34 31 38
rect 41 34 42 38
rect 46 34 47 38
rect 51 34 54 38
rect 58 34 59 38
rect 41 30 47 34
rect 2 29 8 30
rect 2 25 4 29
rect 17 26 47 30
rect 2 22 8 25
rect 2 18 4 22
rect 8 18 40 22
rect 44 18 47 22
rect 56 18 57 22
rect 61 18 62 22
rect 56 15 62 18
rect 21 12 22 15
rect -2 11 22 12
rect 26 12 27 15
rect 56 12 57 15
rect 26 11 57 12
rect 61 12 62 15
rect 61 11 66 12
rect -2 2 66 11
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
<< ntransistor >>
rect 10 13 12 30
rect 17 13 19 30
rect 29 10 31 30
rect 36 10 38 30
rect 46 10 48 30
rect 53 10 55 30
<< ptransistor >>
rect 9 48 11 65
rect 19 48 21 65
rect 29 48 31 65
rect 39 48 41 65
<< polycontact >>
rect 10 40 14 44
rect 26 34 30 38
rect 42 34 46 38
rect 54 34 58 38
<< ndcontact >>
rect 4 25 8 29
rect 4 18 8 22
rect 22 11 26 15
rect 40 18 44 22
rect 57 18 61 22
rect 57 11 61 15
<< pdcontact >>
rect 3 60 7 64
rect 13 58 17 62
rect 13 50 17 54
rect 23 60 27 64
rect 33 58 37 62
rect 33 50 37 54
rect 43 60 47 64
rect 43 52 47 56
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
<< psubstratepdiff >>
rect 0 2 64 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 64 2
rect 0 -3 64 -2
<< nsubstratendiff >>
rect 0 82 64 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 64 82
rect 0 77 64 78
<< labels >>
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 20 12 20 6 z
rlabel metal1 20 20 20 20 6 z
rlabel metal1 20 28 20 28 6 b
rlabel metal1 20 52 20 52 6 z
rlabel metal1 12 52 12 52 6 z
rlabel metal1 32 6 32 6 6 vss
rlabel metal1 28 20 28 20 6 z
rlabel metal1 28 28 28 28 6 b
rlabel metal1 36 20 36 20 6 z
rlabel metal1 36 28 36 28 6 b
rlabel metal1 28 40 28 40 6 a
rlabel metal1 36 44 36 44 6 a
rlabel metal1 28 52 28 52 6 z
rlabel pdcontact 36 60 36 60 6 z
rlabel metal1 32 74 32 74 6 vdd
rlabel metal1 44 20 44 20 6 z
rlabel metal1 44 32 44 32 6 b
rlabel metal1 44 44 44 44 6 a
rlabel metal1 52 44 52 44 6 a
<< end >>
