.subckt nr2v0x2 a b vdd vss z
*   SPICE3 file   created from nr2v0x2.ext -      technology: scmos
m00 w1     a      vdd    vdd p w=27u  l=2.3636u ad=67.5p    pd=32u      as=189p     ps=68u
m01 z      b      w1     vdd p w=27u  l=2.3636u ad=108p     pd=35u      as=67.5p    ps=32u
m02 w2     b      z      vdd p w=27u  l=2.3636u ad=67.5p    pd=32u      as=108p     ps=35u
m03 vdd    a      w2     vdd p w=27u  l=2.3636u ad=189p     pd=68u      as=67.5p    ps=32u
m04 z      a      vss    vss n w=15u  l=2.3636u ad=60p      pd=23u      as=120p     ps=46u
m05 vss    b      z      vss n w=15u  l=2.3636u ad=120p     pd=46u      as=60p      ps=23u
C0  z      vdd    0.062f
C1  b      vdd    0.039f
C2  z      w1     0.006f
C3  vss    a      0.152f
C4  z      a      0.160f
C5  w2     vdd    0.005f
C6  b      a      0.306f
C7  w1     vdd    0.005f
C8  a      vdd    0.030f
C9  vss    z      0.196f
C10 vss    b      0.034f
C11 vss    vdd    0.003f
C12 z      b      0.058f
C14 z      vss    0.011f
C15 b      vss    0.030f
C16 a      vss    0.044f
.ends
