.subckt nr2av0x1 a b vdd vss z
*   SPICE3 file   created from nr2av0x1.ext -      technology: scmos
m00 w1     b      z      vdd p w=28u  l=2.3636u ad=70p      pd=33u      as=166p     ps=70u
m01 vdd    an     w1     vdd p w=28u  l=2.3636u ad=198.545p pd=50.9091u as=70p      ps=33u
m02 an     a      vdd    vdd p w=16u  l=2.3636u ad=106p     pd=46u      as=113.455p ps=29.0909u
m03 an     a      vss    vss n w=8u   l=2.3636u ad=52p      pd=30u      as=72.6667p ps=32.6667u
m04 z      b      vss    vss n w=8u   l=2.3636u ad=32p      pd=16u      as=72.6667p ps=32.6667u
m05 vss    an     z      vss n w=8u   l=2.3636u ad=72.6667p pd=32.6667u as=32p      ps=16u
C0  vdd    an     0.045f
C1  z      b      0.190f
C2  an     b      0.140f
C3  a      z      0.041f
C4  vss    vdd    0.004f
C5  vss    b      0.017f
C6  w1     vdd    0.005f
C7  a      an     0.240f
C8  z      an     0.084f
C9  w1     b      0.016f
C10 vdd    b      0.057f
C11 vss    a      0.027f
C12 vss    z      0.188f
C13 w1     z      0.003f
C14 a      vdd    0.049f
C15 vss    an     0.090f
C16 z      vdd    0.088f
C17 a      b      0.128f
C19 a      vss    0.022f
C20 z      vss    0.016f
C22 an     vss    0.025f
C23 b      vss    0.018f
.ends
