magic
tech scmos
timestamp 1179385938
<< checkpaint >>
rect -22 -22 46 94
<< ab >>
rect 0 0 24 72
<< pwell >>
rect -4 -4 28 32
<< nwell >>
rect -4 32 28 76
<< polysilicon >>
rect 9 62 11 67
rect 9 35 11 38
rect 9 34 15 35
rect 9 30 10 34
rect 14 30 15 34
rect 9 29 15 30
rect 9 25 11 29
rect 9 14 11 19
<< ndiffusion >>
rect 2 24 9 25
rect 2 20 3 24
rect 7 20 9 24
rect 2 19 9 20
rect 11 19 19 25
rect 13 18 19 19
rect 13 14 14 18
rect 18 14 19 18
rect 13 13 19 14
<< pdiffusion >>
rect 2 61 9 62
rect 2 57 3 61
rect 7 57 9 61
rect 2 38 9 57
rect 11 51 16 62
rect 11 50 18 51
rect 11 46 13 50
rect 17 46 18 50
rect 11 43 18 46
rect 11 39 13 43
rect 17 39 18 43
rect 11 38 18 39
<< metal1 >>
rect -2 64 26 72
rect 3 61 7 64
rect 3 56 7 57
rect 2 50 22 51
rect 2 46 13 50
rect 17 46 22 50
rect 2 45 22 46
rect 2 25 6 45
rect 13 43 17 45
rect 13 38 17 39
rect 10 34 22 35
rect 14 30 22 34
rect 10 29 22 30
rect 2 24 7 25
rect 2 20 3 24
rect 18 21 22 29
rect 2 19 7 20
rect 13 14 14 18
rect 18 14 19 18
rect 13 8 19 14
rect -2 4 4 8
rect 8 4 13 8
rect 17 4 26 8
rect -2 0 26 4
<< ntransistor >>
rect 9 19 11 25
<< ptransistor >>
rect 9 38 11 62
<< polycontact >>
rect 10 30 14 34
<< ndcontact >>
rect 3 20 7 24
rect 14 14 18 18
<< pdcontact >>
rect 3 57 7 61
rect 13 46 17 50
rect 13 39 17 43
<< psubstratepcontact >>
rect 4 4 8 8
rect 13 4 17 8
<< psubstratepdiff >>
rect 3 8 18 9
rect 3 4 4 8
rect 8 4 13 8
rect 17 4 18 8
rect 3 3 18 4
<< labels >>
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 4 12 4 6 vss
rlabel polycontact 12 32 12 32 6 a
rlabel metal1 12 48 12 48 6 z
rlabel metal1 12 68 12 68 6 vdd
rlabel metal1 20 28 20 28 6 a
rlabel metal1 20 48 20 48 6 z
<< end >>
