magic
tech scmos
timestamp 1179387686
<< checkpaint >>
rect -22 -22 94 94
<< ab >>
rect 0 0 72 72
<< pwell >>
rect -4 -4 76 32
<< nwell >>
rect -4 32 76 76
<< polysilicon >>
rect 6 68 30 70
rect 6 59 8 68
rect 18 60 20 64
rect 28 60 30 68
rect 38 68 60 70
rect 38 60 40 68
rect 48 60 50 64
rect 58 60 60 68
rect 2 58 8 59
rect 2 54 3 58
rect 7 54 8 58
rect 2 53 8 54
rect 18 35 20 38
rect 8 34 20 35
rect 8 30 9 34
rect 13 33 20 34
rect 28 33 30 38
rect 38 34 40 38
rect 48 34 50 38
rect 58 35 60 38
rect 58 34 64 35
rect 48 33 54 34
rect 13 30 14 33
rect 28 31 34 33
rect 8 29 14 30
rect 12 26 14 29
rect 22 25 24 29
rect 32 25 34 31
rect 48 30 49 33
rect 42 29 49 30
rect 53 29 54 33
rect 58 30 59 34
rect 63 30 64 34
rect 58 29 64 30
rect 42 28 54 29
rect 42 25 44 28
rect 61 25 63 29
rect 12 10 14 15
rect 22 6 24 14
rect 32 10 34 14
rect 42 10 44 14
rect 61 6 63 14
rect 22 4 63 6
<< ndiffusion >>
rect 2 20 12 26
rect 2 16 3 20
rect 7 16 12 20
rect 2 15 12 16
rect 14 25 19 26
rect 14 23 22 25
rect 14 19 16 23
rect 20 19 22 23
rect 14 15 22 19
rect 17 14 22 15
rect 24 24 32 25
rect 24 20 26 24
rect 30 20 32 24
rect 24 14 32 20
rect 34 24 42 25
rect 34 20 36 24
rect 40 20 42 24
rect 34 14 42 20
rect 44 19 61 25
rect 44 15 55 19
rect 59 15 61 19
rect 44 14 61 15
rect 63 24 70 25
rect 63 20 65 24
rect 69 20 70 24
rect 63 19 70 20
rect 63 14 68 19
<< pdiffusion >>
rect 11 59 18 60
rect 11 55 12 59
rect 16 55 18 59
rect 11 38 18 55
rect 20 43 28 60
rect 20 39 22 43
rect 26 39 28 43
rect 20 38 28 39
rect 30 43 38 60
rect 30 39 32 43
rect 36 39 38 43
rect 30 38 38 39
rect 40 43 48 60
rect 40 39 42 43
rect 46 39 48 43
rect 40 38 48 39
rect 50 59 58 60
rect 50 55 52 59
rect 56 55 58 59
rect 50 38 58 55
rect 60 52 65 60
rect 60 51 67 52
rect 60 47 62 51
rect 66 47 67 51
rect 60 46 67 47
rect 60 38 65 46
<< metal1 >>
rect -2 64 74 72
rect 11 59 17 64
rect 3 58 7 59
rect 11 55 12 59
rect 16 55 17 59
rect 51 59 57 64
rect 51 55 52 59
rect 56 55 57 59
rect 3 51 7 54
rect 3 47 62 51
rect 42 43 46 44
rect 2 35 6 43
rect 17 39 22 43
rect 26 39 27 43
rect 30 39 32 43
rect 36 39 38 43
rect 2 34 14 35
rect 2 30 9 34
rect 13 30 14 34
rect 2 29 14 30
rect 17 24 21 39
rect 30 37 38 39
rect 30 34 34 37
rect 42 34 46 39
rect 50 37 62 43
rect 58 35 62 37
rect 58 34 63 35
rect 16 23 21 24
rect 3 20 7 21
rect 20 19 21 23
rect 25 30 34 34
rect 38 30 46 34
rect 49 33 53 34
rect 25 24 31 30
rect 38 24 42 30
rect 58 30 59 34
rect 58 29 63 30
rect 49 27 53 29
rect 25 20 26 24
rect 30 20 31 24
rect 35 20 36 24
rect 40 20 42 24
rect 47 23 53 27
rect 66 25 70 51
rect 65 24 70 25
rect 16 18 21 19
rect 3 8 7 16
rect 17 17 21 18
rect 47 17 51 23
rect 69 20 70 24
rect 17 13 51 17
rect 55 19 59 20
rect 65 19 70 20
rect 55 8 59 15
rect -2 4 4 8
rect 8 4 74 8
rect -2 0 74 4
<< ntransistor >>
rect 12 15 14 26
rect 22 14 24 25
rect 32 14 34 25
rect 42 14 44 25
rect 61 14 63 25
<< ptransistor >>
rect 18 38 20 60
rect 28 38 30 60
rect 38 38 40 60
rect 48 38 50 60
rect 58 38 60 60
<< polycontact >>
rect 3 54 7 58
rect 9 30 13 34
rect 49 29 53 33
rect 59 30 63 34
<< ndcontact >>
rect 3 16 7 20
rect 16 19 20 23
rect 26 20 30 24
rect 36 20 40 24
rect 55 15 59 19
rect 65 20 69 24
<< pdcontact >>
rect 12 55 16 59
rect 22 39 26 43
rect 32 39 36 43
rect 42 39 46 43
rect 52 55 56 59
rect 62 47 66 51
<< psubstratepcontact >>
rect 4 4 8 8
<< psubstratepdiff >>
rect 3 8 9 9
rect 3 4 4 8
rect 8 4 9 8
rect 3 3 9 4
<< labels >>
rlabel polycontact 5 56 5 56 6 bn
rlabel polycontact 51 31 51 31 6 an
rlabel polycontact 12 32 12 32 6 a
rlabel metal1 4 36 4 36 6 a
rlabel metal1 5 53 5 53 6 bn
rlabel metal1 28 28 28 28 6 z
rlabel metal1 19 28 19 28 6 an
rlabel metal1 22 41 22 41 6 an
rlabel metal1 36 4 36 4 6 vss
rlabel ndcontact 38 22 38 22 6 ai
rlabel metal1 51 28 51 28 6 an
rlabel metal1 52 40 52 40 6 b
rlabel metal1 44 37 44 37 6 ai
rlabel metal1 36 40 36 40 6 z
rlabel metal1 36 68 36 68 6 vdd
rlabel metal1 60 36 60 36 6 b
rlabel metal1 68 35 68 35 6 bn
rlabel metal1 36 49 36 49 6 bn
<< end >>
