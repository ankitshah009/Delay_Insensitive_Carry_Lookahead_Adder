.subckt oa2a2a2a24_x4 i0 i1 i2 i3 i4 i5 i6 i7 q vdd vss
*   SPICE3 file   created from oa2a2a2a24_x4.ext -      technology: scmos
m00 w1     i7     w2     vdd p w=38u  l=2.3636u ad=190p     pd=48u      as=247p     ps=70u
m01 w2     i6     w1     vdd p w=38u  l=2.3636u ad=247p     pd=70u      as=190p     ps=48u
m02 w2     i5     w3     vdd p w=38u  l=2.3636u ad=247p     pd=70u      as=247p     ps=70u
m03 w3     i4     w2     vdd p w=38u  l=2.3636u ad=247p     pd=70u      as=247p     ps=70u
m04 w4     i3     w3     vdd p w=38u  l=2.3636u ad=190p     pd=48u      as=247p     ps=70u
m05 w3     i2     w4     vdd p w=38u  l=2.3636u ad=247p     pd=70u      as=190p     ps=48u
m06 w4     i1     vdd    vdd p w=38u  l=2.3636u ad=190p     pd=48u      as=247p     ps=70.0779u
m07 vdd    i0     w4     vdd p w=38u  l=2.3636u ad=247p     pd=70.0779u as=190p     ps=48u
m08 q      w1     vdd    vdd p w=39u  l=2.3636u ad=195p     pd=49u      as=253.5p   ps=71.9221u
m09 vdd    w1     q      vdd p w=39u  l=2.3636u ad=253.5p   pd=71.9221u as=195p     ps=49u
m10 w5     i7     vss    vss n w=19u  l=2.3636u ad=95p      pd=29u      as=133.336p ps=46.0708u
m11 w1     i6     w5     vss n w=19u  l=2.3636u ad=123.12p  pd=41.5467u as=95p      ps=29u
m12 w6     i5     vss    vss n w=19u  l=2.3636u ad=57p      pd=25u      as=133.336p ps=46.0708u
m13 w1     i4     w6     vss n w=19u  l=2.3636u ad=123.12p  pd=41.5467u as=57p      ps=25u
m14 w7     i3     w1     vss n w=19u  l=2.3636u ad=57p      pd=25u      as=123.12p  ps=41.5467u
m15 vss    i2     w7     vss n w=19u  l=2.3636u ad=133.336p pd=46.0708u as=57p      ps=25u
m16 w8     i1     w1     vss n w=18u  l=2.3636u ad=54p      pd=24u      as=116.64p  ps=39.36u
m17 vss    i0     w8     vss n w=18u  l=2.3636u ad=126.319p pd=43.646u  as=54p      ps=24u
m18 q      w1     vss    vss n w=19u  l=2.3636u ad=95p      pd=29u      as=133.336p ps=46.0708u
m19 vss    w1     q      vss n w=19u  l=2.3636u ad=133.336p pd=46.0708u as=95p      ps=29u
C0  vss    i3     0.013f
C1  w3     w1     0.004f
C2  w4     i0     0.019f
C3  vdd    i1     0.020f
C4  i3     i4     0.261f
C5  i2     i5     0.066f
C6  vss    q      0.082f
C7  w4     i2     0.045f
C8  vss    i5     0.013f
C9  vdd    i3     0.010f
C10 i3     i6     0.033f
C11 i4     i5     0.290f
C12 w7     w1     0.012f
C13 q      vdd    0.163f
C14 w1     i1     0.150f
C15 vdd    i5     0.010f
C16 w3     i3     0.023f
C17 vss    i7     0.040f
C18 i5     i6     0.097f
C19 w5     w1     0.016f
C20 vdd    w4     0.232f
C21 w2     i4     0.006f
C22 i0     i2     0.016f
C23 w3     i5     0.013f
C24 w1     i3     0.057f
C25 vdd    i7     0.010f
C26 w8     vss    0.011f
C27 i6     i7     0.133f
C28 vss    i0     0.027f
C29 q      w1     0.026f
C30 w4     w3     0.149f
C31 vdd    w2     0.246f
C32 w1     i5     0.086f
C33 i1     i3     0.041f
C34 w2     i6     0.051f
C35 w6     vss    0.011f
C36 w4     w1     0.005f
C37 w3     w2     0.167f
C38 vdd    i0     0.085f
C39 q      i1     0.043f
C40 vss    i2     0.013f
C41 i2     i4     0.105f
C42 w1     i7     0.228f
C43 w2     w1     0.101f
C44 vss    i4     0.013f
C45 w4     i1     0.034f
C46 vdd    i2     0.010f
C47 i3     i5     0.105f
C48 vss    i6     0.013f
C49 w1     i0     0.130f
C50 vdd    i4     0.010f
C51 w3     i2     0.013f
C52 i4     i6     0.062f
C53 q      w4     0.025f
C54 w6     w1     0.012f
C55 vdd    i6     0.010f
C56 w3     i4     0.019f
C57 i0     i1     0.142f
C58 w1     i2     0.078f
C59 i5     i7     0.048f
C60 vss    w1     0.578f
C61 vdd    w3     0.338f
C62 i1     i2     0.057f
C63 w1     i4     0.078f
C64 w2     i5     0.039f
C65 w7     vss    0.011f
C66 q      i0     0.233f
C67 w4     w2     0.007f
C68 vdd    w1     0.042f
C69 vss    i1     0.022f
C70 w2     i7     0.023f
C71 i2     i3     0.290f
C72 w1     i6     0.212f
C73 w5     vss    0.019f
C75 q      vss    0.014f
C77 w4     vss    0.005f
C78 w2     vss    0.003f
C79 w1     vss    0.095f
C80 i0     vss    0.032f
C81 i1     vss    0.030f
C82 i2     vss    0.029f
C83 i3     vss    0.030f
C84 i4     vss    0.027f
C85 i5     vss    0.030f
C86 i6     vss    0.038f
C87 i7     vss    0.031f
.ends
