magic
tech scmos
timestamp 1180600611
<< checkpaint >>
rect -22 -22 92 122
<< ab >>
rect 0 0 70 100
<< pwell >>
rect -4 -4 74 48
<< nwell >>
rect -4 48 74 104
<< polysilicon >>
rect 45 94 47 98
rect 57 94 59 98
rect 11 81 13 85
rect 23 81 25 85
rect 35 82 37 86
rect 11 33 13 61
rect 23 53 25 61
rect 35 59 37 62
rect 17 52 25 53
rect 17 48 18 52
rect 22 48 25 52
rect 17 47 25 48
rect 31 57 37 59
rect 7 32 13 33
rect 7 28 8 32
rect 12 28 13 32
rect 7 27 13 28
rect 11 24 13 27
rect 19 24 21 47
rect 31 43 33 57
rect 45 43 47 55
rect 57 43 59 55
rect 27 42 33 43
rect 27 38 28 42
rect 32 38 33 42
rect 27 37 33 38
rect 37 42 59 43
rect 37 38 38 42
rect 42 38 59 42
rect 37 37 59 38
rect 27 24 29 37
rect 45 25 47 37
rect 57 25 59 37
rect 11 2 13 6
rect 19 2 21 6
rect 27 2 29 6
rect 45 2 47 6
rect 57 2 59 6
<< ndiffusion >>
rect 35 24 45 25
rect 3 22 11 24
rect 3 18 4 22
rect 8 18 11 22
rect 3 6 11 18
rect 13 6 19 24
rect 21 6 27 24
rect 29 12 45 24
rect 29 8 38 12
rect 42 8 45 12
rect 29 6 45 8
rect 47 22 57 25
rect 47 18 50 22
rect 54 18 57 22
rect 47 6 57 18
rect 59 22 67 25
rect 59 18 62 22
rect 66 18 67 22
rect 59 12 67 18
rect 59 8 62 12
rect 66 8 67 12
rect 59 6 67 8
<< pdiffusion >>
rect 37 94 43 95
rect 15 92 21 93
rect 15 88 16 92
rect 20 88 21 92
rect 37 90 38 94
rect 42 90 45 94
rect 37 89 45 90
rect 3 82 9 83
rect 3 78 4 82
rect 8 81 9 82
rect 15 81 21 88
rect 27 82 33 83
rect 39 82 45 89
rect 27 81 28 82
rect 8 78 11 81
rect 3 61 11 78
rect 13 61 23 81
rect 25 78 28 81
rect 32 78 35 82
rect 25 62 35 78
rect 37 62 45 82
rect 25 61 30 62
rect 39 55 45 62
rect 47 82 57 94
rect 47 78 50 82
rect 54 78 57 82
rect 47 72 57 78
rect 47 68 50 72
rect 54 68 57 72
rect 47 62 57 68
rect 47 58 50 62
rect 54 58 57 62
rect 47 55 57 58
rect 59 92 67 94
rect 59 88 62 92
rect 66 88 67 92
rect 59 82 67 88
rect 59 78 62 82
rect 66 78 67 82
rect 59 72 67 78
rect 59 68 62 72
rect 66 68 67 72
rect 59 62 67 68
rect 59 58 62 62
rect 66 58 67 62
rect 59 55 67 58
<< metal1 >>
rect -2 94 72 100
rect -2 92 38 94
rect -2 88 16 92
rect 20 90 38 92
rect 42 92 72 94
rect 42 90 62 92
rect 20 88 62 90
rect 66 88 72 92
rect 48 82 52 83
rect 62 82 66 88
rect 3 78 4 82
rect 8 78 28 82
rect 32 78 42 82
rect 8 32 12 73
rect 8 27 12 28
rect 18 52 22 73
rect 18 27 22 48
rect 28 42 32 73
rect 28 27 32 38
rect 38 42 42 78
rect 38 22 42 38
rect 3 18 4 22
rect 8 18 42 22
rect 48 78 50 82
rect 54 78 55 82
rect 48 72 52 78
rect 62 72 66 78
rect 48 68 50 72
rect 54 68 55 72
rect 48 62 52 68
rect 62 62 66 68
rect 48 58 50 62
rect 54 58 55 62
rect 48 22 52 58
rect 62 57 66 58
rect 62 22 66 23
rect 48 18 50 22
rect 54 18 55 22
rect 48 17 52 18
rect 62 12 66 18
rect -2 8 38 12
rect 42 8 62 12
rect 66 8 72 12
rect -2 0 72 8
<< ntransistor >>
rect 11 6 13 24
rect 19 6 21 24
rect 27 6 29 24
rect 45 6 47 25
rect 57 6 59 25
<< ptransistor >>
rect 11 61 13 81
rect 23 61 25 81
rect 35 62 37 82
rect 45 55 47 94
rect 57 55 59 94
<< polycontact >>
rect 18 48 22 52
rect 8 28 12 32
rect 28 38 32 42
rect 38 38 42 42
<< ndcontact >>
rect 4 18 8 22
rect 38 8 42 12
rect 50 18 54 22
rect 62 18 66 22
rect 62 8 66 12
<< pdcontact >>
rect 16 88 20 92
rect 38 90 42 94
rect 4 78 8 82
rect 28 78 32 82
rect 50 78 54 82
rect 50 68 54 72
rect 50 58 54 62
rect 62 88 66 92
rect 62 78 66 82
rect 62 68 66 72
rect 62 58 66 62
<< labels >>
rlabel metal1 10 50 10 50 6 i0
rlabel metal1 30 50 30 50 6 i2
rlabel polycontact 20 50 20 50 6 i1
rlabel metal1 35 6 35 6 6 vss
rlabel metal1 50 50 50 50 6 q
rlabel metal1 35 94 35 94 6 vdd
<< end >>
