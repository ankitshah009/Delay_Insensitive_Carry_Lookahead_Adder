magic
tech scmos
timestamp 1179385563
<< checkpaint >>
rect -22 -25 54 105
<< ab >>
rect 0 0 32 80
<< pwell >>
rect -4 -7 36 36
<< nwell >>
rect -4 36 36 87
<< polysilicon >>
rect 9 60 11 65
rect 21 61 27 62
rect 21 57 22 61
rect 26 57 27 61
rect 21 56 27 57
rect 21 48 23 56
rect 9 39 11 42
rect 9 38 16 39
rect 9 34 11 38
rect 15 34 16 38
rect 9 33 16 34
rect 9 30 11 33
rect 21 30 23 42
rect 9 16 11 21
rect 21 19 23 24
<< ndiffusion >>
rect 2 29 9 30
rect 2 25 3 29
rect 7 25 9 29
rect 2 24 9 25
rect 4 21 9 24
rect 11 29 21 30
rect 11 25 14 29
rect 18 25 21 29
rect 11 24 21 25
rect 23 29 30 30
rect 23 25 25 29
rect 29 25 30 29
rect 23 24 30 25
rect 11 21 19 24
<< pdiffusion >>
rect 13 72 19 73
rect 13 68 14 72
rect 18 68 19 72
rect 13 60 19 68
rect 4 55 9 60
rect 2 54 9 55
rect 2 50 3 54
rect 7 50 9 54
rect 2 47 9 50
rect 2 43 3 47
rect 7 43 9 47
rect 2 42 9 43
rect 11 48 19 60
rect 11 42 21 48
rect 23 47 30 48
rect 23 43 25 47
rect 29 43 30 47
rect 23 42 30 43
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect -2 72 34 78
rect -2 68 14 72
rect 18 68 34 72
rect 18 61 30 63
rect 2 54 14 55
rect 2 50 3 54
rect 7 50 14 54
rect 2 49 14 50
rect 18 49 22 61
rect 26 57 30 61
rect 2 47 7 49
rect 2 43 3 47
rect 2 42 7 43
rect 25 47 29 48
rect 2 29 6 42
rect 25 38 29 43
rect 10 34 11 38
rect 15 34 30 38
rect 14 29 18 30
rect 2 25 3 29
rect 7 25 8 29
rect 24 29 30 34
rect 24 25 25 29
rect 29 25 30 29
rect 14 12 18 25
rect -2 2 34 12
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
<< ntransistor >>
rect 9 21 11 30
rect 21 24 23 30
<< ptransistor >>
rect 9 42 11 60
rect 21 42 23 48
<< polycontact >>
rect 22 57 26 61
rect 11 34 15 38
<< ndcontact >>
rect 3 25 7 29
rect 14 25 18 29
rect 25 25 29 29
<< pdcontact >>
rect 14 68 18 72
rect 3 50 7 54
rect 3 43 7 47
rect 25 43 29 47
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
<< psubstratepdiff >>
rect 0 2 32 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 32 2
rect 0 -3 32 -2
<< nsubstratendiff >>
rect 0 82 32 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 32 82
rect 0 77 32 78
<< labels >>
rlabel polycontact 12 36 12 36 6 an
rlabel metal1 4 40 4 40 6 z
rlabel metal1 12 52 12 52 6 z
rlabel metal1 16 6 16 6 6 vss
rlabel metal1 20 56 20 56 6 a
rlabel metal1 16 74 16 74 6 vdd
rlabel metal1 20 36 20 36 6 an
rlabel metal1 27 36 27 36 6 an
rlabel metal1 28 60 28 60 6 a
<< end >>
