.subckt nxr2_x4 i0 i1 nq vdd vss
*   SPICE3 file   created from nxr2_x4.ext -      technology: scmos
m00 vdd    i0     w1     vdd p w=20u  l=2.3636u ad=131.546p pd=39.1753u as=160p     ps=56u
m01 w2     i0     vdd    vdd p w=38u  l=2.3636u ad=190p     pd=48.183u  as=249.938p ps=74.433u
m02 w3     w4     w2     vdd p w=38u  l=2.3636u ad=190p     pd=48.3636u as=190p     ps=48.183u
m03 w2     w1     w3     vdd p w=39u  l=2.3636u ad=195p     pd=49.451u  as=195p     ps=49.6364u
m04 vdd    i1     w2     vdd p w=38u  l=2.3636u ad=249.938p pd=74.433u  as=190p     ps=48.183u
m05 w4     i1     vdd    vdd p w=20u  l=2.3636u ad=176p     pd=62u      as=131.546p ps=39.1753u
m06 nq     w3     vdd    vdd p w=39u  l=2.3636u ad=195p     pd=49u      as=256.515p ps=76.3918u
m07 vdd    w3     nq     vdd p w=39u  l=2.3636u ad=256.515p pd=76.3918u as=195p     ps=49u
m08 vss    i0     w1     vss n w=10u  l=2.3636u ad=65.7895p pd=23.3684u as=80p      ps=36u
m09 w5     i0     vss    vss n w=18u  l=2.3636u ad=90p      pd=28u      as=118.421p ps=42.0632u
m10 w3     i1     w5     vss n w=18u  l=2.3636u ad=90p      pd=28.2162u as=90p      ps=28u
m11 w6     w1     w3     vss n w=19u  l=2.3636u ad=95p      pd=29u      as=95p      ps=29.7838u
m12 vss    w4     w6     vss n w=19u  l=2.3636u ad=125p     pd=44.4u    as=95p      ps=29u
m13 w4     i1     vss    vss n w=10u  l=2.3636u ad=146p     pd=58u      as=65.7895p ps=23.3684u
m14 nq     w3     vss    vss n w=19u  l=2.3636u ad=95p      pd=29u      as=125p     ps=44.4u
m15 vss    w3     nq     vss n w=19u  l=2.3636u ad=125p     pd=44.4u    as=95p      ps=29u
C0  w1     vdd    0.011f
C1  w4     i0     0.047f
C2  nq     w2     0.003f
C3  vss    i1     0.074f
C4  i0     vdd    0.084f
C5  vss    w4     0.040f
C6  w3     i1     0.312f
C7  w2     w1     0.005f
C8  w3     w4     0.272f
C9  vss    vdd    0.004f
C10 w5     vss    0.019f
C11 w3     vdd    0.069f
C12 w2     i0     0.024f
C13 i1     w4     0.424f
C14 vss    nq     0.082f
C15 w5     w3     0.018f
C16 i1     vdd    0.109f
C17 w1     i0     0.227f
C18 nq     w3     0.143f
C19 w4     vdd    0.027f
C20 w3     w2     0.142f
C21 nq     i1     0.065f
C22 vss    w1     0.029f
C23 w3     w1     0.082f
C24 w2     i1     0.011f
C25 nq     w4     0.068f
C26 vss    i0     0.047f
C27 w6     vss    0.019f
C28 i1     w1     0.091f
C29 w3     i0     0.273f
C30 nq     vdd    0.243f
C31 w2     w4     0.027f
C32 w6     w3     0.019f
C33 i1     i0     0.035f
C34 w2     vdd    0.193f
C35 w1     w4     0.126f
C36 vss    w3     0.391f
C38 nq     vss    0.012f
C39 w3     vss    0.079f
C40 i1     vss    0.057f
C41 w1     vss    0.052f
C42 w4     vss    0.056f
C43 i0     vss    0.042f
.ends
