.subckt iv1v4x8 a vdd vss z
*   SPICE3 file   created from iv1v4x8.ext -      technology: scmos
m00 z      a      vdd    vdd p w=28u  l=2.3636u ad=121.188p pd=41.5625u as=135.625p ps=46.8125u
m01 vdd    a      z      vdd p w=28u  l=2.3636u ad=135.625p pd=46.8125u as=121.188p ps=41.5625u
m02 z      a      vdd    vdd p w=28u  l=2.3636u ad=121.188p pd=41.5625u as=135.625p ps=46.8125u
m03 vdd    a      z      vdd p w=28u  l=2.3636u ad=135.625p pd=46.8125u as=121.188p ps=41.5625u
m04 z      a      vdd    vdd p w=16u  l=2.3636u ad=69.25p   pd=23.75u   as=77.5p    ps=26.75u
m05 z      a      vss    vss n w=16u  l=2.3636u ad=64p      pd=24u      as=128p     ps=48u
m06 vss    a      z      vss n w=16u  l=2.3636u ad=128p     pd=48u      as=64p      ps=24u
C0  vss    vdd    0.009f
C1  z      a      0.235f
C2  vss    z      0.193f
C3  vss    a      0.061f
C4  z      vdd    0.188f
C5  vdd    a      0.040f
C7  z      vss    0.005f
C9  a      vss    0.067f
.ends
