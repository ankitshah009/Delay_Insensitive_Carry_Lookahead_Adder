.subckt inv_x2 i nq vdd vss
*   SPICE3 file   created from inv_x2.ext -      technology: scmos
m00 nq     i      vdd    vdd p w=30u  l=2.3636u ad=240p     pd=76u      as=364p     ps=96u
m01 nq     i      vss    vss n w=20u  l=2.3636u ad=160p     pd=56u      as=256p     ps=74u
C0  nq     i      0.334f
C1  i      vdd    0.083f
C2  vss    i      0.062f
C3  nq     vdd    0.024f
C4  vss    nq     0.024f
C6  nq     vss    0.010f
C7  i      vss    0.027f
.ends
