.subckt mxi2v2x05 a0 a1 s vdd vss z
*   SPICE3 file   created from mxi2v2x05.ext -      technology: scmos
m00 sn     s      vdd    vdd p w=6u   l=2.3636u ad=42p      pd=26u      as=70.4p    ps=27.6u
m01 a0n    a0     vdd    vdd p w=12u  l=2.3636u ad=48p      pd=20u      as=140.8p   ps=55.2u
m02 z      s      a0n    vdd p w=12u  l=2.3636u ad=48p      pd=20u      as=48p      ps=20u
m03 a1n    sn     z      vdd p w=12u  l=2.3636u ad=48p      pd=20u      as=48p      ps=20u
m04 vdd    a1     a1n    vdd p w=12u  l=2.3636u ad=140.8p   pd=55.2u    as=48p      ps=20u
m05 a0n    a0     vss    vss n w=6u   l=2.3636u ad=24p      pd=14u      as=44.6667p ps=23.3333u
m06 z      sn     a0n    vss n w=6u   l=2.3636u ad=24p      pd=14u      as=24p      ps=14u
m07 a1n    s      z      vss n w=6u   l=2.3636u ad=24p      pd=14u      as=24p      ps=14u
m08 vss    a1     a1n    vss n w=6u   l=2.3636u ad=44.6667p pd=23.3333u as=24p      ps=14u
m09 sn     s      vss    vss n w=6u   l=2.3636u ad=42p      pd=26u      as=44.6667p ps=23.3333u
C0  z      vdd    0.012f
C1  a1     a0     0.022f
C2  a0n    s      0.017f
C3  vss    a1n    0.068f
C4  sn     s      0.332f
C5  a1     vdd    0.012f
C6  a1n    z      0.293f
C7  vss    a0n    0.067f
C8  a0     vdd    0.075f
C9  z      a0n    0.172f
C10 vss    sn     0.028f
C11 a1n    a1     0.094f
C12 z      sn     0.065f
C13 a1n    a0     0.016f
C14 a0n    a1     0.020f
C15 vss    s      0.027f
C16 a1n    vdd    0.009f
C17 a1     sn     0.137f
C18 a0n    a0     0.078f
C19 z      s      0.038f
C20 a1     s      0.137f
C21 sn     a0     0.048f
C22 a0n    vdd    0.010f
C23 vss    z      0.061f
C24 a0     s      0.042f
C25 sn     vdd    0.216f
C26 a1n    a0n    0.068f
C27 vss    a1     0.085f
C28 s      vdd    0.064f
C29 a1n    sn     0.057f
C30 vss    a0     0.023f
C31 z      a1     0.037f
C32 a0n    sn     0.038f
C33 vss    vdd    0.007f
C34 z      a0     0.038f
C35 a1n    s      0.018f
C37 a1n    vss    0.009f
C38 z      vss    0.009f
C39 a0n    vss    0.009f
C40 a1     vss    0.024f
C41 sn     vss    0.041f
C42 a0     vss    0.024f
C43 s      vss    0.070f
.ends
