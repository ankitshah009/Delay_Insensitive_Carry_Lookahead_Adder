magic
tech scmos
timestamp 1170759844
<< checkpaint >>
rect -22 -26 54 114
<< ab >>
rect 0 0 32 88
<< pwell >>
rect -4 -8 36 40
<< nwell >>
rect -4 40 36 96
<< polysilicon >>
rect 2 77 11 83
rect 9 74 11 77
rect 21 77 30 83
rect 21 74 23 77
rect 9 43 11 46
rect 21 43 23 46
rect 2 37 14 43
rect 18 37 30 43
rect 9 34 11 37
rect 21 34 23 37
rect 9 11 11 14
rect 2 5 11 11
rect 21 11 23 14
rect 21 5 30 11
<< ndiffusion >>
rect 2 26 9 34
rect 2 22 3 26
rect 7 22 9 26
rect 2 19 9 22
rect 2 15 3 19
rect 7 15 9 19
rect 2 14 9 15
rect 11 30 21 34
rect 11 26 14 30
rect 18 26 21 30
rect 11 22 21 26
rect 11 18 14 22
rect 18 18 21 22
rect 11 14 21 18
rect 23 26 30 34
rect 23 22 25 26
rect 29 22 30 26
rect 23 19 30 22
rect 23 15 25 19
rect 29 15 30 19
rect 23 14 30 15
rect 13 2 19 14
<< pdiffusion >>
rect 13 74 19 86
rect 2 46 9 74
rect 11 70 21 74
rect 11 66 14 70
rect 18 66 21 70
rect 11 62 21 66
rect 11 58 14 62
rect 18 58 21 62
rect 11 54 21 58
rect 11 50 14 54
rect 18 50 21 54
rect 11 46 21 50
rect 23 46 30 74
<< metal1 >>
rect -2 86 2 90
rect 10 86 22 90
rect 30 86 34 90
rect 5 78 6 82
rect 10 78 22 82
rect 26 78 27 82
rect 14 70 18 71
rect 14 62 18 66
rect 14 54 18 58
rect 14 30 18 50
rect 3 26 7 27
rect 3 19 7 22
rect 14 22 18 26
rect 14 17 18 18
rect 25 26 29 27
rect 25 19 29 22
rect 3 10 7 15
rect 3 2 7 6
rect 25 10 29 15
rect 25 2 29 6
rect -2 -2 2 2
rect 10 -2 22 2
rect 30 -2 34 2
<< metal2 >>
rect -2 86 6 90
rect 10 86 22 90
rect 26 86 34 90
rect -2 82 34 86
rect -2 78 6 82
rect 10 78 22 82
rect 26 78 34 82
rect -2 76 34 78
rect -2 10 34 12
rect -2 6 3 10
rect 7 6 25 10
rect 29 6 34 10
rect -2 2 34 6
rect -2 -2 6 2
rect 10 -2 22 2
rect 26 -2 34 2
<< ntransistor >>
rect 9 14 11 34
rect 21 14 23 34
<< ptransistor >>
rect 9 46 11 74
rect 21 46 23 74
<< ndcontact >>
rect 3 22 7 26
rect 3 15 7 19
rect 14 26 18 30
rect 14 18 18 22
rect 25 22 29 26
rect 25 15 29 19
<< pdcontact >>
rect 14 66 18 70
rect 14 58 18 62
rect 14 50 18 54
<< m2contact >>
rect 6 86 10 90
rect 22 86 26 90
rect 6 78 10 82
rect 22 78 26 82
rect 3 6 7 10
rect 25 6 29 10
rect 6 -2 10 2
rect 22 -2 26 2
<< psubstratepcontact >>
rect 2 -2 6 2
rect 26 -2 30 2
<< nsubstratencontact >>
rect 2 86 6 90
rect 26 86 30 90
<< psubstratepdiff >>
rect 0 2 7 3
rect 25 2 32 3
rect 0 -2 2 2
rect 6 -2 7 2
rect 0 -3 7 -2
rect 25 -2 26 2
rect 30 -2 32 2
rect 25 -3 32 -2
<< nsubstratendiff >>
rect 0 90 7 91
rect 0 86 2 90
rect 6 86 7 90
rect 25 90 32 91
rect 25 86 26 90
rect 30 86 32 90
rect 0 85 7 86
rect 25 85 32 86
<< labels >>
rlabel metal1 16 44 16 44 6 z
rlabel metal2 16 6 16 6 6 vss
rlabel metal2 16 82 16 82 6 vdd
<< end >>
