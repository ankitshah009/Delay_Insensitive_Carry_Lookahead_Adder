.subckt mxi2_x05 a0 a1 s vdd vss z
*   SPICE3 file   created from mxi2_x05.ext -      technology: scmos
m00 w1     s      vdd    vdd p w=20u  l=2.3636u ad=60p      pd=26u      as=179.655p ps=51.7241u
m01 z      a0     w1     vdd p w=20u  l=2.3636u ad=100p     pd=30u      as=60p      ps=26u
m02 w2     a1     z      vdd p w=20u  l=2.3636u ad=60p      pd=26u      as=100p     ps=30u
m03 vdd    sn     w2     vdd p w=20u  l=2.3636u ad=179.655p pd=51.7241u as=60p      ps=26u
m04 sn     s      vdd    vdd p w=18u  l=2.3636u ad=132p     pd=52u      as=161.69p  ps=46.5517u
m05 w3     a1     vss    vss n w=9u   l=2.3636u ad=27p      pd=15u      as=94p      ps=35.3333u
m06 z      s      w3     vss n w=9u   l=2.3636u ad=45p      pd=19u      as=27p      ps=15u
m07 w4     a0     z      vss n w=9u   l=2.3636u ad=27p      pd=15u      as=45p      ps=19u
m08 vss    sn     w4     vss n w=9u   l=2.3636u ad=94p      pd=35.3333u as=27p      ps=15u
m09 sn     s      vss    vss n w=9u   l=2.3636u ad=63p      pd=34u      as=94p      ps=35.3333u
C0  a1     vdd    0.021f
C1  a0     s      0.169f
C2  vss    sn     0.058f
C3  s      vdd    0.216f
C4  z      sn     0.098f
C5  vss    a0     0.093f
C6  w1     a1     0.016f
C7  z      a0     0.177f
C8  w2     s      0.012f
C9  z      vdd    0.017f
C10 sn     a0     0.087f
C11 w1     s      0.012f
C12 a1     s      0.368f
C13 sn     vdd    0.010f
C14 w2     z      0.015f
C15 vss    a1     0.034f
C16 w3     a0     0.004f
C17 z      a1     0.167f
C18 vss    s      0.020f
C19 z      s      0.226f
C20 sn     a1     0.073f
C21 w4     z      0.012f
C22 sn     s      0.234f
C23 a1     a0     0.276f
C24 vss    z      0.157f
C26 z      vss    0.013f
C27 sn     vss    0.046f
C28 a1     vss    0.042f
C29 a0     vss    0.037f
C30 s      vss    0.061f
.ends
