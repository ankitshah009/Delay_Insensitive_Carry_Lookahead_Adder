.subckt bsi2v2x1 a0 a1 s vdd vss z0 z1
*   SPICE3 file   created from bsi2v2x1.ext -      technology: scmos
m00 a0n    a0     vdd    vdd p w=21u  l=2.3636u ad=99.8308p pd=38.1231u as=202.246p ps=48.4615u
m01 z0     s      a0n    vdd p w=22u  l=2.3636u ad=88p      pd=30u      as=104.585p ps=39.9385u
m02 a1n    sn     z0     vdd p w=22u  l=2.3636u ad=104p     pd=39.3333u as=88p      ps=30u
m03 vdd    s      sn     vdd p w=22u  l=2.3636u ad=211.877p pd=50.7692u as=122p     ps=58u
m04 a1n    a1     vdd    vdd p w=22u  l=2.3636u ad=104p     pd=39.3333u as=211.877p ps=50.7692u
m05 z1     s      a1n    vdd p w=22u  l=2.3636u ad=88p      pd=30u      as=104p     ps=39.3333u
m06 a0n    sn     z1     vdd p w=22u  l=2.3636u ad=104.585p pd=39.9385u as=88p      ps=30u
m07 a0n    a0     vss    vss n w=10u  l=2.3636u ad=47.3333p pd=23.3333u as=98.6667p ps=34u
m08 z0     sn     a0n    vss n w=10u  l=2.3636u ad=40p      pd=18u      as=47.3333p ps=23.3333u
m09 a1n    s      z0     vss n w=10u  l=2.3636u ad=48p      pd=23.3333u as=40p      ps=18u
m10 vss    s      sn     vss n w=10u  l=2.3636u ad=98.6667p pd=34u      as=62p      ps=34u
m11 a1n    a1     vss    vss n w=10u  l=2.3636u ad=48p      pd=23.3333u as=98.6667p ps=34u
m12 z1     sn     a1n    vss n w=10u  l=2.3636u ad=40p      pd=18u      as=48p      ps=23.3333u
m13 a0n    s      z1     vss n w=10u  l=2.3636u ad=47.3333p pd=23.3333u as=40p      ps=18u
C0  z0     sn     0.051f
C1  a1n    a0     0.022f
C2  a1     s      0.151f
C3  z1     vdd    0.019f
C4  vss    z1     0.070f
C5  a1n    vdd    0.047f
C6  z0     s      0.045f
C7  a0n    a0     0.095f
C8  z1     a1     0.053f
C9  vss    a1n    0.373f
C10 a0n    vdd    0.647f
C11 sn     s      0.378f
C12 vss    a0n    0.050f
C13 a1     a1n    0.295f
C14 a0     vdd    0.068f
C15 vss    a0     0.042f
C16 a1n    z0     0.221f
C17 a1     a0n    0.156f
C18 z1     sn     0.030f
C19 a1n    sn     0.332f
C20 z0     a0n    0.361f
C21 z1     s      0.037f
C22 vss    vdd    0.003f
C23 a0n    sn     0.087f
C24 a1n    s      0.160f
C25 a1     vdd    0.066f
C26 z0     a0     0.041f
C27 vss    a1     0.017f
C28 a0n    s      0.101f
C29 z0     vdd    0.035f
C30 sn     a0     0.055f
C31 vss    z0     0.058f
C32 z1     a1n    0.178f
C33 sn     vdd    0.022f
C34 a0     s      0.043f
C35 a1     z0     0.010f
C36 z1     a0n    0.299f
C37 vss    sn     0.050f
C38 s      vdd    0.053f
C39 vss    s      0.021f
C40 a1n    a0n    0.259f
C41 a1     sn     0.095f
C43 z1     vss    0.011f
C44 a1     vss    0.019f
C45 a1n    vss    0.023f
C46 z0     vss    0.008f
C47 a0n    vss    0.023f
C48 sn     vss    0.088f
C49 a0     vss    0.037f
C50 s      vss    0.105f
.ends
