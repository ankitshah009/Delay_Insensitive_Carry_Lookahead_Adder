magic
tech scmos
timestamp 1179387067
<< checkpaint >>
rect -22 -25 214 105
<< ab >>
rect 0 0 192 80
<< pwell >>
rect -4 -7 196 36
<< nwell >>
rect -4 36 196 87
<< polysilicon >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 39 70 41 74
rect 49 70 51 74
rect 56 70 58 74
rect 66 70 68 74
rect 73 70 75 74
rect 83 70 85 74
rect 90 70 92 74
rect 100 70 102 74
rect 107 70 109 74
rect 117 70 119 74
rect 124 70 126 74
rect 134 70 136 74
rect 141 70 143 74
rect 151 70 153 74
rect 158 70 160 74
rect 168 63 170 68
rect 175 63 177 68
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 39 39 41 42
rect 49 39 51 42
rect 9 38 41 39
rect 9 34 26 38
rect 30 37 41 38
rect 30 34 31 37
rect 9 33 31 34
rect 9 30 11 33
rect 19 30 21 33
rect 29 30 31 33
rect 39 30 41 37
rect 45 38 51 39
rect 45 34 46 38
rect 50 34 51 38
rect 56 39 58 42
rect 66 39 68 42
rect 56 37 68 39
rect 73 39 75 42
rect 83 39 85 42
rect 73 38 85 39
rect 73 37 77 38
rect 45 33 51 34
rect 59 29 61 37
rect 76 34 77 37
rect 81 37 85 38
rect 90 39 92 42
rect 100 39 102 42
rect 90 38 102 39
rect 81 34 82 37
rect 76 33 82 34
rect 70 29 72 33
rect 80 29 82 33
rect 90 34 91 38
rect 95 37 102 38
rect 107 39 109 42
rect 117 39 119 42
rect 124 39 126 42
rect 134 39 136 42
rect 107 38 119 39
rect 95 34 96 37
rect 90 33 96 34
rect 107 34 111 38
rect 115 37 119 38
rect 123 37 136 39
rect 141 39 143 42
rect 151 39 153 42
rect 141 38 153 39
rect 115 34 116 37
rect 107 33 116 34
rect 123 36 129 37
rect 123 33 124 36
rect 49 25 51 29
rect 90 28 92 33
rect 100 31 116 33
rect 122 32 124 33
rect 128 32 129 36
rect 141 34 142 38
rect 146 37 153 38
rect 158 39 160 42
rect 168 39 170 42
rect 158 38 170 39
rect 146 34 147 37
rect 141 33 147 34
rect 158 34 161 38
rect 165 37 170 38
rect 175 39 177 42
rect 175 38 183 39
rect 165 34 168 37
rect 158 33 168 34
rect 175 34 178 38
rect 182 34 183 38
rect 175 33 183 34
rect 122 31 129 32
rect 134 31 147 33
rect 156 31 168 33
rect 100 28 102 31
rect 112 28 114 31
rect 122 28 124 31
rect 134 28 136 31
rect 144 28 146 31
rect 156 28 158 31
rect 166 28 168 31
rect 177 30 179 33
rect 80 12 82 16
rect 9 6 11 10
rect 19 6 21 10
rect 29 6 31 10
rect 39 8 41 11
rect 49 8 51 11
rect 39 6 51 8
rect 59 8 61 11
rect 70 8 72 11
rect 90 8 92 16
rect 59 6 92 8
rect 100 6 102 10
rect 112 6 114 10
rect 122 6 124 10
rect 177 15 179 19
rect 134 6 136 10
rect 144 6 146 10
rect 156 8 158 13
rect 166 8 168 13
<< ndiffusion >>
rect 2 29 9 30
rect 2 25 3 29
rect 7 25 9 29
rect 2 22 9 25
rect 2 18 3 22
rect 7 18 9 22
rect 2 17 9 18
rect 4 10 9 17
rect 11 29 19 30
rect 11 25 13 29
rect 17 25 19 29
rect 11 10 19 25
rect 21 21 29 30
rect 21 17 23 21
rect 27 17 29 21
rect 21 10 29 17
rect 31 29 39 30
rect 31 25 33 29
rect 37 25 39 29
rect 31 11 39 25
rect 41 25 46 30
rect 54 25 59 29
rect 41 21 49 25
rect 41 17 43 21
rect 47 17 49 21
rect 41 11 49 17
rect 51 24 59 25
rect 51 20 53 24
rect 57 20 59 24
rect 51 11 59 20
rect 61 16 70 29
rect 61 12 64 16
rect 68 12 70 16
rect 61 11 70 12
rect 72 26 80 29
rect 72 22 74 26
rect 78 22 80 26
rect 72 16 80 22
rect 82 28 87 29
rect 170 28 177 30
rect 82 21 90 28
rect 82 17 84 21
rect 88 17 90 21
rect 82 16 90 17
rect 92 26 100 28
rect 92 22 94 26
rect 98 22 100 26
rect 92 16 100 22
rect 72 11 77 16
rect 31 10 36 11
rect 95 10 100 16
rect 102 12 112 28
rect 102 10 105 12
rect 104 8 105 10
rect 109 10 112 12
rect 114 21 122 28
rect 114 17 116 21
rect 120 17 122 21
rect 114 10 122 17
rect 124 12 134 28
rect 124 10 127 12
rect 109 8 110 10
rect 104 7 110 8
rect 126 8 127 10
rect 131 10 134 12
rect 136 21 144 28
rect 136 17 138 21
rect 142 17 144 21
rect 136 10 144 17
rect 146 13 156 28
rect 158 21 166 28
rect 158 17 160 21
rect 164 17 166 21
rect 158 13 166 17
rect 168 19 177 28
rect 179 29 186 30
rect 179 25 181 29
rect 185 25 186 29
rect 179 24 186 25
rect 179 19 184 24
rect 168 18 175 19
rect 168 14 170 18
rect 174 14 175 18
rect 168 13 175 14
rect 146 12 154 13
rect 146 10 149 12
rect 131 8 132 10
rect 126 7 132 8
rect 148 8 149 10
rect 153 8 154 12
rect 148 7 154 8
<< pdiffusion >>
rect 2 69 9 70
rect 2 65 3 69
rect 7 65 9 69
rect 2 62 9 65
rect 2 58 3 62
rect 7 58 9 62
rect 2 42 9 58
rect 11 54 19 70
rect 11 50 13 54
rect 17 50 19 54
rect 11 47 19 50
rect 11 43 13 47
rect 17 43 19 47
rect 11 42 19 43
rect 21 69 29 70
rect 21 65 23 69
rect 27 65 29 69
rect 21 62 29 65
rect 21 58 23 62
rect 27 58 29 62
rect 21 42 29 58
rect 31 62 39 70
rect 31 58 33 62
rect 37 58 39 62
rect 31 54 39 58
rect 31 50 33 54
rect 37 50 39 54
rect 31 42 39 50
rect 41 69 49 70
rect 41 65 43 69
rect 47 65 49 69
rect 41 62 49 65
rect 41 58 43 62
rect 47 58 49 62
rect 41 42 49 58
rect 51 42 56 70
rect 58 62 66 70
rect 58 58 60 62
rect 64 58 66 62
rect 58 54 66 58
rect 58 50 60 54
rect 64 50 66 54
rect 58 42 66 50
rect 68 42 73 70
rect 75 69 83 70
rect 75 65 77 69
rect 81 65 83 69
rect 75 62 83 65
rect 75 58 77 62
rect 81 58 83 62
rect 75 42 83 58
rect 85 42 90 70
rect 92 61 100 70
rect 92 57 94 61
rect 98 57 100 61
rect 92 54 100 57
rect 92 50 94 54
rect 98 50 100 54
rect 92 42 100 50
rect 102 42 107 70
rect 109 69 117 70
rect 109 65 111 69
rect 115 65 117 69
rect 109 62 117 65
rect 109 58 111 62
rect 115 58 117 62
rect 109 42 117 58
rect 119 42 124 70
rect 126 62 134 70
rect 126 58 128 62
rect 132 58 134 62
rect 126 54 134 58
rect 126 50 128 54
rect 132 50 134 54
rect 126 42 134 50
rect 136 42 141 70
rect 143 69 151 70
rect 143 65 145 69
rect 149 65 151 69
rect 143 62 151 65
rect 143 58 145 62
rect 149 58 151 62
rect 143 42 151 58
rect 153 42 158 70
rect 160 63 165 70
rect 160 62 168 63
rect 160 58 162 62
rect 166 58 168 62
rect 160 55 168 58
rect 160 51 162 55
rect 166 51 168 55
rect 160 42 168 51
rect 170 42 175 63
rect 177 62 185 63
rect 177 58 179 62
rect 183 58 185 62
rect 177 55 185 58
rect 177 51 179 55
rect 183 51 185 55
rect 177 42 185 51
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect 118 78 122 82
rect 126 78 130 82
rect 134 78 138 82
rect 142 78 146 82
rect 150 78 154 82
rect 158 78 162 82
rect 166 78 170 82
rect 174 78 178 82
rect 182 78 186 82
rect 190 78 194 82
rect -2 69 194 78
rect -2 68 3 69
rect 2 65 3 68
rect 7 68 23 69
rect 7 65 8 68
rect 2 62 8 65
rect 2 58 3 62
rect 7 58 8 62
rect 22 65 23 68
rect 27 68 43 69
rect 27 65 28 68
rect 22 62 28 65
rect 42 65 43 68
rect 47 68 77 69
rect 47 65 48 68
rect 22 58 23 62
rect 27 58 28 62
rect 33 62 38 63
rect 37 58 38 62
rect 42 62 48 65
rect 76 65 77 68
rect 81 68 111 69
rect 81 65 82 68
rect 42 58 43 62
rect 47 58 48 62
rect 58 62 64 63
rect 58 58 60 62
rect 76 62 82 65
rect 110 65 111 68
rect 115 68 145 69
rect 115 65 116 68
rect 110 62 116 65
rect 144 65 145 68
rect 149 68 194 69
rect 149 65 150 68
rect 76 58 77 62
rect 81 58 82 62
rect 94 61 98 62
rect 33 54 38 58
rect 58 54 64 58
rect 110 58 111 62
rect 115 58 116 62
rect 128 62 134 63
rect 132 58 134 62
rect 144 62 150 65
rect 144 58 145 62
rect 149 58 150 62
rect 162 62 166 63
rect 94 54 98 57
rect 128 54 134 58
rect 162 55 166 58
rect 179 62 183 68
rect 179 55 183 58
rect 12 50 13 54
rect 17 50 33 54
rect 37 50 60 54
rect 64 50 94 54
rect 98 50 128 54
rect 132 51 162 54
rect 132 50 166 51
rect 12 47 17 50
rect 2 43 13 47
rect 170 46 174 55
rect 179 50 183 51
rect 2 42 17 43
rect 25 42 39 46
rect 78 42 183 46
rect 2 29 7 42
rect 25 38 31 42
rect 78 38 82 42
rect 110 38 116 42
rect 17 34 26 38
rect 30 34 31 38
rect 41 34 46 38
rect 50 34 77 38
rect 81 34 82 38
rect 89 34 91 38
rect 95 34 106 38
rect 110 34 111 38
rect 115 34 116 38
rect 141 38 147 42
rect 177 38 183 42
rect 124 36 128 37
rect 102 30 106 34
rect 141 34 142 38
rect 146 34 147 38
rect 153 34 161 38
rect 165 34 167 38
rect 177 34 178 38
rect 182 34 183 38
rect 124 30 128 32
rect 153 30 159 34
rect 2 25 3 29
rect 12 25 13 29
rect 17 25 33 29
rect 37 26 98 29
rect 102 26 159 30
rect 37 25 74 26
rect 2 22 7 25
rect 2 18 3 22
rect 53 24 57 25
rect 7 18 23 21
rect 2 17 23 18
rect 27 17 43 21
rect 47 17 48 21
rect 78 25 94 26
rect 74 21 78 22
rect 94 21 98 22
rect 162 25 181 29
rect 185 25 186 29
rect 162 21 166 25
rect 53 19 57 20
rect 83 17 84 21
rect 88 17 89 21
rect 94 17 116 21
rect 120 17 138 21
rect 142 17 160 21
rect 164 17 166 21
rect 170 18 174 19
rect 64 16 68 17
rect 83 12 89 17
rect 170 12 174 14
rect -2 8 105 12
rect 109 8 127 12
rect 131 8 149 12
rect 153 8 194 12
rect -2 2 194 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 122 2
rect 126 -2 130 2
rect 134 -2 138 2
rect 142 -2 146 2
rect 150 -2 154 2
rect 158 -2 162 2
rect 166 -2 170 2
rect 174 -2 178 2
rect 182 -2 186 2
rect 190 -2 194 2
<< ntransistor >>
rect 9 10 11 30
rect 19 10 21 30
rect 29 10 31 30
rect 39 11 41 30
rect 49 11 51 25
rect 59 11 61 29
rect 70 11 72 29
rect 80 16 82 29
rect 90 16 92 28
rect 100 10 102 28
rect 112 10 114 28
rect 122 10 124 28
rect 134 10 136 28
rect 144 10 146 28
rect 156 13 158 28
rect 166 13 168 28
rect 177 19 179 30
<< ptransistor >>
rect 9 42 11 70
rect 19 42 21 70
rect 29 42 31 70
rect 39 42 41 70
rect 49 42 51 70
rect 56 42 58 70
rect 66 42 68 70
rect 73 42 75 70
rect 83 42 85 70
rect 90 42 92 70
rect 100 42 102 70
rect 107 42 109 70
rect 117 42 119 70
rect 124 42 126 70
rect 134 42 136 70
rect 141 42 143 70
rect 151 42 153 70
rect 158 42 160 70
rect 168 42 170 63
rect 175 42 177 63
<< polycontact >>
rect 26 34 30 38
rect 46 34 50 38
rect 77 34 81 38
rect 91 34 95 38
rect 111 34 115 38
rect 124 32 128 36
rect 142 34 146 38
rect 161 34 165 38
rect 178 34 182 38
<< ndcontact >>
rect 3 25 7 29
rect 3 18 7 22
rect 13 25 17 29
rect 23 17 27 21
rect 33 25 37 29
rect 43 17 47 21
rect 53 20 57 24
rect 64 12 68 16
rect 74 22 78 26
rect 84 17 88 21
rect 94 22 98 26
rect 105 8 109 12
rect 116 17 120 21
rect 127 8 131 12
rect 138 17 142 21
rect 160 17 164 21
rect 181 25 185 29
rect 170 14 174 18
rect 149 8 153 12
<< pdcontact >>
rect 3 65 7 69
rect 3 58 7 62
rect 13 50 17 54
rect 13 43 17 47
rect 23 65 27 69
rect 23 58 27 62
rect 33 58 37 62
rect 33 50 37 54
rect 43 65 47 69
rect 43 58 47 62
rect 60 58 64 62
rect 60 50 64 54
rect 77 65 81 69
rect 77 58 81 62
rect 94 57 98 61
rect 94 50 98 54
rect 111 65 115 69
rect 111 58 115 62
rect 128 58 132 62
rect 128 50 132 54
rect 145 65 149 69
rect 145 58 149 62
rect 162 58 166 62
rect 162 51 166 55
rect 179 58 183 62
rect 179 51 183 55
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
rect 90 -2 94 2
rect 98 -2 102 2
rect 106 -2 110 2
rect 114 -2 118 2
rect 122 -2 126 2
rect 130 -2 134 2
rect 138 -2 142 2
rect 146 -2 150 2
rect 154 -2 158 2
rect 162 -2 166 2
rect 170 -2 174 2
rect 178 -2 182 2
rect 186 -2 190 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
rect 90 78 94 82
rect 98 78 102 82
rect 106 78 110 82
rect 114 78 118 82
rect 122 78 126 82
rect 130 78 134 82
rect 138 78 142 82
rect 146 78 150 82
rect 154 78 158 82
rect 162 78 166 82
rect 170 78 174 82
rect 178 78 182 82
rect 186 78 190 82
<< psubstratepdiff >>
rect 0 2 192 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 122 2
rect 126 -2 130 2
rect 134 -2 138 2
rect 142 -2 146 2
rect 150 -2 154 2
rect 158 -2 162 2
rect 166 -2 170 2
rect 174 -2 178 2
rect 182 -2 186 2
rect 190 -2 192 2
rect 0 -3 192 -2
<< nsubstratendiff >>
rect 0 82 192 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect 118 78 122 82
rect 126 78 130 82
rect 134 78 138 82
rect 142 78 146 82
rect 150 78 154 82
rect 158 78 162 82
rect 166 78 170 82
rect 174 78 178 82
rect 182 78 186 82
rect 190 78 192 82
rect 0 77 192 78
<< labels >>
rlabel metal1 4 32 4 32 6 z
rlabel metal1 20 36 20 36 6 b
rlabel metal1 12 44 12 44 6 z
rlabel metal1 20 52 20 52 6 z
rlabel metal1 55 24 55 24 6 n1
rlabel metal1 60 36 60 36 6 a1
rlabel metal1 52 36 52 36 6 a1
rlabel metal1 44 36 44 36 6 a1
rlabel metal1 36 44 36 44 6 b
rlabel metal1 28 40 28 40 6 b
rlabel metal1 28 52 28 52 6 z
rlabel metal1 44 52 44 52 6 z
rlabel metal1 60 56 60 56 6 z
rlabel metal1 36 56 36 56 6 z
rlabel polycontact 92 36 92 36 6 a2
rlabel metal1 76 36 76 36 6 a1
rlabel metal1 68 36 68 36 6 a1
rlabel metal1 92 44 92 44 6 a1
rlabel metal1 84 44 84 44 6 a1
rlabel metal1 92 52 92 52 6 z
rlabel metal1 84 52 84 52 6 z
rlabel metal1 76 52 76 52 6 z
rlabel metal1 68 52 68 52 6 z
rlabel metal1 96 6 96 6 6 vss
rlabel metal1 124 28 124 28 6 a2
rlabel metal1 116 28 116 28 6 a2
rlabel metal1 108 28 108 28 6 a2
rlabel ndcontact 96 23 96 23 6 n1
rlabel metal1 55 27 55 27 6 n1
rlabel metal1 100 36 100 36 6 a2
rlabel metal1 124 44 124 44 6 a1
rlabel metal1 116 44 116 44 6 a1
rlabel metal1 108 44 108 44 6 a1
rlabel metal1 100 44 100 44 6 a1
rlabel metal1 100 52 100 52 6 z
rlabel metal1 124 52 124 52 6 z
rlabel metal1 116 52 116 52 6 z
rlabel metal1 108 52 108 52 6 z
rlabel metal1 96 74 96 74 6 vdd
rlabel metal1 148 28 148 28 6 a2
rlabel metal1 140 28 140 28 6 a2
rlabel metal1 132 28 132 28 6 a2
rlabel metal1 156 32 156 32 6 a2
rlabel metal1 156 44 156 44 6 a1
rlabel metal1 148 44 148 44 6 a1
rlabel metal1 140 44 140 44 6 a1
rlabel metal1 132 44 132 44 6 a1
rlabel metal1 156 52 156 52 6 z
rlabel metal1 148 52 148 52 6 z
rlabel metal1 140 52 140 52 6 z
rlabel metal1 132 56 132 56 6 z
rlabel metal1 130 19 130 19 6 n1
rlabel metal1 174 27 174 27 6 n1
rlabel polycontact 164 36 164 36 6 a2
rlabel metal1 180 40 180 40 6 a1
rlabel metal1 164 44 164 44 6 a1
rlabel metal1 172 48 172 48 6 a1
rlabel pdcontact 164 60 164 60 6 z
<< end >>
