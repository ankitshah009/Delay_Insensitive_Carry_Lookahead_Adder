magic
tech scmos
timestamp 1179384986
<< checkpaint >>
rect -22 -22 78 94
<< ab >>
rect 0 0 56 72
<< pwell >>
rect -4 -4 60 32
<< nwell >>
rect -4 32 60 76
<< polysilicon >>
rect 9 66 11 70
rect 19 66 21 70
rect 29 63 31 68
rect 39 63 41 68
rect 9 35 11 38
rect 19 35 21 38
rect 29 35 31 38
rect 39 35 41 38
rect 9 34 22 35
rect 9 30 15 34
rect 19 30 22 34
rect 9 29 22 30
rect 28 34 34 35
rect 28 30 29 34
rect 33 30 34 34
rect 28 29 34 30
rect 10 26 12 29
rect 20 26 22 29
rect 32 26 34 29
rect 39 34 47 35
rect 39 30 42 34
rect 46 30 47 34
rect 39 29 47 30
rect 39 26 41 29
rect 10 7 12 12
rect 20 7 22 12
rect 32 2 34 6
rect 39 2 41 6
<< ndiffusion >>
rect 2 12 10 26
rect 12 18 20 26
rect 12 14 14 18
rect 18 14 20 18
rect 12 12 20 14
rect 22 12 32 26
rect 2 8 8 12
rect 2 4 3 8
rect 7 4 8 8
rect 24 11 32 12
rect 24 7 25 11
rect 29 7 32 11
rect 24 6 32 7
rect 34 6 39 26
rect 41 19 46 26
rect 41 18 48 19
rect 41 14 43 18
rect 47 14 48 18
rect 41 13 48 14
rect 41 6 46 13
rect 2 3 8 4
<< pdiffusion >>
rect 2 65 9 66
rect 2 61 3 65
rect 7 61 9 65
rect 2 58 9 61
rect 2 54 3 58
rect 7 54 9 58
rect 2 38 9 54
rect 11 58 19 66
rect 11 54 13 58
rect 17 54 19 58
rect 11 51 19 54
rect 11 47 13 51
rect 17 47 19 51
rect 11 38 19 47
rect 21 63 27 66
rect 21 62 29 63
rect 21 58 23 62
rect 27 58 29 62
rect 21 38 29 58
rect 31 58 39 63
rect 31 54 33 58
rect 37 54 39 58
rect 31 51 39 54
rect 31 47 33 51
rect 37 47 39 51
rect 31 38 39 47
rect 41 62 48 63
rect 41 58 43 62
rect 47 58 48 62
rect 41 54 48 58
rect 41 50 43 54
rect 47 50 48 54
rect 41 38 48 50
<< metal1 >>
rect -2 65 58 72
rect -2 64 3 65
rect 2 61 3 64
rect 7 64 58 65
rect 7 61 8 64
rect 2 58 8 61
rect 23 62 27 64
rect 2 54 3 58
rect 7 54 8 58
rect 13 58 17 59
rect 43 62 47 64
rect 23 57 27 58
rect 33 58 37 59
rect 13 51 17 54
rect 2 47 13 51
rect 33 51 37 54
rect 2 46 17 47
rect 23 47 33 50
rect 43 54 47 58
rect 43 49 47 50
rect 23 46 37 47
rect 2 18 6 46
rect 23 42 27 46
rect 15 38 27 42
rect 33 38 47 42
rect 15 34 19 38
rect 41 34 47 38
rect 25 30 29 34
rect 15 26 19 30
rect 33 26 37 34
rect 41 30 42 34
rect 46 30 47 34
rect 15 22 28 26
rect 33 22 47 26
rect 24 18 28 22
rect 2 14 14 18
rect 18 14 19 18
rect 24 14 43 18
rect 47 14 48 18
rect 2 13 19 14
rect 24 8 25 11
rect -2 4 3 8
rect 7 7 25 8
rect 29 8 30 11
rect 29 7 58 8
rect 7 4 58 7
rect -2 0 58 4
<< ntransistor >>
rect 10 12 12 26
rect 20 12 22 26
rect 32 6 34 26
rect 39 6 41 26
<< ptransistor >>
rect 9 38 11 66
rect 19 38 21 66
rect 29 38 31 63
rect 39 38 41 63
<< polycontact >>
rect 15 30 19 34
rect 29 30 33 34
rect 42 30 46 34
<< ndcontact >>
rect 14 14 18 18
rect 3 4 7 8
rect 25 7 29 11
rect 43 14 47 18
<< pdcontact >>
rect 3 61 7 65
rect 3 54 7 58
rect 13 54 17 58
rect 13 47 17 51
rect 23 58 27 62
rect 33 54 37 58
rect 33 47 37 51
rect 43 58 47 62
rect 43 50 47 54
<< labels >>
rlabel polysilicon 15 32 15 32 6 zn
rlabel metal1 4 32 4 32 6 z
rlabel metal1 12 16 12 16 6 z
rlabel polycontact 17 32 17 32 6 zn
rlabel metal1 12 48 12 48 6 z
rlabel metal1 28 4 28 4 6 vss
rlabel metal1 28 32 28 32 6 a
rlabel metal1 36 24 36 24 6 a
rlabel metal1 36 40 36 40 6 b
rlabel metal1 35 52 35 52 6 zn
rlabel metal1 28 68 28 68 6 vdd
rlabel metal1 36 16 36 16 6 zn
rlabel metal1 44 24 44 24 6 a
rlabel metal1 44 36 44 36 6 b
<< end >>
