magic
tech scmos
timestamp 1182081787
<< checkpaint >>
rect -25 -26 121 114
<< ab >>
rect 0 0 96 88
<< pwell >>
rect -7 -8 103 40
<< nwell >>
rect -7 40 103 96
<< polysilicon >>
rect 5 80 14 86
rect 18 80 27 86
rect 37 85 46 86
rect 37 81 41 85
rect 45 81 46 85
rect 37 80 46 81
rect 50 80 59 86
rect 69 80 78 86
rect 82 85 91 86
rect 82 81 86 85
rect 90 81 91 85
rect 82 80 91 81
rect 9 77 11 80
rect 21 77 23 80
rect 41 77 43 80
rect 53 77 55 80
rect 73 77 75 80
rect 85 77 87 80
rect 9 48 11 51
rect 21 48 23 51
rect 41 48 43 51
rect 53 48 55 51
rect 73 48 75 51
rect 85 48 87 51
rect 2 47 11 48
rect 2 43 6 47
rect 10 43 11 47
rect 2 42 11 43
rect 15 47 30 48
rect 15 43 22 47
rect 26 43 30 47
rect 15 42 30 43
rect 34 47 43 48
rect 34 43 38 47
rect 42 43 43 47
rect 34 42 43 43
rect 47 47 62 48
rect 47 43 54 47
rect 58 43 62 47
rect 47 42 62 43
rect 66 47 75 48
rect 66 43 70 47
rect 74 43 75 47
rect 66 42 75 43
rect 79 42 94 48
rect 2 37 17 38
rect 2 33 6 37
rect 10 33 17 37
rect 2 32 17 33
rect 21 37 30 38
rect 21 33 22 37
rect 26 33 30 37
rect 21 32 30 33
rect 34 37 49 38
rect 34 33 38 37
rect 42 33 49 37
rect 34 32 49 33
rect 53 37 62 38
rect 53 33 54 37
rect 58 33 62 37
rect 53 32 62 33
rect 66 37 81 38
rect 66 33 70 37
rect 74 33 81 37
rect 66 32 81 33
rect 85 32 94 38
rect 9 29 11 32
rect 21 29 23 32
rect 41 29 43 32
rect 53 29 55 32
rect 73 29 75 32
rect 85 29 87 32
rect 9 8 11 11
rect 21 8 23 11
rect 41 8 43 11
rect 53 8 55 11
rect 73 8 75 11
rect 85 8 87 11
rect 5 2 14 8
rect 18 2 27 8
rect 37 2 46 8
rect 50 2 59 8
rect 69 2 78 8
rect 82 7 91 8
rect 82 3 86 7
rect 90 3 91 7
rect 82 2 91 3
<< ndiffusion >>
rect 2 25 9 29
rect 2 21 3 25
rect 7 21 9 25
rect 2 18 9 21
rect 2 14 3 18
rect 7 14 9 18
rect 2 11 9 14
rect 11 16 21 29
rect 11 12 14 16
rect 18 12 21 16
rect 11 11 21 12
rect 23 18 30 29
rect 23 14 25 18
rect 29 14 30 18
rect 23 11 30 14
rect 34 26 41 29
rect 34 22 35 26
rect 39 22 41 26
rect 34 11 41 22
rect 43 26 53 29
rect 43 22 46 26
rect 50 22 53 26
rect 43 11 53 22
rect 55 26 62 29
rect 55 22 57 26
rect 61 22 62 26
rect 55 19 62 22
rect 55 15 57 19
rect 61 15 62 19
rect 55 11 62 15
rect 66 25 73 29
rect 66 21 67 25
rect 71 21 73 25
rect 66 18 73 21
rect 66 14 67 18
rect 71 14 73 18
rect 66 11 73 14
rect 75 17 85 29
rect 75 13 78 17
rect 82 13 85 17
rect 75 11 85 13
rect 87 11 94 29
<< pdiffusion >>
rect 2 66 9 77
rect 2 62 3 66
rect 7 62 9 66
rect 2 59 9 62
rect 2 55 3 59
rect 7 55 9 59
rect 2 51 9 55
rect 11 74 21 77
rect 11 70 14 74
rect 18 70 21 74
rect 11 67 21 70
rect 11 63 14 67
rect 18 63 21 67
rect 11 51 21 63
rect 23 73 30 77
rect 23 69 25 73
rect 29 69 30 73
rect 23 66 30 69
rect 23 62 25 66
rect 29 62 30 66
rect 23 51 30 62
rect 34 74 41 77
rect 34 70 35 74
rect 39 70 41 74
rect 34 51 41 70
rect 43 58 53 77
rect 43 54 46 58
rect 50 54 53 58
rect 43 51 53 54
rect 55 66 62 77
rect 55 62 57 66
rect 61 62 62 66
rect 55 51 62 62
rect 66 73 73 77
rect 66 69 67 73
rect 71 69 73 73
rect 66 66 73 69
rect 66 62 67 66
rect 71 62 73 66
rect 66 59 73 62
rect 66 55 67 59
rect 71 55 73 59
rect 66 51 73 55
rect 75 74 85 77
rect 75 70 78 74
rect 82 70 85 74
rect 75 67 85 70
rect 75 63 78 67
rect 82 63 85 67
rect 75 51 85 63
rect 87 51 94 77
<< metal1 >>
rect -2 86 2 90
rect 30 86 34 90
rect 2 82 30 85
rect 62 86 66 90
rect -2 81 34 82
rect 40 81 41 85
rect 45 81 58 85
rect 94 86 98 90
rect 66 82 86 85
rect 62 81 86 82
rect 90 82 94 85
rect 90 81 98 82
rect 14 74 18 81
rect 54 74 58 81
rect 78 74 82 81
rect 14 67 18 70
rect 3 66 7 67
rect 14 62 18 63
rect 25 73 35 74
rect 29 70 35 73
rect 39 70 40 74
rect 54 73 71 74
rect 54 70 67 73
rect 25 66 29 69
rect 67 66 71 69
rect 3 59 7 62
rect 25 61 29 62
rect 38 62 57 66
rect 61 62 62 66
rect 78 67 82 70
rect 78 62 82 63
rect 38 58 42 62
rect 67 59 71 62
rect 7 55 42 58
rect 3 54 42 55
rect 46 58 50 59
rect 6 47 10 51
rect 6 37 10 43
rect 6 29 10 33
rect 22 47 26 51
rect 22 37 26 43
rect 22 29 26 33
rect 38 47 42 48
rect 38 37 42 43
rect 38 32 42 33
rect 46 26 50 54
rect 54 50 58 59
rect 71 55 82 58
rect 67 54 82 55
rect 54 47 74 50
rect 58 46 70 47
rect 54 37 58 43
rect 54 32 58 33
rect 70 37 74 43
rect 70 32 74 33
rect 3 25 35 26
rect 7 22 35 25
rect 39 22 40 26
rect 46 21 50 22
rect 57 26 61 27
rect 78 26 82 54
rect 3 18 7 21
rect 57 19 61 22
rect 3 13 7 14
rect 14 16 18 17
rect 24 14 25 18
rect 29 15 57 18
rect 29 14 61 15
rect 67 25 82 26
rect 71 22 82 25
rect 67 18 71 21
rect 67 13 71 14
rect 78 17 82 18
rect 14 7 18 12
rect 78 7 82 13
rect -2 6 34 7
rect 2 3 30 6
rect -2 -2 2 2
rect 30 -2 34 2
rect 62 6 86 7
rect 66 3 86 6
rect 90 6 98 7
rect 90 3 94 6
rect 62 -2 66 2
rect 94 -2 98 2
<< metal2 >>
rect -2 86 98 90
rect 2 82 30 86
rect 34 82 62 86
rect 66 82 94 86
rect -2 80 98 82
rect -2 6 98 8
rect 2 2 30 6
rect 34 2 62 6
rect 66 2 94 6
rect -2 -2 98 2
<< ntransistor >>
rect 9 11 11 29
rect 21 11 23 29
rect 41 11 43 29
rect 53 11 55 29
rect 73 11 75 29
rect 85 11 87 29
<< ptransistor >>
rect 9 51 11 77
rect 21 51 23 77
rect 41 51 43 77
rect 53 51 55 77
rect 73 51 75 77
rect 85 51 87 77
<< polycontact >>
rect 41 81 45 85
rect 86 81 90 85
rect 6 43 10 47
rect 22 43 26 47
rect 38 43 42 47
rect 54 43 58 47
rect 70 43 74 47
rect 6 33 10 37
rect 22 33 26 37
rect 38 33 42 37
rect 54 33 58 37
rect 70 33 74 37
rect 86 3 90 7
<< ndcontact >>
rect 3 21 7 25
rect 3 14 7 18
rect 14 12 18 16
rect 25 14 29 18
rect 35 22 39 26
rect 46 22 50 26
rect 57 22 61 26
rect 57 15 61 19
rect 67 21 71 25
rect 67 14 71 18
rect 78 13 82 17
<< pdcontact >>
rect 3 62 7 66
rect 3 55 7 59
rect 14 70 18 74
rect 14 63 18 67
rect 25 69 29 73
rect 25 62 29 66
rect 35 70 39 74
rect 46 54 50 58
rect 57 62 61 66
rect 67 69 71 73
rect 67 62 71 66
rect 67 55 71 59
rect 78 70 82 74
rect 78 63 82 67
<< m2contact >>
rect -2 82 2 86
rect 30 82 34 86
rect 62 82 66 86
rect 94 82 98 86
rect -2 2 2 6
rect 30 2 34 6
rect 62 2 66 6
rect 94 2 98 6
<< psubstratepcontact >>
rect -2 2 2 6
rect 30 2 34 6
rect 62 2 66 6
rect 94 2 98 6
<< nsubstratencontact >>
rect -2 82 2 86
rect 30 82 34 86
rect 62 82 66 86
rect 94 82 98 86
<< psubstratepdiff >>
rect -3 6 3 7
rect -3 2 -2 6
rect 2 2 3 6
rect 29 6 35 7
rect 29 2 30 6
rect 34 2 35 6
rect 61 6 67 7
rect 61 2 62 6
rect 66 2 67 6
rect 93 6 99 7
rect 93 2 94 6
rect 98 2 99 6
rect -3 0 3 2
rect 29 0 35 2
rect 61 0 67 2
rect 93 0 99 2
<< nsubstratendiff >>
rect -3 86 3 88
rect 29 86 35 88
rect 61 86 67 88
rect 93 86 99 88
rect -3 82 -2 86
rect 2 82 3 86
rect -3 81 3 82
rect 29 82 30 86
rect 34 82 35 86
rect 29 81 35 82
rect 61 82 62 86
rect 66 82 67 86
rect 61 81 67 82
rect 93 82 94 86
rect 98 82 99 86
rect 93 81 99 82
<< labels >>
rlabel metal1 8 40 8 40 6 a1
rlabel metal1 24 40 24 40 6 a2
rlabel metal1 48 40 48 40 6 z
rlabel metal1 56 48 56 48 6 s
rlabel metal1 72 40 72 40 6 s
rlabel metal1 64 48 64 48 6 s
rlabel metal2 48 4 48 4 6 vss
rlabel metal2 48 84 48 84 6 vdd
<< end >>
