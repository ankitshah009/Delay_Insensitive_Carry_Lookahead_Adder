magic
tech scmos
timestamp 1179386141
<< checkpaint >>
rect -22 -25 86 105
<< ab >>
rect 0 0 64 80
<< pwell >>
rect -4 -7 68 36
<< nwell >>
rect -4 36 68 87
<< polysilicon >>
rect 9 62 11 67
rect 19 62 21 67
rect 26 62 28 67
rect 36 62 38 67
rect 43 62 45 67
rect 56 56 62 57
rect 56 53 57 56
rect 9 31 11 50
rect 19 41 21 50
rect 16 40 22 41
rect 16 36 17 40
rect 21 36 22 40
rect 16 35 22 36
rect 26 37 28 50
rect 36 47 38 50
rect 33 46 39 47
rect 33 42 34 46
rect 38 42 39 46
rect 33 41 39 42
rect 43 39 45 50
rect 53 52 57 53
rect 61 52 62 56
rect 53 51 62 52
rect 53 48 55 51
rect 43 38 49 39
rect 26 35 38 37
rect 8 30 14 31
rect 8 26 9 30
rect 13 26 14 30
rect 8 25 14 26
rect 9 22 11 25
rect 19 22 21 35
rect 26 30 32 31
rect 26 26 27 30
rect 31 26 32 30
rect 26 25 32 26
rect 26 22 28 25
rect 36 22 38 35
rect 43 34 44 38
rect 48 34 49 38
rect 43 33 49 34
rect 43 22 45 33
rect 53 22 55 42
rect 9 11 11 16
rect 19 11 21 16
rect 26 11 28 16
rect 36 8 38 16
rect 43 12 45 16
rect 53 8 55 16
rect 36 6 55 8
<< ndiffusion >>
rect 2 21 9 22
rect 2 17 3 21
rect 7 17 9 21
rect 2 16 9 17
rect 11 21 19 22
rect 11 17 13 21
rect 17 17 19 21
rect 11 16 19 17
rect 21 16 26 22
rect 28 21 36 22
rect 28 17 30 21
rect 34 17 36 21
rect 28 16 36 17
rect 38 16 43 22
rect 45 21 53 22
rect 45 17 47 21
rect 51 17 53 21
rect 45 16 53 17
rect 55 21 62 22
rect 55 17 57 21
rect 61 17 62 21
rect 55 16 62 17
<< pdiffusion >>
rect 4 56 9 62
rect 2 55 9 56
rect 2 51 3 55
rect 7 51 9 55
rect 2 50 9 51
rect 11 61 19 62
rect 11 57 13 61
rect 17 57 19 61
rect 11 50 19 57
rect 21 50 26 62
rect 28 55 36 62
rect 28 51 30 55
rect 34 51 36 55
rect 28 50 36 51
rect 38 50 43 62
rect 45 61 52 62
rect 45 57 47 61
rect 51 57 52 61
rect 45 56 52 57
rect 45 50 51 56
rect 47 48 51 50
rect 47 42 53 48
rect 55 47 62 48
rect 55 43 57 47
rect 61 43 62 47
rect 55 42 62 43
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect -2 68 66 78
rect 12 61 18 68
rect 12 57 13 61
rect 17 57 18 61
rect 46 61 52 68
rect 46 57 47 61
rect 51 57 52 61
rect 57 56 62 63
rect 2 51 3 55
rect 7 54 8 55
rect 29 54 30 55
rect 7 51 15 54
rect 2 50 15 51
rect 18 51 30 54
rect 34 51 35 55
rect 18 50 35 51
rect 49 52 57 54
rect 61 52 62 56
rect 49 50 62 52
rect 2 21 6 50
rect 18 47 22 50
rect 9 43 22 47
rect 34 46 57 47
rect 9 30 13 43
rect 25 40 31 46
rect 16 36 17 40
rect 21 36 31 40
rect 16 34 31 36
rect 38 43 57 46
rect 61 43 62 47
rect 34 31 38 42
rect 27 30 38 31
rect 13 26 24 29
rect 9 25 24 26
rect 31 26 38 30
rect 27 25 38 26
rect 42 38 48 39
rect 42 34 44 38
rect 42 31 48 34
rect 42 25 54 31
rect 13 21 17 22
rect 2 17 3 21
rect 7 17 8 21
rect 20 21 24 25
rect 58 21 62 43
rect 20 17 30 21
rect 34 17 35 21
rect 46 17 47 21
rect 51 17 52 21
rect 56 17 57 21
rect 61 17 62 21
rect 13 12 17 17
rect 46 12 52 17
rect -2 2 66 12
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
<< ntransistor >>
rect 9 16 11 22
rect 19 16 21 22
rect 26 16 28 22
rect 36 16 38 22
rect 43 16 45 22
rect 53 16 55 22
<< ptransistor >>
rect 9 50 11 62
rect 19 50 21 62
rect 26 50 28 62
rect 36 50 38 62
rect 43 50 45 62
rect 53 42 55 48
<< polycontact >>
rect 17 36 21 40
rect 34 42 38 46
rect 57 52 61 56
rect 9 26 13 30
rect 27 26 31 30
rect 44 34 48 38
<< ndcontact >>
rect 3 17 7 21
rect 13 17 17 21
rect 30 17 34 21
rect 47 17 51 21
rect 57 17 61 21
<< pdcontact >>
rect 3 51 7 55
rect 13 57 17 61
rect 30 51 34 55
rect 47 57 51 61
rect 57 43 61 47
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
<< psubstratepdiff >>
rect 0 2 64 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 64 2
rect 0 -3 64 -2
<< nsubstratendiff >>
rect 0 82 64 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 64 82
rect 0 77 64 78
<< labels >>
rlabel polysilicon 10 39 10 39 6 zn
rlabel polycontact 29 28 29 28 6 sn
rlabel ptransistor 37 54 37 54 6 sn
rlabel metal1 4 36 4 36 6 z
rlabel metal1 11 36 11 36 6 zn
rlabel metal1 20 36 20 36 6 a0
rlabel metal1 12 52 12 52 6 z
rlabel metal1 32 6 32 6 6 vss
rlabel metal1 27 19 27 19 6 zn
rlabel metal1 36 36 36 36 6 sn
rlabel metal1 32 28 32 28 6 sn
rlabel metal1 28 40 28 40 6 a0
rlabel metal1 26 52 26 52 6 zn
rlabel metal1 32 74 32 74 6 vdd
rlabel metal1 44 32 44 32 6 a1
rlabel metal1 52 28 52 28 6 a1
rlabel metal1 60 32 60 32 6 sn
rlabel metal1 48 45 48 45 6 sn
rlabel metal1 52 52 52 52 6 s
rlabel metal1 60 60 60 60 6 s
<< end >>
