magic
tech scmos
timestamp 1179387560
<< checkpaint >>
rect -22 -22 206 94
<< ab >>
rect 0 0 184 72
<< pwell >>
rect -4 -4 188 32
<< nwell >>
rect -4 32 188 76
<< polysilicon >>
rect 9 65 11 70
rect 19 65 21 70
rect 29 68 53 70
rect 29 65 31 68
rect 39 65 41 68
rect 51 51 53 68
rect 63 66 65 70
rect 73 66 75 70
rect 83 66 85 70
rect 93 66 95 70
rect 116 66 118 70
rect 123 66 125 70
rect 133 66 135 70
rect 151 66 153 70
rect 161 66 163 70
rect 48 50 54 51
rect 48 46 49 50
rect 53 46 54 50
rect 48 45 54 46
rect 9 35 11 38
rect 19 35 21 38
rect 29 35 31 38
rect 39 35 41 38
rect 63 37 65 40
rect 73 37 75 40
rect 9 34 22 35
rect 9 33 17 34
rect 16 30 17 33
rect 21 30 22 34
rect 29 33 41 35
rect 61 35 75 37
rect 83 35 85 38
rect 93 35 95 38
rect 116 35 118 38
rect 61 34 67 35
rect 16 29 22 30
rect 9 24 11 29
rect 16 27 28 29
rect 16 24 18 27
rect 26 24 28 27
rect 33 24 35 33
rect 61 31 62 34
rect 45 26 47 31
rect 55 30 62 31
rect 66 30 67 34
rect 80 34 108 35
rect 80 33 103 34
rect 80 31 82 33
rect 55 29 67 30
rect 55 26 57 29
rect 65 26 67 29
rect 75 29 82 31
rect 102 30 103 33
rect 107 30 108 34
rect 102 29 108 30
rect 112 34 118 35
rect 112 30 113 34
rect 117 30 118 34
rect 123 35 125 38
rect 133 35 135 38
rect 151 35 153 38
rect 161 35 163 38
rect 123 32 126 35
rect 133 34 153 35
rect 133 33 138 34
rect 112 29 118 30
rect 75 26 77 29
rect 86 27 92 28
rect 86 23 87 27
rect 91 23 92 27
rect 114 26 116 29
rect 124 26 126 32
rect 137 30 138 33
rect 142 33 153 34
rect 157 34 163 35
rect 142 30 148 33
rect 137 29 148 30
rect 157 30 158 34
rect 162 30 163 34
rect 157 29 163 30
rect 146 26 148 29
rect 85 21 97 23
rect 85 18 87 21
rect 95 18 97 21
rect 9 4 11 12
rect 16 8 18 12
rect 26 8 28 12
rect 33 4 35 12
rect 9 2 35 4
rect 45 4 47 12
rect 55 8 57 12
rect 65 8 67 12
rect 75 4 77 12
rect 133 17 139 18
rect 133 13 134 17
rect 138 13 139 17
rect 158 23 160 29
rect 133 12 139 13
rect 45 2 77 4
rect 85 2 87 6
rect 95 2 97 6
rect 114 7 116 12
rect 124 9 126 12
rect 133 9 135 12
rect 146 10 148 15
rect 124 7 135 9
rect 158 7 160 12
<< ndiffusion >>
rect 37 24 45 26
rect 4 18 9 24
rect 2 17 9 18
rect 2 13 3 17
rect 7 13 9 17
rect 2 12 9 13
rect 11 12 16 24
rect 18 23 26 24
rect 18 19 20 23
rect 24 19 26 23
rect 18 12 26 19
rect 28 12 33 24
rect 35 12 45 24
rect 47 25 55 26
rect 47 21 49 25
rect 53 21 55 25
rect 47 12 55 21
rect 57 17 65 26
rect 57 13 59 17
rect 63 13 65 17
rect 57 12 65 13
rect 67 25 75 26
rect 67 21 69 25
rect 73 21 75 25
rect 67 18 75 21
rect 67 14 69 18
rect 73 14 75 18
rect 67 12 75 14
rect 77 18 82 26
rect 109 19 114 26
rect 107 18 114 19
rect 77 17 85 18
rect 77 13 79 17
rect 83 13 85 17
rect 77 12 85 13
rect 37 8 43 12
rect 37 4 38 8
rect 42 4 43 8
rect 37 3 43 4
rect 80 6 85 12
rect 87 17 95 18
rect 87 13 89 17
rect 93 13 95 17
rect 87 6 95 13
rect 97 9 103 18
rect 107 14 108 18
rect 112 14 114 18
rect 107 13 114 14
rect 109 12 114 13
rect 116 25 124 26
rect 116 21 118 25
rect 122 21 124 25
rect 116 12 124 21
rect 126 25 133 26
rect 126 21 128 25
rect 132 21 133 25
rect 126 20 133 21
rect 139 25 146 26
rect 139 21 140 25
rect 144 21 146 25
rect 139 20 146 21
rect 126 12 131 20
rect 141 15 146 20
rect 148 23 156 26
rect 148 15 158 23
rect 97 8 105 9
rect 97 6 100 8
rect 99 4 100 6
rect 104 4 105 8
rect 150 12 158 15
rect 160 18 165 23
rect 160 17 167 18
rect 160 13 162 17
rect 166 13 167 17
rect 160 12 167 13
rect 99 3 105 4
rect 150 8 156 12
rect 150 4 151 8
rect 155 4 156 8
rect 150 3 156 4
<< pdiffusion >>
rect 4 59 9 65
rect 2 58 9 59
rect 2 54 3 58
rect 7 54 9 58
rect 2 51 9 54
rect 2 47 3 51
rect 7 47 9 51
rect 2 46 9 47
rect 4 38 9 46
rect 11 50 19 65
rect 11 46 13 50
rect 17 46 19 50
rect 11 43 19 46
rect 11 39 13 43
rect 17 39 19 43
rect 11 38 19 39
rect 21 58 29 65
rect 21 54 23 58
rect 27 54 29 58
rect 21 38 29 54
rect 31 43 39 65
rect 31 39 33 43
rect 37 39 39 43
rect 31 38 39 39
rect 41 59 46 65
rect 41 58 48 59
rect 41 54 43 58
rect 47 54 48 58
rect 41 53 48 54
rect 41 38 46 53
rect 56 65 63 66
rect 56 61 57 65
rect 61 61 63 65
rect 56 58 63 61
rect 56 54 57 58
rect 61 54 63 58
rect 56 40 63 54
rect 65 58 73 66
rect 65 54 67 58
rect 71 54 73 58
rect 65 51 73 54
rect 65 47 67 51
rect 71 47 73 51
rect 65 40 73 47
rect 75 65 83 66
rect 75 61 77 65
rect 81 61 83 65
rect 75 40 83 61
rect 78 38 83 40
rect 85 45 93 66
rect 85 41 87 45
rect 91 41 93 45
rect 85 38 93 41
rect 95 65 116 66
rect 95 61 97 65
rect 101 61 105 65
rect 109 61 116 65
rect 95 58 116 61
rect 95 54 105 58
rect 109 54 116 58
rect 95 38 116 54
rect 118 38 123 66
rect 125 59 133 66
rect 125 55 127 59
rect 131 55 133 59
rect 125 38 133 55
rect 135 60 140 66
rect 135 59 142 60
rect 135 55 137 59
rect 141 55 142 59
rect 135 54 142 55
rect 135 38 140 54
rect 146 50 151 66
rect 144 49 151 50
rect 144 45 145 49
rect 149 45 151 49
rect 144 44 151 45
rect 146 38 151 44
rect 153 65 161 66
rect 153 61 155 65
rect 159 61 161 65
rect 153 38 161 61
rect 163 51 168 66
rect 163 50 170 51
rect 163 46 165 50
rect 169 46 170 50
rect 163 43 170 46
rect 163 39 165 43
rect 169 39 170 43
rect 163 38 170 39
<< metal1 >>
rect -2 68 186 72
rect -2 65 173 68
rect -2 64 57 65
rect 56 61 57 64
rect 61 64 77 65
rect 61 61 62 64
rect 56 58 62 61
rect 81 64 97 65
rect 77 60 81 61
rect 101 64 105 65
rect 97 60 101 61
rect 109 64 155 65
rect 154 61 155 64
rect 159 64 173 65
rect 177 64 186 68
rect 159 61 160 64
rect 2 54 3 58
rect 7 54 23 58
rect 27 54 43 58
rect 47 54 48 58
rect 56 54 57 58
rect 61 54 62 58
rect 67 58 71 59
rect 105 58 109 61
rect 2 51 7 54
rect 2 47 3 51
rect 67 51 99 54
rect 105 53 109 54
rect 113 55 127 59
rect 131 55 132 59
rect 136 55 137 59
rect 141 58 142 59
rect 141 55 169 58
rect 2 46 7 47
rect 12 46 13 50
rect 17 46 49 50
rect 53 47 67 50
rect 71 50 99 51
rect 53 46 71 47
rect 2 26 6 46
rect 12 43 17 46
rect 87 45 91 46
rect 12 39 13 43
rect 12 38 17 39
rect 32 39 33 43
rect 37 39 38 43
rect 32 34 38 39
rect 48 41 87 42
rect 48 38 91 41
rect 48 34 52 38
rect 16 30 17 34
rect 21 30 52 34
rect 57 30 62 34
rect 66 30 87 34
rect 2 23 24 26
rect 2 22 20 23
rect 48 25 52 30
rect 81 28 87 30
rect 81 27 91 28
rect 48 21 49 25
rect 53 21 69 25
rect 73 21 74 25
rect 81 23 87 27
rect 81 22 91 23
rect 20 18 24 19
rect 69 18 74 21
rect 3 17 7 18
rect 20 17 64 18
rect 20 14 59 17
rect 58 13 59 14
rect 63 13 64 17
rect 73 14 74 18
rect 95 17 99 50
rect 113 49 117 55
rect 136 54 169 55
rect 103 45 117 49
rect 121 45 145 49
rect 149 45 150 49
rect 103 34 107 45
rect 121 34 125 45
rect 129 38 142 42
rect 138 34 142 38
rect 154 35 158 51
rect 165 50 169 54
rect 165 43 169 46
rect 112 30 113 34
rect 117 30 131 34
rect 103 25 107 30
rect 127 25 131 30
rect 138 29 142 30
rect 146 34 162 35
rect 146 30 158 34
rect 146 29 162 30
rect 103 21 118 25
rect 122 21 123 25
rect 127 21 128 25
rect 132 21 140 25
rect 144 21 145 25
rect 154 21 158 29
rect 69 13 74 14
rect 78 13 79 17
rect 83 13 84 17
rect 88 13 89 17
rect 93 13 99 17
rect 107 14 108 18
rect 112 17 113 18
rect 165 17 169 39
rect 112 14 134 17
rect 107 13 134 14
rect 138 13 162 17
rect 166 13 169 17
rect 3 8 7 13
rect 78 8 84 13
rect -2 4 38 8
rect 42 4 100 8
rect 104 4 138 8
rect 142 4 151 8
rect 155 4 172 8
rect 176 4 186 8
rect -2 0 186 4
<< ntransistor >>
rect 9 12 11 24
rect 16 12 18 24
rect 26 12 28 24
rect 33 12 35 24
rect 45 12 47 26
rect 55 12 57 26
rect 65 12 67 26
rect 75 12 77 26
rect 85 6 87 18
rect 95 6 97 18
rect 114 12 116 26
rect 124 12 126 26
rect 146 15 148 26
rect 158 12 160 23
<< ptransistor >>
rect 9 38 11 65
rect 19 38 21 65
rect 29 38 31 65
rect 39 38 41 65
rect 63 40 65 66
rect 73 40 75 66
rect 83 38 85 66
rect 93 38 95 66
rect 116 38 118 66
rect 123 38 125 66
rect 133 38 135 66
rect 151 38 153 66
rect 161 38 163 66
<< polycontact >>
rect 49 46 53 50
rect 17 30 21 34
rect 62 30 66 34
rect 103 30 107 34
rect 113 30 117 34
rect 87 23 91 27
rect 138 30 142 34
rect 158 30 162 34
rect 134 13 138 17
<< ndcontact >>
rect 3 13 7 17
rect 20 19 24 23
rect 49 21 53 25
rect 59 13 63 17
rect 69 21 73 25
rect 69 14 73 18
rect 79 13 83 17
rect 38 4 42 8
rect 89 13 93 17
rect 108 14 112 18
rect 118 21 122 25
rect 128 21 132 25
rect 140 21 144 25
rect 100 4 104 8
rect 162 13 166 17
rect 151 4 155 8
<< pdcontact >>
rect 3 54 7 58
rect 3 47 7 51
rect 13 46 17 50
rect 13 39 17 43
rect 23 54 27 58
rect 33 39 37 43
rect 43 54 47 58
rect 57 61 61 65
rect 57 54 61 58
rect 67 54 71 58
rect 67 47 71 51
rect 77 61 81 65
rect 87 41 91 45
rect 97 61 101 65
rect 105 61 109 65
rect 105 54 109 58
rect 127 55 131 59
rect 137 55 141 59
rect 145 45 149 49
rect 155 61 159 65
rect 165 46 169 50
rect 165 39 169 43
<< psubstratepcontact >>
rect 138 4 142 8
rect 172 4 176 8
<< nsubstratencontact >>
rect 173 64 177 68
<< psubstratepdiff >>
rect 137 8 143 9
rect 137 4 138 8
rect 142 4 143 8
rect 137 3 143 4
rect 171 8 177 26
rect 171 4 172 8
rect 176 4 177 8
rect 171 3 177 4
<< nsubstratendiff >>
rect 172 68 178 69
rect 172 64 173 68
rect 177 64 178 68
rect 172 55 178 64
<< labels >>
rlabel ptransistor 20 48 20 48 6 zn
rlabel polysilicon 52 57 52 57 6 cn
rlabel ntransistor 115 21 115 21 6 bn
rlabel polycontact 105 32 105 32 6 iz
rlabel polycontact 136 15 136 15 6 an
rlabel metal1 28 16 28 16 6 z
rlabel metal1 20 24 20 24 6 z
rlabel metal1 12 24 12 24 6 z
rlabel metal1 4 40 4 40 6 z
rlabel metal1 14 44 14 44 6 cn
rlabel metal1 28 56 28 56 6 z
rlabel metal1 20 56 20 56 6 z
rlabel metal1 12 56 12 56 6 z
rlabel ndcontact 60 16 60 16 6 z
rlabel metal1 52 16 52 16 6 z
rlabel metal1 44 16 44 16 6 z
rlabel metal1 36 16 36 16 6 z
rlabel metal1 68 32 68 32 6 c
rlabel metal1 60 32 60 32 6 c
rlabel metal1 35 36 35 36 6 zn
rlabel metal1 41 48 41 48 6 cn
rlabel pdcontact 44 56 44 56 6 z
rlabel metal1 36 56 36 56 6 z
rlabel metal1 92 4 92 4 6 vss
rlabel metal1 93 15 93 15 6 cn
rlabel metal1 71 19 71 19 6 zn
rlabel metal1 61 23 61 23 6 zn
rlabel metal1 84 28 84 28 6 c
rlabel metal1 76 32 76 32 6 c
rlabel pdcontact 89 42 89 42 6 zn
rlabel metal1 105 35 105 35 6 iz
rlabel metal1 83 52 83 52 6 cn
rlabel metal1 92 68 92 68 6 vdd
rlabel metal1 113 23 113 23 6 iz
rlabel metal1 136 23 136 23 6 bn
rlabel polycontact 140 32 140 32 6 b
rlabel metal1 132 40 132 40 6 b
rlabel metal1 123 39 123 39 6 bn
rlabel pdcontact 139 56 139 56 6 an
rlabel metal1 122 57 122 57 6 iz
rlabel metal1 138 15 138 15 6 an
rlabel metal1 156 24 156 24 6 a
rlabel metal1 148 32 148 32 6 a
rlabel metal1 156 36 156 36 6 a
rlabel metal1 135 47 135 47 6 bn
rlabel metal1 167 35 167 35 6 an
<< end >>
