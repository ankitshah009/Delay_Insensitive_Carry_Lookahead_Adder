magic
tech scmos
timestamp 1179386522
<< checkpaint >>
rect -22 -25 78 105
<< ab >>
rect 0 0 56 80
<< pwell >>
rect -4 -7 60 36
<< nwell >>
rect -4 36 60 87
<< polysilicon >>
rect 9 60 11 65
rect 21 60 23 65
rect 31 60 33 65
rect 45 64 47 69
rect 9 32 11 50
rect 21 39 23 50
rect 31 39 33 50
rect 45 49 47 52
rect 41 48 47 49
rect 41 44 42 48
rect 46 44 47 48
rect 41 43 47 44
rect 19 38 25 39
rect 19 34 20 38
rect 24 34 25 38
rect 19 33 25 34
rect 31 38 41 39
rect 31 34 36 38
rect 40 34 41 38
rect 31 33 41 34
rect 9 31 15 32
rect 9 27 10 31
rect 14 29 15 31
rect 14 27 17 29
rect 9 26 17 27
rect 15 23 17 26
rect 22 23 24 33
rect 31 29 33 33
rect 45 30 47 43
rect 29 26 33 29
rect 29 23 31 26
rect 45 19 47 24
rect 15 8 17 13
rect 22 8 24 13
rect 29 8 31 13
<< ndiffusion >>
rect 35 24 45 30
rect 47 29 54 30
rect 47 25 49 29
rect 53 25 54 29
rect 47 24 54 25
rect 35 23 43 24
rect 8 21 15 23
rect 8 17 9 21
rect 13 17 15 21
rect 8 16 15 17
rect 10 13 15 16
rect 17 13 22 23
rect 24 13 29 23
rect 31 20 43 23
rect 31 16 36 20
rect 40 16 43 20
rect 31 13 43 16
<< pdiffusion >>
rect 35 60 45 64
rect 4 56 9 60
rect 2 55 9 56
rect 2 51 3 55
rect 7 51 9 55
rect 2 50 9 51
rect 11 59 21 60
rect 11 55 14 59
rect 18 55 21 59
rect 11 50 21 55
rect 23 55 31 60
rect 23 51 25 55
rect 29 51 31 55
rect 23 50 31 51
rect 33 59 45 60
rect 33 55 35 59
rect 39 55 45 59
rect 33 52 45 55
rect 47 58 52 64
rect 47 57 54 58
rect 47 53 49 57
rect 53 53 54 57
rect 47 52 54 53
rect 33 50 39 52
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect -2 68 58 78
rect 14 59 18 68
rect 2 55 7 56
rect 2 51 3 55
rect 35 59 39 68
rect 14 54 18 55
rect 25 55 29 56
rect 2 46 7 51
rect 35 54 39 55
rect 25 46 29 51
rect 42 48 46 63
rect 2 42 29 46
rect 33 44 42 46
rect 33 42 46 44
rect 49 57 53 58
rect 2 21 6 42
rect 49 38 53 53
rect 19 34 20 38
rect 24 34 31 38
rect 35 34 36 38
rect 40 34 53 38
rect 10 31 14 32
rect 26 31 31 34
rect 14 27 22 29
rect 10 25 22 27
rect 26 25 38 31
rect 49 29 53 34
rect 2 17 9 21
rect 13 17 14 21
rect 18 17 22 25
rect 49 24 53 25
rect 36 20 40 21
rect 36 12 40 16
rect -2 2 58 12
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
<< ntransistor >>
rect 45 24 47 30
rect 15 13 17 23
rect 22 13 24 23
rect 29 13 31 23
<< ptransistor >>
rect 9 50 11 60
rect 21 50 23 60
rect 31 50 33 60
rect 45 52 47 64
<< polycontact >>
rect 42 44 46 48
rect 20 34 24 38
rect 36 34 40 38
rect 10 27 14 31
<< ndcontact >>
rect 49 25 53 29
rect 9 17 13 21
rect 36 16 40 20
<< pdcontact >>
rect 3 51 7 55
rect 14 55 18 59
rect 25 51 29 55
rect 35 55 39 59
rect 49 53 53 57
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
<< psubstratepdiff >>
rect 0 2 56 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 56 2
rect 0 -3 56 -2
<< nsubstratendiff >>
rect 0 82 56 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 56 82
rect 0 77 56 78
<< labels >>
rlabel polysilicon 36 36 36 36 6 an
rlabel metal1 4 36 4 36 6 z
rlabel metal1 20 20 20 20 6 c
rlabel polycontact 12 28 12 28 6 c
rlabel metal1 20 44 20 44 6 z
rlabel metal1 12 44 12 44 6 z
rlabel metal1 28 6 28 6 6 vss
rlabel metal1 28 32 28 32 6 b
rlabel metal1 36 28 36 28 6 b
rlabel metal1 36 44 36 44 6 a
rlabel metal1 28 74 28 74 6 vdd
rlabel metal1 44 36 44 36 6 an
rlabel metal1 51 41 51 41 6 an
rlabel metal1 44 56 44 56 6 a
<< end >>
