magic
tech scmos
timestamp 1185038975
<< checkpaint >>
rect -22 -24 112 124
<< ab >>
rect 0 0 90 100
<< pwell >>
rect -2 -4 92 49
<< nwell >>
rect -2 49 92 104
<< polysilicon >>
rect 75 95 77 98
rect 11 85 13 88
rect 23 85 25 88
rect 31 85 33 88
rect 47 85 49 88
rect 55 85 57 88
rect 11 41 13 65
rect 23 63 25 65
rect 17 62 25 63
rect 17 58 18 62
rect 22 61 25 62
rect 22 58 23 61
rect 17 57 23 58
rect 31 43 33 65
rect 47 57 49 65
rect 55 63 57 65
rect 55 62 63 63
rect 55 61 58 62
rect 57 58 58 61
rect 62 58 63 62
rect 57 57 63 58
rect 47 56 53 57
rect 47 52 48 56
rect 52 52 53 56
rect 47 51 53 52
rect 37 50 43 51
rect 37 46 38 50
rect 42 47 43 50
rect 75 47 77 55
rect 42 46 77 47
rect 37 45 77 46
rect 27 42 33 43
rect 27 41 28 42
rect 11 39 28 41
rect 11 15 13 39
rect 27 38 28 39
rect 32 41 33 42
rect 32 39 49 41
rect 32 38 33 39
rect 27 37 33 38
rect 17 32 23 33
rect 17 28 18 32
rect 22 29 23 32
rect 22 28 25 29
rect 17 27 25 28
rect 23 15 25 27
rect 29 22 35 23
rect 29 18 30 22
rect 34 18 35 22
rect 29 17 35 18
rect 31 15 33 17
rect 47 15 49 39
rect 57 32 63 33
rect 57 29 58 32
rect 55 28 58 29
rect 62 28 63 32
rect 55 27 63 28
rect 55 15 57 27
rect 75 25 77 45
rect 11 2 13 5
rect 23 2 25 5
rect 31 2 33 5
rect 47 2 49 5
rect 55 2 57 5
rect 75 2 77 5
<< ndiffusion >>
rect 3 22 9 25
rect 3 18 4 22
rect 8 18 9 22
rect 3 15 9 18
rect 37 32 45 33
rect 37 28 38 32
rect 42 28 45 32
rect 37 15 45 28
rect 59 22 75 25
rect 59 18 68 22
rect 72 18 75 22
rect 59 15 75 18
rect 3 5 11 15
rect 13 12 23 15
rect 13 8 16 12
rect 20 8 23 12
rect 13 5 23 8
rect 25 5 31 15
rect 33 5 47 15
rect 49 5 55 15
rect 57 12 75 15
rect 57 8 68 12
rect 72 8 75 12
rect 57 5 75 8
rect 77 22 85 25
rect 77 18 80 22
rect 84 18 85 22
rect 77 5 85 18
<< pdiffusion >>
rect 15 92 21 93
rect 15 88 16 92
rect 20 88 21 92
rect 59 92 75 95
rect 59 88 68 92
rect 72 88 75 92
rect 15 85 21 88
rect 59 85 75 88
rect 3 82 11 85
rect 3 78 4 82
rect 8 78 11 82
rect 3 72 11 78
rect 3 68 4 72
rect 8 68 11 72
rect 3 65 11 68
rect 13 65 23 85
rect 25 65 31 85
rect 33 82 47 85
rect 33 78 38 82
rect 42 78 47 82
rect 33 72 47 78
rect 33 68 38 72
rect 42 68 47 72
rect 33 65 47 68
rect 49 65 55 85
rect 57 82 75 85
rect 57 78 68 82
rect 72 78 75 82
rect 57 72 75 78
rect 57 68 68 72
rect 72 68 75 72
rect 57 65 75 68
rect 67 62 75 65
rect 67 58 68 62
rect 72 58 75 62
rect 67 55 75 58
rect 77 82 85 95
rect 77 78 80 82
rect 84 78 85 82
rect 77 72 85 78
rect 77 68 80 72
rect 84 68 85 72
rect 77 62 85 68
rect 77 58 80 62
rect 84 58 85 62
rect 77 55 85 58
<< metal1 >>
rect -2 96 92 101
rect -2 92 28 96
rect 32 92 38 96
rect 42 92 48 96
rect 52 92 92 96
rect -2 88 16 92
rect 20 88 68 92
rect 72 88 92 92
rect -2 87 92 88
rect 3 82 9 83
rect 37 82 43 83
rect 67 82 73 87
rect 3 78 4 82
rect 8 78 9 82
rect 3 77 9 78
rect 4 73 8 77
rect 3 72 9 73
rect 3 68 4 72
rect 8 68 9 72
rect 3 67 9 68
rect 4 23 8 67
rect 17 62 23 82
rect 17 58 18 62
rect 22 58 23 62
rect 17 32 23 58
rect 17 28 18 32
rect 22 28 23 32
rect 27 42 33 82
rect 37 78 38 82
rect 42 78 43 82
rect 37 77 43 78
rect 38 73 42 77
rect 37 72 43 73
rect 37 68 38 72
rect 42 68 43 72
rect 37 67 43 68
rect 38 51 42 67
rect 57 62 63 82
rect 57 58 58 62
rect 62 58 63 62
rect 47 56 53 57
rect 47 52 48 56
rect 52 52 53 56
rect 47 51 53 52
rect 37 50 43 51
rect 37 46 38 50
rect 42 46 43 50
rect 37 45 43 46
rect 27 38 28 42
rect 32 38 33 42
rect 27 28 33 38
rect 38 33 42 45
rect 37 32 43 33
rect 37 28 38 32
rect 42 28 43 32
rect 17 27 23 28
rect 37 27 43 28
rect 3 22 9 23
rect 29 22 35 23
rect 48 22 52 51
rect 3 18 4 22
rect 8 18 30 22
rect 34 18 52 22
rect 57 32 63 58
rect 67 78 68 82
rect 72 78 73 82
rect 67 72 73 78
rect 67 68 68 72
rect 72 68 73 72
rect 67 62 73 68
rect 67 58 68 62
rect 72 58 73 62
rect 67 57 73 58
rect 77 82 85 83
rect 77 78 80 82
rect 84 78 85 82
rect 77 77 85 78
rect 77 73 83 77
rect 77 72 85 73
rect 77 68 80 72
rect 84 68 85 72
rect 77 67 85 68
rect 77 63 83 67
rect 77 62 85 63
rect 77 58 80 62
rect 84 58 85 62
rect 77 57 85 58
rect 57 28 58 32
rect 62 28 63 32
rect 57 18 63 28
rect 77 23 83 57
rect 67 22 73 23
rect 67 18 68 22
rect 72 18 73 22
rect 3 17 9 18
rect 29 17 35 18
rect 67 13 73 18
rect 77 22 85 23
rect 77 18 80 22
rect 84 18 85 22
rect 77 17 85 18
rect -2 12 92 13
rect -2 8 16 12
rect 20 8 68 12
rect 72 8 92 12
rect -2 -1 92 8
<< ntransistor >>
rect 11 5 13 15
rect 23 5 25 15
rect 31 5 33 15
rect 47 5 49 15
rect 55 5 57 15
rect 75 5 77 25
<< ptransistor >>
rect 11 65 13 85
rect 23 65 25 85
rect 31 65 33 85
rect 47 65 49 85
rect 55 65 57 85
rect 75 55 77 95
<< polycontact >>
rect 18 58 22 62
rect 58 58 62 62
rect 48 52 52 56
rect 38 46 42 50
rect 28 38 32 42
rect 18 28 22 32
rect 30 18 34 22
rect 58 28 62 32
<< ndcontact >>
rect 4 18 8 22
rect 38 28 42 32
rect 68 18 72 22
rect 16 8 20 12
rect 68 8 72 12
rect 80 18 84 22
<< pdcontact >>
rect 16 88 20 92
rect 68 88 72 92
rect 4 78 8 82
rect 4 68 8 72
rect 38 78 42 82
rect 38 68 42 72
rect 68 78 72 82
rect 68 68 72 72
rect 68 58 72 62
rect 80 78 84 82
rect 80 68 84 72
rect 80 58 84 62
<< nsubstratencontact >>
rect 28 92 32 96
rect 38 92 42 96
rect 48 92 52 96
<< nsubstratendiff >>
rect 27 96 53 97
rect 27 92 28 96
rect 32 92 38 96
rect 42 92 48 96
rect 52 92 53 96
rect 27 91 53 92
<< labels >>
rlabel metal1 20 55 20 55 6 i0
rlabel metal1 20 55 20 55 6 i0
rlabel metal1 30 55 30 55 6 cmd
rlabel metal1 30 55 30 55 6 cmd
rlabel metal1 45 6 45 6 6 vss
rlabel metal1 45 6 45 6 6 vss
rlabel metal1 60 50 60 50 6 i1
rlabel metal1 60 50 60 50 6 i1
rlabel metal1 45 94 45 94 6 vdd
rlabel metal1 45 94 45 94 6 vdd
rlabel metal1 80 50 80 50 6 q
rlabel metal1 80 50 80 50 6 q
<< end >>
