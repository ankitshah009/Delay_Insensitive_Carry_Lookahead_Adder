magic
tech scmos
timestamp 1180640107
<< checkpaint >>
rect -24 -26 84 126
<< ab >>
rect 0 0 60 100
<< pwell >>
rect -4 -6 64 49
<< nwell >>
rect -4 49 64 106
<< polysilicon >>
rect 23 94 25 98
rect 31 94 33 98
rect 39 94 41 98
rect 47 94 49 98
rect 23 52 25 55
rect 19 51 25 52
rect 19 48 20 51
rect 11 47 20 48
rect 24 47 25 51
rect 11 46 25 47
rect 11 23 13 46
rect 31 43 33 55
rect 29 42 35 43
rect 29 39 30 42
rect 23 38 30 39
rect 34 38 35 42
rect 23 37 35 38
rect 23 23 25 37
rect 39 33 41 55
rect 47 52 49 55
rect 47 51 53 52
rect 47 47 48 51
rect 52 47 53 51
rect 47 46 53 47
rect 35 32 43 33
rect 35 28 38 32
rect 42 28 43 32
rect 35 27 43 28
rect 35 23 37 27
rect 47 23 49 46
rect 11 12 13 17
rect 23 12 25 17
rect 35 12 37 17
rect 47 12 49 17
<< ndiffusion >>
rect 3 17 11 23
rect 13 22 23 23
rect 13 18 16 22
rect 20 18 23 22
rect 13 17 23 18
rect 25 17 35 23
rect 37 22 47 23
rect 37 18 40 22
rect 44 18 47 22
rect 37 17 47 18
rect 49 22 57 23
rect 49 18 52 22
rect 56 18 57 22
rect 49 17 57 18
rect 3 12 9 17
rect 27 12 33 17
rect 3 8 4 12
rect 8 8 9 12
rect 3 7 9 8
rect 27 8 28 12
rect 32 8 33 12
rect 27 7 33 8
<< pdiffusion >>
rect 18 73 23 94
rect 15 72 23 73
rect 15 68 16 72
rect 20 68 23 72
rect 15 62 23 68
rect 15 58 16 62
rect 20 58 23 62
rect 15 57 23 58
rect 18 55 23 57
rect 25 55 31 94
rect 33 55 39 94
rect 41 55 47 94
rect 49 92 57 94
rect 49 88 52 92
rect 56 88 57 92
rect 49 82 57 88
rect 49 78 52 82
rect 56 78 57 82
rect 49 55 57 78
<< metal1 >>
rect -2 92 62 100
rect -2 88 52 92
rect 56 88 62 92
rect 52 82 56 88
rect 52 77 56 78
rect 16 72 22 73
rect 20 68 22 72
rect 37 68 53 72
rect 16 63 22 68
rect 8 62 22 63
rect 8 58 16 62
rect 20 58 22 62
rect 8 57 22 58
rect 8 22 12 57
rect 28 53 32 63
rect 18 51 32 53
rect 18 47 20 51
rect 24 47 32 51
rect 18 37 22 47
rect 38 43 42 53
rect 47 51 53 68
rect 47 47 48 51
rect 52 47 53 51
rect 28 42 42 43
rect 28 38 30 42
rect 34 38 42 42
rect 28 37 42 38
rect 28 27 32 37
rect 48 32 52 43
rect 37 28 38 32
rect 42 28 52 32
rect 37 27 52 28
rect 52 22 56 23
rect 8 18 16 22
rect 20 18 40 22
rect 44 18 45 22
rect 8 17 45 18
rect 52 12 56 18
rect -2 8 4 12
rect 8 8 28 12
rect 32 8 62 12
rect -2 0 62 8
<< ntransistor >>
rect 11 17 13 23
rect 23 17 25 23
rect 35 17 37 23
rect 47 17 49 23
<< ptransistor >>
rect 23 55 25 94
rect 31 55 33 94
rect 39 55 41 94
rect 47 55 49 94
<< polycontact >>
rect 20 47 24 51
rect 30 38 34 42
rect 48 47 52 51
rect 38 28 42 32
<< ndcontact >>
rect 16 18 20 22
rect 40 18 44 22
rect 52 18 56 22
rect 4 8 8 12
rect 28 8 32 12
<< pdcontact >>
rect 16 68 20 72
rect 16 58 20 62
rect 52 88 56 92
rect 52 78 56 82
<< psubstratepcontact >>
rect 40 4 44 8
rect 50 4 54 8
<< nsubstratencontact >>
rect 4 92 8 96
<< psubstratepdiff >>
rect 39 8 55 9
rect 39 4 40 8
rect 44 4 50 8
rect 54 4 55 8
rect 39 3 55 4
<< nsubstratendiff >>
rect 3 96 9 97
rect 3 92 4 96
rect 8 92 9 96
rect 3 91 9 92
<< labels >>
rlabel metal1 20 20 20 20 6 z
rlabel metal1 20 20 20 20 6 z
rlabel metal1 10 40 10 40 6 z
rlabel metal1 10 40 10 40 6 z
rlabel metal1 20 45 20 45 6 d
rlabel metal1 20 45 20 45 6 d
rlabel metal1 20 65 20 65 6 z
rlabel metal1 20 65 20 65 6 z
rlabel metal1 30 6 30 6 6 vss
rlabel metal1 30 6 30 6 6 vss
rlabel metal1 30 20 30 20 6 z
rlabel metal1 30 20 30 20 6 z
rlabel metal1 30 35 30 35 6 c
rlabel metal1 30 35 30 35 6 c
rlabel metal1 30 55 30 55 6 d
rlabel metal1 30 55 30 55 6 d
rlabel metal1 30 94 30 94 6 vdd
rlabel metal1 30 94 30 94 6 vdd
rlabel metal1 40 20 40 20 6 z
rlabel metal1 40 20 40 20 6 z
rlabel polycontact 40 30 40 30 6 b
rlabel polycontact 40 30 40 30 6 b
rlabel metal1 40 45 40 45 6 c
rlabel metal1 40 45 40 45 6 c
rlabel metal1 40 70 40 70 6 a
rlabel metal1 40 70 40 70 6 a
rlabel metal1 50 35 50 35 6 b
rlabel metal1 50 35 50 35 6 b
rlabel metal1 50 60 50 60 6 a
rlabel metal1 50 60 50 60 6 a
<< end >>
