magic
tech scmos
timestamp 1179385078
<< checkpaint >>
rect -22 -22 78 94
<< ab >>
rect 0 0 56 72
<< pwell >>
rect -4 -4 60 32
<< nwell >>
rect -4 32 60 76
<< polysilicon >>
rect 9 66 11 70
rect 19 63 21 68
rect 29 63 31 68
rect 41 63 43 68
rect 9 35 11 38
rect 19 35 21 46
rect 29 43 31 46
rect 29 42 35 43
rect 29 38 30 42
rect 34 38 35 42
rect 29 37 35 38
rect 9 34 15 35
rect 9 30 10 34
rect 14 30 15 34
rect 9 29 15 30
rect 19 34 25 35
rect 19 30 20 34
rect 24 30 25 34
rect 19 29 25 30
rect 9 25 11 29
rect 22 25 24 29
rect 29 25 31 37
rect 41 35 43 46
rect 41 34 47 35
rect 41 31 42 34
rect 36 30 42 31
rect 46 30 47 34
rect 36 29 47 30
rect 36 25 38 29
rect 9 6 11 11
rect 22 3 24 8
rect 29 3 31 8
rect 36 3 38 8
<< ndiffusion >>
rect 4 19 9 25
rect 2 18 9 19
rect 2 14 3 18
rect 7 14 9 18
rect 2 13 9 14
rect 4 11 9 13
rect 11 11 22 25
rect 13 8 22 11
rect 24 8 29 25
rect 31 8 36 25
rect 38 18 43 25
rect 38 17 45 18
rect 38 13 40 17
rect 44 13 45 17
rect 38 12 45 13
rect 38 8 43 12
rect 13 4 15 8
rect 19 4 20 8
rect 13 3 20 4
<< pdiffusion >>
rect 33 68 39 69
rect 4 51 9 66
rect 2 50 9 51
rect 2 46 3 50
rect 7 46 9 50
rect 2 43 9 46
rect 2 39 3 43
rect 7 39 9 43
rect 2 38 9 39
rect 11 63 17 66
rect 33 64 34 68
rect 38 64 39 68
rect 33 63 39 64
rect 11 62 19 63
rect 11 58 13 62
rect 17 58 19 62
rect 11 46 19 58
rect 21 58 29 63
rect 21 54 23 58
rect 27 54 29 58
rect 21 51 29 54
rect 21 47 23 51
rect 27 47 29 51
rect 21 46 29 47
rect 31 46 41 63
rect 43 60 48 63
rect 43 59 50 60
rect 43 55 45 59
rect 49 55 50 59
rect 43 54 50 55
rect 43 46 48 54
rect 11 38 17 46
<< metal1 >>
rect -2 68 58 72
rect -2 64 34 68
rect 38 64 58 68
rect 13 62 17 64
rect 13 57 17 58
rect 23 58 45 59
rect 27 55 45 58
rect 49 55 50 59
rect 27 54 28 55
rect 23 51 28 54
rect 2 50 7 51
rect 2 46 3 50
rect 2 43 7 46
rect 2 39 3 43
rect 2 38 7 39
rect 10 47 23 51
rect 27 47 28 51
rect 2 18 6 38
rect 10 34 14 47
rect 18 34 22 43
rect 42 42 46 51
rect 29 38 30 42
rect 34 38 46 42
rect 18 30 20 34
rect 24 30 31 34
rect 41 30 42 34
rect 46 30 47 34
rect 10 26 14 30
rect 41 26 47 30
rect 10 22 26 26
rect 33 22 47 26
rect 2 14 3 18
rect 7 14 15 18
rect 2 13 15 14
rect 22 17 26 22
rect 22 13 40 17
rect 44 13 45 17
rect -2 4 15 8
rect 19 4 58 8
rect -2 0 58 4
<< ntransistor >>
rect 9 11 11 25
rect 22 8 24 25
rect 29 8 31 25
rect 36 8 38 25
<< ptransistor >>
rect 9 38 11 66
rect 19 46 21 63
rect 29 46 31 63
rect 41 46 43 63
<< polycontact >>
rect 30 38 34 42
rect 10 30 14 34
rect 20 30 24 34
rect 42 30 46 34
<< ndcontact >>
rect 3 14 7 18
rect 40 13 44 17
rect 15 4 19 8
<< pdcontact >>
rect 3 46 7 50
rect 3 39 7 43
rect 34 64 38 68
rect 13 58 17 62
rect 23 54 27 58
rect 23 47 27 51
rect 45 55 49 59
<< labels >>
rlabel polycontact 12 32 12 32 6 zn
rlabel metal1 4 32 4 32 6 z
rlabel metal1 12 16 12 16 6 z
rlabel metal1 20 40 20 40 6 a
rlabel metal1 12 36 12 36 6 zn
rlabel metal1 28 4 28 4 6 vss
rlabel metal1 28 32 28 32 6 a
rlabel metal1 36 24 36 24 6 c
rlabel metal1 36 40 36 40 6 b
rlabel metal1 19 49 19 49 6 zn
rlabel metal1 25 53 25 53 6 zn
rlabel metal1 28 68 28 68 6 vdd
rlabel metal1 33 15 33 15 6 zn
rlabel metal1 44 28 44 28 6 c
rlabel metal1 44 48 44 48 6 b
rlabel metal1 36 57 36 57 6 zn
<< end >>
