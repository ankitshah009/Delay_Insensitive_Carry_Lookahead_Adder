magic
tech scmos
timestamp 1180640099
<< checkpaint >>
rect -24 -26 84 126
<< ab >>
rect 0 0 60 100
<< pwell >>
rect -4 -6 64 49
<< nwell >>
rect -4 49 64 106
<< polysilicon >>
rect 15 94 17 98
rect 23 94 25 98
rect 35 94 37 98
rect 43 94 45 98
rect 15 43 17 55
rect 23 52 25 55
rect 35 52 37 55
rect 23 51 37 52
rect 23 50 28 51
rect 27 47 28 50
rect 32 50 37 51
rect 32 47 33 50
rect 27 46 33 47
rect 15 42 23 43
rect 15 38 18 42
rect 22 38 23 42
rect 15 37 23 38
rect 15 34 17 37
rect 27 34 29 46
rect 43 43 45 55
rect 37 42 45 43
rect 37 38 38 42
rect 42 38 45 42
rect 37 37 45 38
rect 15 8 17 13
rect 27 8 29 13
<< ndiffusion >>
rect 6 22 15 34
rect 6 18 8 22
rect 12 18 15 22
rect 6 13 15 18
rect 17 32 27 34
rect 17 28 20 32
rect 24 28 27 32
rect 17 22 27 28
rect 17 18 20 22
rect 24 18 27 22
rect 17 13 27 18
rect 29 32 38 34
rect 29 28 32 32
rect 36 28 38 32
rect 29 22 38 28
rect 29 18 32 22
rect 36 18 38 22
rect 29 13 38 18
<< pdiffusion >>
rect 6 92 15 94
rect 6 88 8 92
rect 12 88 15 92
rect 6 82 15 88
rect 6 78 8 82
rect 12 78 15 82
rect 6 72 15 78
rect 6 68 8 72
rect 12 68 15 72
rect 6 55 15 68
rect 17 55 23 94
rect 25 72 35 94
rect 25 68 28 72
rect 32 68 35 72
rect 25 62 35 68
rect 25 58 28 62
rect 32 58 35 62
rect 25 55 35 58
rect 37 55 43 94
rect 45 92 54 94
rect 45 88 48 92
rect 52 88 54 92
rect 45 82 54 88
rect 45 78 48 82
rect 52 78 54 82
rect 45 72 54 78
rect 45 68 48 72
rect 52 68 54 72
rect 45 55 54 68
<< metal1 >>
rect -2 92 62 100
rect -2 88 8 92
rect 12 88 48 92
rect 52 88 62 92
rect 8 82 12 88
rect 8 72 12 78
rect 48 82 52 88
rect 48 72 52 78
rect 8 67 12 68
rect 27 68 28 72
rect 32 68 33 72
rect 27 63 33 68
rect 48 67 52 68
rect 8 62 33 63
rect 8 58 28 62
rect 32 58 33 62
rect 8 33 12 58
rect 38 53 42 63
rect 17 42 22 53
rect 27 51 42 53
rect 27 47 28 51
rect 32 47 42 51
rect 17 38 18 42
rect 22 38 38 42
rect 42 38 43 42
rect 8 32 24 33
rect 8 28 20 32
rect 8 27 24 28
rect 8 22 12 23
rect 8 12 12 18
rect 18 22 24 27
rect 18 18 20 22
rect 18 17 24 18
rect 32 32 36 33
rect 32 22 36 28
rect 32 12 36 18
rect -2 0 62 12
<< ntransistor >>
rect 15 13 17 34
rect 27 13 29 34
<< ptransistor >>
rect 15 55 17 94
rect 23 55 25 94
rect 35 55 37 94
rect 43 55 45 94
<< polycontact >>
rect 28 47 32 51
rect 18 38 22 42
rect 38 38 42 42
<< ndcontact >>
rect 8 18 12 22
rect 20 28 24 32
rect 20 18 24 22
rect 32 28 36 32
rect 32 18 36 22
<< pdcontact >>
rect 8 88 12 92
rect 8 78 12 82
rect 8 68 12 72
rect 28 68 32 72
rect 28 58 32 62
rect 48 88 52 92
rect 48 78 52 82
rect 48 68 52 72
<< psubstratepcontact >>
rect 48 4 52 8
<< psubstratepdiff >>
rect 47 8 53 37
rect 47 4 48 8
rect 52 4 53 8
rect 47 3 53 4
<< labels >>
rlabel metal1 10 45 10 45 6 z
rlabel metal1 10 45 10 45 6 z
rlabel metal1 20 25 20 25 6 z
rlabel metal1 20 25 20 25 6 z
rlabel metal1 20 45 20 45 6 a
rlabel metal1 20 45 20 45 6 a
rlabel metal1 20 60 20 60 6 z
rlabel metal1 20 60 20 60 6 z
rlabel metal1 30 6 30 6 6 vss
rlabel metal1 30 6 30 6 6 vss
rlabel metal1 30 40 30 40 6 a
rlabel metal1 30 40 30 40 6 a
rlabel polycontact 40 40 40 40 6 a
rlabel polycontact 40 40 40 40 6 a
rlabel polycontact 30 50 30 50 6 b
rlabel polycontact 30 50 30 50 6 b
rlabel metal1 30 65 30 65 6 z
rlabel metal1 30 65 30 65 6 z
rlabel metal1 40 55 40 55 6 b
rlabel metal1 40 55 40 55 6 b
rlabel metal1 30 94 30 94 6 vdd
rlabel metal1 30 94 30 94 6 vdd
<< end >>
