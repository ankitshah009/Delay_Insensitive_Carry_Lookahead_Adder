magic
tech scmos
timestamp 1180640144
<< checkpaint >>
rect -22 -22 92 122
<< ab >>
rect 0 0 70 100
<< metal1 >>
rect -2 98 38 102
rect 42 98 48 102
rect 52 98 58 102
rect 62 98 72 102
rect -2 92 72 98
rect -2 88 38 92
rect 42 88 48 92
rect 52 88 58 92
rect 62 88 72 92
rect -2 8 8 12
rect 12 8 18 12
rect 22 8 28 12
rect 32 8 72 12
rect -2 2 72 8
rect -2 -2 8 2
rect 12 -2 18 2
rect 22 -2 28 2
rect 32 -2 72 2
<< metal2 >>
rect 7 98 8 102
rect 12 98 18 102
rect 22 98 28 102
rect 32 98 38 102
rect 42 98 48 102
rect 52 98 58 102
rect 62 98 63 102
rect 7 92 63 98
rect 7 88 8 92
rect 12 88 18 92
rect 22 88 28 92
rect 32 88 38 92
rect 42 88 48 92
rect 52 88 58 92
rect 62 88 63 92
rect 7 8 8 12
rect 12 8 18 12
rect 22 8 28 12
rect 32 8 38 12
rect 42 8 48 12
rect 52 8 58 12
rect 62 8 63 12
rect 7 2 63 8
rect 7 -2 8 2
rect 12 -2 18 2
rect 22 -2 28 2
rect 32 -2 38 2
rect 42 -2 48 2
rect 52 -2 58 2
rect 62 -2 63 2
<< metal3 >>
rect 7 98 8 102
rect 12 98 18 102
rect 22 98 28 102
rect 32 98 33 102
rect 7 92 33 98
rect 7 88 8 92
rect 12 88 18 92
rect 22 88 28 92
rect 32 88 33 92
rect 7 -2 33 88
rect 37 12 63 102
rect 37 8 38 12
rect 42 8 48 12
rect 52 8 58 12
rect 62 8 63 12
rect 37 2 63 8
rect 37 -2 38 2
rect 42 -2 48 2
rect 52 -2 58 2
rect 62 -2 63 2
<< m2contact >>
rect 38 98 42 102
rect 48 98 52 102
rect 58 98 62 102
rect 38 88 42 92
rect 48 88 52 92
rect 58 88 62 92
rect 8 8 12 12
rect 18 8 22 12
rect 28 8 32 12
rect 8 -2 12 2
rect 18 -2 22 2
rect 28 -2 32 2
<< m3contact >>
rect 8 98 12 102
rect 18 98 22 102
rect 28 98 32 102
rect 8 88 12 92
rect 18 88 22 92
rect 28 88 32 92
rect 38 8 42 12
rect 48 8 52 12
rect 58 8 62 12
rect 38 -2 42 2
rect 48 -2 52 2
rect 58 -2 62 2
<< labels >>
rlabel metal1 35 6 35 6 6 vss
rlabel metal1 35 6 35 6 6 vss
rlabel metal1 35 94 35 94 6 vdd
rlabel metal1 35 94 35 94 6 vdd
rlabel metal2 35 6 35 6 6 vss
rlabel metal2 35 94 35 94 6 vdd
<< end >>
