magic
tech scmos
timestamp 1180600712
<< checkpaint >>
rect -22 -22 62 122
<< ab >>
rect 0 0 40 100
<< pwell >>
rect -4 -4 44 48
<< nwell >>
rect -4 48 44 104
<< polysilicon >>
rect 19 94 21 98
rect 27 94 29 98
rect 19 53 21 56
rect 17 52 23 53
rect 17 49 18 52
rect 13 48 18 49
rect 22 48 23 52
rect 13 47 23 48
rect 13 25 15 47
rect 27 43 29 56
rect 27 42 33 43
rect 27 41 28 42
rect 25 38 28 41
rect 32 38 33 42
rect 25 37 33 38
rect 25 25 27 37
rect 13 11 15 15
rect 25 11 27 15
<< ndiffusion >>
rect 5 15 13 25
rect 15 22 25 25
rect 15 18 18 22
rect 22 18 25 22
rect 15 15 25 18
rect 27 15 35 25
rect 5 12 11 15
rect 5 8 6 12
rect 10 8 11 12
rect 29 12 35 15
rect 5 7 11 8
rect 29 8 30 12
rect 34 8 35 12
rect 29 7 35 8
<< pdiffusion >>
rect 14 85 19 94
rect 7 82 19 85
rect 7 78 8 82
rect 12 78 19 82
rect 7 72 19 78
rect 7 68 8 72
rect 12 68 19 72
rect 7 62 19 68
rect 7 58 8 62
rect 12 58 19 62
rect 7 56 19 58
rect 21 56 27 94
rect 29 92 37 94
rect 29 88 32 92
rect 36 88 37 92
rect 29 56 37 88
rect 7 55 13 56
<< metal1 >>
rect -2 92 42 100
rect -2 88 32 92
rect 36 88 42 92
rect 8 82 12 83
rect 8 72 12 78
rect 8 62 12 68
rect 8 22 12 58
rect 18 52 22 83
rect 18 27 22 48
rect 28 42 32 83
rect 8 18 18 22
rect 22 18 23 22
rect 8 17 12 18
rect 28 17 32 38
rect -2 8 6 12
rect 10 8 30 12
rect 34 8 42 12
rect -2 0 42 8
<< ntransistor >>
rect 13 15 15 25
rect 25 15 27 25
<< ptransistor >>
rect 19 56 21 94
rect 27 56 29 94
<< polycontact >>
rect 18 48 22 52
rect 28 38 32 42
<< ndcontact >>
rect 18 18 22 22
rect 6 8 10 12
rect 30 8 34 12
<< pdcontact >>
rect 8 78 12 82
rect 8 68 12 72
rect 8 58 12 62
rect 32 88 36 92
<< labels >>
rlabel metal1 10 50 10 50 6 nq
rlabel ndcontact 20 20 20 20 6 nq
rlabel metal1 20 6 20 6 6 vss
rlabel metal1 20 55 20 55 6 i1
rlabel metal1 20 94 20 94 6 vdd
rlabel metal1 30 50 30 50 6 i0
<< end >>
