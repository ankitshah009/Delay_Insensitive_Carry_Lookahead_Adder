.subckt nmx3_x1 cmd0 cmd1 i0 i1 i2 nq vdd vss
*   SPICE3 file   created from nmx3_x1.ext -      technology: scmos
m00 w1     i2     w2     vdd p w=20u  l=2.3636u ad=100p     pd=30u      as=120p     ps=38.6667u
m01 nq     cmd1   w1     vdd p w=20u  l=2.3636u ad=136p     pd=44u      as=100p     ps=30u
m02 w3     w4     nq     vdd p w=20u  l=2.3636u ad=60p      pd=26u      as=136p     ps=44u
m03 w2     i1     w3     vdd p w=20u  l=2.3636u ad=120p     pd=38.6667u as=60p      ps=26u
m04 vdd    w5     w2     vdd p w=20u  l=2.3636u ad=174.118p pd=60u      as=120p     ps=38.6667u
m05 w6     cmd0   vdd    vdd p w=20u  l=2.3636u ad=60p      pd=26u      as=174.118p ps=60u
m06 nq     i0     w6     vdd p w=20u  l=2.3636u ad=136p     pd=44u      as=60p      ps=26u
m07 w4     cmd1   vdd    vdd p w=14u  l=2.3636u ad=112p     pd=44u      as=121.882p ps=42u
m08 w4     cmd1   vss    vss n w=8u   l=2.3636u ad=64p      pd=32u      as=90.4p    ps=35.2u
m09 vdd    cmd0   w5     vdd p w=14u  l=2.3636u ad=121.882p pd=42u      as=112p     ps=44u
m10 w7     i2     w8     vss n w=12u  l=2.3636u ad=60p      pd=22u      as=80p      ps=30.6667u
m11 nq     w4     w7     vss n w=12u  l=2.3636u ad=100p     pd=37.3333u as=60p      ps=22u
m12 w9     cmd1   nq     vss n w=12u  l=2.3636u ad=36p      pd=18u      as=100p     ps=37.3333u
m13 w8     i1     w9     vss n w=12u  l=2.3636u ad=80p      pd=30.6667u as=36p      ps=18u
m14 vss    cmd0   w5     vss n w=8u   l=2.3636u ad=90.4p    pd=35.2u    as=64p      ps=32u
m15 vss    cmd0   w8     vss n w=12u  l=2.3636u ad=135.6p   pd=52.8u    as=80p      ps=30.6667u
m16 w10    w5     vss    vss n w=12u  l=2.3636u ad=36p      pd=18u      as=135.6p   ps=52.8u
m17 nq     i0     w10    vss n w=12u  l=2.3636u ad=100p     pd=37.3333u as=36p      ps=18u
C0  w1     vdd    0.023f
C1  nq     i0     0.209f
C2  w8     w4     0.184f
C3  vss    i1     0.017f
C4  w5     cmd1   0.044f
C5  cmd0   i2     0.014f
C6  i1     w4     0.224f
C7  w8     i2     0.017f
C8  nq     w5     0.466f
C9  vss    cmd1   0.059f
C10 w4     cmd1   0.577f
C11 i1     i2     0.075f
C12 vss    nq     0.225f
C13 vdd    cmd0   0.019f
C14 nq     w4     0.222f
C15 cmd1   i2     0.187f
C16 w2     w4     0.081f
C17 i0     w5     0.369f
C18 nq     i2     0.021f
C19 vdd    i1     0.018f
C20 w10    vss    0.011f
C21 w9     w8     0.011f
C22 w8     cmd0   0.004f
C23 w3     w2     0.014f
C24 w6     vdd    0.014f
C25 vss    i0     0.022f
C26 cmd0   i1     0.080f
C27 i0     w4     0.017f
C28 vdd    cmd1   0.142f
C29 w2     i2     0.013f
C30 w7     vss    0.010f
C31 w8     i1     0.025f
C32 w1     w2     0.024f
C33 nq     vdd    0.324f
C34 vss    w5     0.087f
C35 cmd0   cmd1   0.030f
C36 w5     w4     0.041f
C37 w2     vdd    0.457f
C38 w8     cmd1   0.006f
C39 nq     cmd0   0.269f
C40 vss    w4     0.051f
C41 i1     cmd1   0.152f
C42 w5     i2     0.022f
C43 w8     nq     0.105f
C44 nq     i1     0.159f
C45 vdd    i0     0.022f
C46 vss    i2     0.010f
C47 w2     cmd0   0.004f
C48 w4     i2     0.236f
C49 i0     cmd0   0.361f
C50 nq     cmd1   0.068f
C51 vdd    w5     0.015f
C52 w2     i1     0.025f
C53 i0     i1     0.030f
C54 cmd0   w5     0.361f
C55 vdd    w4     0.050f
C56 w2     cmd1   0.157f
C57 w9     vss    0.006f
C58 w7     w8     0.019f
C59 nq     w2     0.241f
C60 w3     vdd    0.014f
C61 w8     w5     0.030f
C62 vss    cmd0   0.019f
C63 i0     cmd1   0.008f
C64 vdd    i2     0.010f
C65 cmd0   w4     0.029f
C66 w5     i1     0.128f
C67 w8     vss    0.434f
C69 nq     vss    0.073f
C71 i0     vss    0.052f
C72 cmd0   vss    0.069f
C73 w5     vss    0.063f
C74 i1     vss    0.040f
C75 w4     vss    0.059f
C76 cmd1   vss    0.076f
C77 i2     vss    0.033f
.ends
