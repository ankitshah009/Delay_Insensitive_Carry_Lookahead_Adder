magic
tech scmos
timestamp 1185094809
<< checkpaint >>
rect -20 -20 90 120
<< metal1 >>
rect -2 98 72 102
rect -2 94 38 98
rect 42 94 46 98
rect 50 94 54 98
rect 58 94 72 98
rect -2 88 72 94
rect -2 10 72 12
rect -2 6 14 10
rect 18 6 22 10
rect 26 6 72 10
rect -2 2 72 6
rect -2 -2 14 2
rect 18 -2 22 2
rect 26 -2 72 2
<< metal2 >>
rect 7 98 63 102
rect 7 94 14 98
rect 18 94 22 98
rect 26 94 38 98
rect 42 94 46 98
rect 50 94 54 98
rect 58 94 63 98
rect 7 88 63 94
rect 7 10 63 12
rect 7 6 14 10
rect 18 6 22 10
rect 26 6 38 10
rect 42 6 46 10
rect 50 6 54 10
rect 58 6 63 10
rect 7 2 63 6
rect 7 -2 14 2
rect 18 -2 22 2
rect 26 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 63 2
<< metal3 >>
rect 7 98 33 102
rect 7 94 14 98
rect 18 94 22 98
rect 26 94 33 98
rect 7 -2 33 94
rect 37 10 63 102
rect 37 6 38 10
rect 42 6 46 10
rect 50 6 54 10
rect 58 6 63 10
rect 37 2 63 6
rect 37 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 63 2
<< m2contact >>
rect 38 94 42 98
rect 46 94 50 98
rect 54 94 58 98
rect 14 6 18 10
rect 22 6 26 10
rect 14 -2 18 2
rect 22 -2 26 2
<< m3contact >>
rect 14 94 18 98
rect 22 94 26 98
rect 38 6 42 10
rect 46 6 50 10
rect 54 6 58 10
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
<< labels >>
rlabel metal1 35 6 35 6 6 vss
rlabel metal1 35 94 35 94 6 vdd
rlabel metal2 35 6 35 6 6 vss
rlabel metal2 35 94 35 94 6 vdd
<< end >>
