magic
tech scmos
timestamp 1185039152
<< checkpaint >>
rect -22 -24 262 124
<< ab >>
rect 0 0 240 100
<< pwell >>
rect -2 -4 242 49
<< nwell >>
rect -2 49 242 104
<< polysilicon >>
rect 119 95 121 98
rect 155 95 157 98
rect 167 95 169 98
rect 179 95 181 98
rect 191 95 193 98
rect 203 95 205 98
rect 215 95 217 98
rect 227 95 229 98
rect 11 85 13 88
rect 23 85 25 88
rect 31 85 33 88
rect 49 85 51 88
rect 57 85 59 88
rect 83 85 85 88
rect 95 85 97 88
rect 131 85 133 88
rect 143 85 145 88
rect 119 73 121 75
rect 115 72 121 73
rect 115 68 116 72
rect 120 68 121 72
rect 115 67 121 68
rect 155 73 157 75
rect 155 72 163 73
rect 155 68 158 72
rect 162 68 163 72
rect 155 67 163 68
rect 11 51 13 65
rect 23 63 25 65
rect 17 62 25 63
rect 17 58 18 62
rect 22 58 25 62
rect 17 57 25 58
rect 31 53 33 65
rect 49 63 51 65
rect 57 63 59 65
rect 83 63 85 65
rect 47 62 53 63
rect 47 58 48 62
rect 52 58 53 62
rect 47 57 53 58
rect 57 62 63 63
rect 57 58 58 62
rect 62 58 63 62
rect 57 57 63 58
rect 83 62 91 63
rect 83 58 86 62
rect 90 58 91 62
rect 83 57 91 58
rect 27 52 33 53
rect 27 51 28 52
rect 11 49 28 51
rect 11 25 13 49
rect 27 48 28 49
rect 32 51 33 52
rect 77 52 83 53
rect 32 49 51 51
rect 32 48 33 49
rect 27 47 33 48
rect 27 42 33 43
rect 27 38 28 42
rect 32 38 33 42
rect 27 37 33 38
rect 17 32 25 33
rect 17 28 18 32
rect 22 28 25 32
rect 17 27 25 28
rect 23 25 25 27
rect 31 25 33 37
rect 49 25 51 49
rect 77 48 78 52
rect 82 51 83 52
rect 95 51 97 65
rect 131 63 133 65
rect 127 62 133 63
rect 127 58 128 62
rect 132 58 133 62
rect 127 57 133 58
rect 127 52 133 53
rect 127 51 128 52
rect 82 49 128 51
rect 82 48 83 49
rect 77 47 83 48
rect 57 32 63 33
rect 57 28 58 32
rect 62 28 63 32
rect 57 27 63 28
rect 83 32 91 33
rect 83 28 86 32
rect 90 28 91 32
rect 83 27 91 28
rect 57 25 59 27
rect 83 25 85 27
rect 95 25 97 49
rect 127 48 128 49
rect 132 51 133 52
rect 143 51 145 65
rect 167 63 169 75
rect 161 62 169 63
rect 161 58 162 62
rect 166 58 169 62
rect 161 57 169 58
rect 179 51 181 75
rect 191 73 193 75
rect 185 72 193 73
rect 185 68 186 72
rect 190 68 193 72
rect 185 67 193 68
rect 203 53 205 75
rect 203 52 211 53
rect 132 49 193 51
rect 132 48 133 49
rect 127 47 133 48
rect 101 42 107 43
rect 101 38 102 42
rect 106 41 107 42
rect 137 42 145 43
rect 137 41 138 42
rect 106 39 138 41
rect 106 38 107 39
rect 101 37 107 38
rect 137 38 138 39
rect 142 41 145 42
rect 179 42 187 43
rect 179 41 182 42
rect 142 39 182 41
rect 142 38 145 39
rect 137 37 145 38
rect 117 32 123 33
rect 117 28 118 32
rect 122 28 123 32
rect 117 27 123 28
rect 127 32 133 33
rect 127 28 128 32
rect 132 28 133 32
rect 127 27 133 28
rect 119 25 121 27
rect 131 25 133 27
rect 143 25 145 37
rect 179 38 182 39
rect 186 38 187 42
rect 179 37 187 38
rect 161 32 169 33
rect 161 28 162 32
rect 166 28 169 32
rect 161 27 169 28
rect 155 22 163 23
rect 155 18 158 22
rect 162 18 163 22
rect 155 17 163 18
rect 155 15 157 17
rect 167 15 169 27
rect 179 25 181 37
rect 191 25 193 49
rect 203 48 206 52
rect 210 48 211 52
rect 203 47 211 48
rect 215 43 217 55
rect 227 43 229 55
rect 205 42 229 43
rect 205 38 206 42
rect 210 38 229 42
rect 205 37 229 38
rect 203 32 211 33
rect 203 28 206 32
rect 210 28 211 32
rect 203 27 211 28
rect 203 25 205 27
rect 215 25 217 37
rect 227 25 229 37
rect 11 12 13 15
rect 23 12 25 15
rect 31 12 33 15
rect 49 12 51 15
rect 57 12 59 15
rect 83 12 85 15
rect 95 12 97 15
rect 119 12 121 15
rect 131 12 133 15
rect 143 12 145 15
rect 179 12 181 15
rect 191 12 193 15
rect 203 12 205 15
rect 155 2 157 5
rect 167 2 169 5
rect 215 2 217 5
rect 227 2 229 5
<< ndiffusion >>
rect 37 32 47 33
rect 37 28 38 32
rect 42 28 47 32
rect 37 25 47 28
rect 3 22 11 25
rect 3 18 4 22
rect 8 18 11 22
rect 3 15 11 18
rect 13 15 23 25
rect 25 15 31 25
rect 33 15 49 25
rect 51 15 57 25
rect 59 15 67 25
rect 75 22 83 25
rect 75 18 76 22
rect 80 18 83 22
rect 75 15 83 18
rect 85 15 95 25
rect 97 22 105 25
rect 97 18 100 22
rect 104 18 105 22
rect 97 15 105 18
rect 111 15 119 25
rect 121 15 131 25
rect 133 22 143 25
rect 133 18 136 22
rect 140 18 143 22
rect 133 15 143 18
rect 145 15 153 25
rect 171 22 179 25
rect 171 18 172 22
rect 176 18 179 22
rect 171 15 179 18
rect 181 22 191 25
rect 181 18 184 22
rect 188 18 191 22
rect 181 15 191 18
rect 193 15 203 25
rect 205 22 215 25
rect 205 18 208 22
rect 212 18 215 22
rect 205 15 215 18
rect 15 12 21 15
rect 61 12 67 15
rect 87 12 93 15
rect 111 12 117 15
rect 15 8 16 12
rect 20 8 21 12
rect 15 7 21 8
rect 61 8 62 12
rect 66 8 67 12
rect 61 7 67 8
rect 87 8 88 12
rect 92 8 93 12
rect 87 7 93 8
rect 111 8 112 12
rect 116 8 117 12
rect 111 7 117 8
rect 147 5 155 15
rect 157 12 167 15
rect 157 8 160 12
rect 164 8 167 12
rect 157 5 167 8
rect 169 5 177 15
rect 207 12 215 15
rect 207 8 208 12
rect 212 8 215 12
rect 207 5 215 8
rect 217 22 227 25
rect 217 18 220 22
rect 224 18 227 22
rect 217 5 227 18
rect 229 22 237 25
rect 229 18 232 22
rect 236 18 237 22
rect 229 12 237 18
rect 229 8 232 12
rect 236 8 237 12
rect 229 5 237 8
<< pdiffusion >>
rect 15 92 21 93
rect 15 88 16 92
rect 20 88 21 92
rect 61 92 67 93
rect 61 88 62 92
rect 66 88 67 92
rect 87 92 93 93
rect 87 88 88 92
rect 92 88 93 92
rect 111 92 119 95
rect 111 88 112 92
rect 116 88 119 92
rect 15 85 21 88
rect 61 85 67 88
rect 87 85 93 88
rect 3 72 11 85
rect 3 68 4 72
rect 8 68 11 72
rect 3 65 11 68
rect 13 65 23 85
rect 25 65 31 85
rect 33 72 49 85
rect 33 68 38 72
rect 42 68 49 72
rect 33 65 49 68
rect 51 65 57 85
rect 59 65 67 85
rect 75 72 83 85
rect 75 68 76 72
rect 80 68 83 72
rect 75 65 83 68
rect 85 65 95 85
rect 97 72 105 85
rect 111 75 119 88
rect 121 85 129 95
rect 147 85 155 95
rect 121 75 131 85
rect 97 68 100 72
rect 104 68 105 72
rect 97 65 105 68
rect 123 65 131 75
rect 133 72 143 85
rect 133 68 136 72
rect 140 68 143 72
rect 133 65 143 68
rect 145 75 155 85
rect 157 92 167 95
rect 157 88 160 92
rect 164 88 167 92
rect 157 75 167 88
rect 169 82 179 95
rect 169 78 172 82
rect 176 78 179 82
rect 169 75 179 78
rect 181 82 191 95
rect 181 78 184 82
rect 188 78 191 82
rect 181 75 191 78
rect 193 75 203 95
rect 205 92 215 95
rect 205 88 208 92
rect 212 88 215 92
rect 205 82 215 88
rect 205 78 208 82
rect 212 78 215 82
rect 205 75 215 78
rect 145 65 153 75
rect 207 72 215 75
rect 207 68 208 72
rect 212 68 215 72
rect 207 62 215 68
rect 207 58 208 62
rect 212 58 215 62
rect 207 55 215 58
rect 217 82 227 95
rect 217 78 220 82
rect 224 78 227 82
rect 217 72 227 78
rect 217 68 220 72
rect 224 68 227 72
rect 217 62 227 68
rect 217 58 220 62
rect 224 58 227 62
rect 217 55 227 58
rect 229 92 237 95
rect 229 88 232 92
rect 236 88 237 92
rect 229 82 237 88
rect 229 78 232 82
rect 236 78 237 82
rect 229 72 237 78
rect 229 68 232 72
rect 236 68 237 72
rect 229 62 237 68
rect 229 58 232 62
rect 236 58 237 62
rect 229 55 237 58
<< metal1 >>
rect -2 96 242 101
rect -2 92 28 96
rect 32 92 48 96
rect 52 92 242 96
rect -2 88 16 92
rect 20 88 62 92
rect 66 88 88 92
rect 92 88 112 92
rect 116 88 160 92
rect 164 88 208 92
rect 212 88 232 92
rect 236 88 242 92
rect -2 87 242 88
rect 171 82 177 83
rect 3 72 9 73
rect 3 68 4 72
rect 8 68 9 72
rect 3 67 9 68
rect 4 23 8 67
rect 17 62 23 82
rect 17 58 18 62
rect 22 58 23 62
rect 17 32 23 58
rect 27 52 33 82
rect 38 78 122 82
rect 38 73 42 78
rect 118 73 122 78
rect 171 78 172 82
rect 176 78 177 82
rect 171 77 177 78
rect 183 82 189 83
rect 207 82 213 87
rect 219 82 225 83
rect 183 78 184 82
rect 188 78 200 82
rect 183 77 189 78
rect 37 72 43 73
rect 75 72 81 73
rect 99 72 105 73
rect 37 68 38 72
rect 42 68 43 72
rect 37 67 43 68
rect 27 48 28 52
rect 32 48 33 52
rect 27 47 33 48
rect 27 42 33 43
rect 27 38 28 42
rect 32 38 33 42
rect 27 37 33 38
rect 17 28 18 32
rect 22 28 23 32
rect 17 27 23 28
rect 3 22 9 23
rect 28 22 32 37
rect 38 33 42 67
rect 47 62 53 63
rect 47 58 48 62
rect 52 58 53 62
rect 47 57 53 58
rect 57 62 63 72
rect 75 68 76 72
rect 80 68 81 72
rect 75 67 81 68
rect 57 58 58 62
rect 62 58 63 62
rect 37 32 43 33
rect 37 28 38 32
rect 42 28 43 32
rect 37 27 43 28
rect 48 22 52 57
rect 3 18 4 22
rect 8 18 52 22
rect 57 32 63 58
rect 57 28 58 32
rect 62 28 63 32
rect 57 18 63 28
rect 76 53 80 67
rect 87 63 93 72
rect 99 68 100 72
rect 104 68 105 72
rect 99 67 105 68
rect 115 72 122 73
rect 115 68 116 72
rect 120 68 122 72
rect 115 67 122 68
rect 135 72 141 73
rect 157 72 163 73
rect 172 72 176 77
rect 185 72 191 73
rect 135 68 136 72
rect 140 68 152 72
rect 135 67 141 68
rect 85 62 93 63
rect 85 58 86 62
rect 90 58 93 62
rect 85 57 93 58
rect 76 52 83 53
rect 76 48 78 52
rect 82 48 83 52
rect 76 47 83 48
rect 76 23 80 47
rect 87 33 93 57
rect 85 32 93 33
rect 85 28 86 32
rect 90 28 93 32
rect 85 27 93 28
rect 75 22 81 23
rect 75 18 76 22
rect 80 18 81 22
rect 87 18 93 27
rect 100 43 104 67
rect 100 42 107 43
rect 100 38 102 42
rect 106 38 107 42
rect 100 37 107 38
rect 100 23 104 37
rect 118 33 122 67
rect 127 62 133 63
rect 148 62 152 68
rect 157 68 158 72
rect 162 68 176 72
rect 157 67 163 68
rect 161 62 167 63
rect 127 58 128 62
rect 132 58 142 62
rect 127 57 133 58
rect 127 52 133 53
rect 127 48 128 52
rect 132 48 133 52
rect 127 47 133 48
rect 128 33 132 47
rect 138 43 142 58
rect 148 58 162 62
rect 166 58 167 62
rect 137 42 143 43
rect 137 38 138 42
rect 142 38 143 42
rect 137 37 143 38
rect 117 32 123 33
rect 117 28 118 32
rect 122 28 123 32
rect 117 27 123 28
rect 127 32 133 33
rect 127 28 128 32
rect 132 28 133 32
rect 127 27 133 28
rect 148 32 152 58
rect 161 57 167 58
rect 161 32 167 33
rect 148 28 162 32
rect 166 28 167 32
rect 99 22 105 23
rect 99 18 100 22
rect 104 18 105 22
rect 3 17 9 18
rect 75 17 81 18
rect 99 17 105 18
rect 135 22 141 23
rect 148 22 152 28
rect 161 27 167 28
rect 172 23 176 68
rect 184 68 186 72
rect 190 68 191 72
rect 184 67 191 68
rect 184 43 188 67
rect 181 42 188 43
rect 181 38 182 42
rect 186 38 188 42
rect 196 42 200 78
rect 207 78 208 82
rect 212 78 213 82
rect 207 72 213 78
rect 207 68 208 72
rect 212 68 213 72
rect 207 62 213 68
rect 207 58 208 62
rect 212 58 213 62
rect 207 57 213 58
rect 217 78 220 82
rect 224 78 225 82
rect 217 77 225 78
rect 231 82 237 87
rect 231 78 232 82
rect 236 78 237 82
rect 217 73 223 77
rect 217 72 225 73
rect 217 68 220 72
rect 224 68 225 72
rect 217 67 225 68
rect 231 72 237 78
rect 231 68 232 72
rect 236 68 237 72
rect 217 63 223 67
rect 217 62 225 63
rect 217 58 220 62
rect 224 58 225 62
rect 217 57 225 58
rect 231 62 237 68
rect 231 58 232 62
rect 236 58 237 62
rect 231 57 237 58
rect 205 52 211 53
rect 217 52 223 57
rect 205 48 206 52
rect 210 48 224 52
rect 205 47 211 48
rect 205 42 211 43
rect 196 38 206 42
rect 210 38 211 42
rect 181 37 187 38
rect 135 18 136 22
rect 140 18 152 22
rect 157 22 163 23
rect 171 22 177 23
rect 157 18 158 22
rect 162 18 172 22
rect 176 18 177 22
rect 135 17 141 18
rect 157 17 163 18
rect 171 17 177 18
rect 183 22 189 23
rect 196 22 200 38
rect 205 37 211 38
rect 205 32 211 33
rect 217 32 223 48
rect 205 28 206 32
rect 210 28 224 32
rect 205 27 211 28
rect 217 23 223 28
rect 183 18 184 22
rect 188 18 200 22
rect 207 22 213 23
rect 207 18 208 22
rect 212 18 213 22
rect 217 22 225 23
rect 217 18 220 22
rect 224 18 225 22
rect 183 17 189 18
rect 207 13 213 18
rect 219 17 225 18
rect 231 22 237 23
rect 231 18 232 22
rect 236 18 237 22
rect 231 13 237 18
rect -2 12 242 13
rect -2 8 16 12
rect 20 8 62 12
rect 66 8 88 12
rect 92 8 112 12
rect 116 8 160 12
rect 164 8 208 12
rect 212 8 232 12
rect 236 8 242 12
rect -2 4 28 8
rect 32 4 48 8
rect 52 4 124 8
rect 128 4 136 8
rect 140 4 184 8
rect 188 4 196 8
rect 200 4 242 8
rect -2 -1 242 4
<< ntransistor >>
rect 11 15 13 25
rect 23 15 25 25
rect 31 15 33 25
rect 49 15 51 25
rect 57 15 59 25
rect 83 15 85 25
rect 95 15 97 25
rect 119 15 121 25
rect 131 15 133 25
rect 143 15 145 25
rect 179 15 181 25
rect 191 15 193 25
rect 203 15 205 25
rect 155 5 157 15
rect 167 5 169 15
rect 215 5 217 25
rect 227 5 229 25
<< ptransistor >>
rect 11 65 13 85
rect 23 65 25 85
rect 31 65 33 85
rect 49 65 51 85
rect 57 65 59 85
rect 83 65 85 85
rect 95 65 97 85
rect 119 75 121 95
rect 131 65 133 85
rect 143 65 145 85
rect 155 75 157 95
rect 167 75 169 95
rect 179 75 181 95
rect 191 75 193 95
rect 203 75 205 95
rect 215 55 217 95
rect 227 55 229 95
<< polycontact >>
rect 116 68 120 72
rect 158 68 162 72
rect 18 58 22 62
rect 48 58 52 62
rect 58 58 62 62
rect 86 58 90 62
rect 28 48 32 52
rect 28 38 32 42
rect 18 28 22 32
rect 78 48 82 52
rect 128 58 132 62
rect 58 28 62 32
rect 86 28 90 32
rect 128 48 132 52
rect 162 58 166 62
rect 186 68 190 72
rect 102 38 106 42
rect 138 38 142 42
rect 118 28 122 32
rect 128 28 132 32
rect 182 38 186 42
rect 162 28 166 32
rect 158 18 162 22
rect 206 48 210 52
rect 206 38 210 42
rect 206 28 210 32
<< ndcontact >>
rect 38 28 42 32
rect 4 18 8 22
rect 76 18 80 22
rect 100 18 104 22
rect 136 18 140 22
rect 172 18 176 22
rect 184 18 188 22
rect 208 18 212 22
rect 16 8 20 12
rect 62 8 66 12
rect 88 8 92 12
rect 112 8 116 12
rect 160 8 164 12
rect 208 8 212 12
rect 220 18 224 22
rect 232 18 236 22
rect 232 8 236 12
<< pdcontact >>
rect 16 88 20 92
rect 62 88 66 92
rect 88 88 92 92
rect 112 88 116 92
rect 4 68 8 72
rect 38 68 42 72
rect 76 68 80 72
rect 100 68 104 72
rect 136 68 140 72
rect 160 88 164 92
rect 172 78 176 82
rect 184 78 188 82
rect 208 88 212 92
rect 208 78 212 82
rect 208 68 212 72
rect 208 58 212 62
rect 220 78 224 82
rect 220 68 224 72
rect 220 58 224 62
rect 232 88 236 92
rect 232 78 236 82
rect 232 68 236 72
rect 232 58 236 62
<< psubstratepcontact >>
rect 28 4 32 8
rect 48 4 52 8
rect 124 4 128 8
rect 136 4 140 8
rect 184 4 188 8
rect 196 4 200 8
<< nsubstratencontact >>
rect 28 92 32 96
rect 48 92 52 96
<< psubstratepdiff >>
rect 27 8 53 9
rect 27 4 28 8
rect 32 4 48 8
rect 52 4 53 8
rect 123 8 141 9
rect 27 3 53 4
rect 123 4 124 8
rect 128 4 136 8
rect 140 4 141 8
rect 183 8 201 9
rect 123 3 141 4
rect 183 4 184 8
rect 188 4 196 8
rect 200 4 201 8
rect 183 3 201 4
<< nsubstratendiff >>
rect 27 96 53 97
rect 27 92 28 96
rect 32 92 48 96
rect 52 92 53 96
rect 27 91 53 92
<< labels >>
rlabel metal1 20 55 20 55 6 i0
rlabel metal1 20 55 20 55 6 i0
rlabel metal1 30 65 30 65 6 cmd
rlabel metal1 30 65 30 65 6 cmd
rlabel metal1 90 45 90 45 6 ck
rlabel metal1 60 45 60 45 6 i1
rlabel metal1 90 45 90 45 6 ck
rlabel metal1 60 45 60 45 6 i1
rlabel metal1 120 6 120 6 6 vss
rlabel metal1 120 6 120 6 6 vss
rlabel metal1 120 94 120 94 6 vdd
rlabel metal1 120 94 120 94 6 vdd
rlabel metal1 220 50 220 50 6 q
rlabel metal1 220 50 220 50 6 q
<< end >>
