magic
tech scmos
timestamp 1170759764
<< checkpaint >>
rect -22 -26 54 114
<< ab >>
rect 0 0 32 88
<< pwell >>
rect -4 -8 36 40
<< nwell >>
rect -4 40 36 96
<< polysilicon >>
rect 2 82 11 83
rect 2 78 6 82
rect 10 78 11 82
rect 2 77 11 78
rect 9 74 11 77
rect 21 77 30 83
rect 21 74 23 77
rect 9 43 11 46
rect 21 43 23 46
rect 2 37 14 43
rect 18 42 30 43
rect 18 38 22 42
rect 26 38 30 42
rect 18 37 30 38
rect 9 34 11 37
rect 21 34 23 37
rect 9 11 11 14
rect 2 5 11 11
rect 21 11 23 14
rect 21 5 30 11
<< ndiffusion >>
rect 2 14 9 34
rect 11 20 21 34
rect 11 16 14 20
rect 18 16 21 20
rect 11 14 21 16
rect 23 29 30 34
rect 23 25 25 29
rect 29 25 30 29
rect 23 21 30 25
rect 23 17 25 21
rect 29 17 30 21
rect 23 14 30 17
rect 13 13 19 14
rect 13 10 14 13
rect 18 10 19 13
rect 13 2 19 10
<< pdiffusion >>
rect 13 78 19 86
rect 13 75 14 78
rect 18 75 19 78
rect 13 74 19 75
rect 2 46 9 74
rect 11 72 21 74
rect 11 68 14 72
rect 18 68 21 72
rect 11 46 21 68
rect 23 71 30 74
rect 23 67 25 71
rect 29 67 30 71
rect 23 63 30 67
rect 23 59 25 63
rect 29 59 30 63
rect 23 46 30 59
<< metal1 >>
rect -2 86 2 90
rect 10 86 22 90
rect 30 86 34 90
rect 6 82 10 86
rect 6 77 10 78
rect 14 82 18 86
rect 14 72 18 75
rect 14 67 18 68
rect 22 67 25 71
rect 29 67 30 71
rect 22 63 26 67
rect 14 59 25 63
rect 29 59 30 63
rect 14 29 18 59
rect 22 42 26 55
rect 22 33 26 38
rect 14 25 25 29
rect 29 25 30 29
rect 22 21 26 25
rect 14 20 18 21
rect 22 17 25 21
rect 29 17 30 21
rect 14 13 18 16
rect 14 2 18 6
rect -2 -2 2 2
rect 10 -2 22 2
rect 30 -2 34 2
<< metal2 >>
rect -2 86 6 90
rect 10 86 22 90
rect 26 86 34 90
rect -2 82 34 86
rect -2 78 14 82
rect 18 78 34 82
rect -2 76 34 78
rect -2 10 34 12
rect -2 6 14 10
rect 18 6 34 10
rect -2 2 34 6
rect -2 -2 6 2
rect 10 -2 22 2
rect 26 -2 34 2
<< ntransistor >>
rect 9 14 11 34
rect 21 14 23 34
<< ptransistor >>
rect 9 46 11 74
rect 21 46 23 74
<< polycontact >>
rect 6 78 10 82
rect 22 38 26 42
<< ndcontact >>
rect 14 16 18 20
rect 25 25 29 29
rect 25 17 29 21
rect 14 10 18 13
<< pdcontact >>
rect 14 75 18 78
rect 14 68 18 72
rect 25 67 29 71
rect 25 59 29 63
<< m2contact >>
rect 6 86 10 90
rect 22 86 26 90
rect 14 78 18 82
rect 14 6 18 10
rect 6 -2 10 2
rect 22 -2 26 2
<< psubstratepcontact >>
rect 2 -2 6 2
rect 26 -2 30 2
<< nsubstratencontact >>
rect 2 86 6 90
rect 26 86 30 90
<< psubstratepdiff >>
rect 0 2 7 3
rect 25 2 32 3
rect 0 -2 2 2
rect 6 -2 7 2
rect 0 -3 7 -2
rect 25 -2 26 2
rect 30 -2 32 2
rect 25 -3 32 -2
<< nsubstratendiff >>
rect 0 90 7 91
rect 0 86 2 90
rect 6 86 7 90
rect 25 90 32 91
rect 25 86 26 90
rect 30 86 32 90
rect 0 85 7 86
rect 25 85 32 86
<< labels >>
rlabel metal1 16 44 16 44 6 z
rlabel metal1 24 20 24 20 6 z
rlabel metal1 24 44 24 44 6 a
rlabel metal1 24 68 24 68 6 z
rlabel metal2 16 6 16 6 6 vss
rlabel metal2 16 82 16 82 6 vdd
<< end >>
