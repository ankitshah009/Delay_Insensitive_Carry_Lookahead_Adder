magic
tech scmos
timestamp 1180600823
<< checkpaint >>
rect -20 -21 90 120
<< metal1 >>
rect 18 100 22 102
rect -2 88 72 100
rect -2 0 72 12
rect 38 -3 62 0
<< metal2 >>
rect 38 2 62 3
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 38 -3 62 -2
<< metal3 >>
rect 8 98 18 102
rect 22 98 32 102
rect 8 -2 32 98
rect 38 2 62 102
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 38 -3 62 -2
<< m3contact >>
rect 18 98 22 102
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
<< labels >>
rlabel metal1 35 6 35 6 6 vss
rlabel metal1 35 94 35 94 6 vdd
<< end >>
