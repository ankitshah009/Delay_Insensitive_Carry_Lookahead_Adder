magic
tech scmos
timestamp 1179387579
<< checkpaint >>
rect -22 -25 118 105
<< ab >>
rect 0 0 96 80
<< pwell >>
rect -4 -7 100 36
<< nwell >>
rect -4 36 100 87
<< polysilicon >>
rect 12 70 14 74
rect 19 70 21 74
rect 31 70 33 74
rect 38 70 40 74
rect 48 70 50 74
rect 58 70 60 74
rect 68 70 70 74
rect 75 70 77 74
rect 85 70 87 74
rect 12 39 14 42
rect 9 38 15 39
rect 9 34 10 38
rect 14 34 15 38
rect 9 33 15 34
rect 9 30 11 33
rect 19 30 21 42
rect 31 39 33 50
rect 38 47 40 50
rect 48 47 50 50
rect 58 47 60 50
rect 68 47 70 50
rect 38 45 43 47
rect 48 46 61 47
rect 48 45 56 46
rect 41 41 43 45
rect 55 42 56 45
rect 60 42 61 46
rect 55 41 61 42
rect 65 45 70 47
rect 41 39 51 41
rect 31 38 37 39
rect 31 34 32 38
rect 36 35 37 38
rect 49 35 51 39
rect 65 35 67 45
rect 75 39 77 50
rect 85 39 87 42
rect 36 34 44 35
rect 31 33 44 34
rect 49 33 67 35
rect 71 38 77 39
rect 71 34 72 38
rect 76 34 77 38
rect 71 33 77 34
rect 81 38 87 39
rect 81 34 82 38
rect 86 34 87 38
rect 81 33 87 34
rect 42 30 44 33
rect 52 30 54 33
rect 61 30 67 33
rect 28 21 34 22
rect 28 17 29 21
rect 33 17 34 21
rect 28 16 34 17
rect 61 26 62 30
rect 66 26 67 30
rect 84 28 86 33
rect 61 25 67 26
rect 9 11 11 16
rect 19 13 21 16
rect 28 13 30 16
rect 19 11 30 13
rect 42 13 44 18
rect 52 13 54 18
rect 84 10 86 15
<< ndiffusion >>
rect 4 22 9 30
rect 2 21 9 22
rect 2 17 3 21
rect 7 17 9 21
rect 2 16 9 17
rect 11 29 19 30
rect 11 25 13 29
rect 17 25 19 29
rect 11 16 19 25
rect 21 29 28 30
rect 21 25 23 29
rect 27 25 28 29
rect 21 24 28 25
rect 21 16 26 24
rect 36 18 42 30
rect 44 29 52 30
rect 44 25 46 29
rect 50 25 52 29
rect 44 18 52 25
rect 54 22 59 30
rect 77 27 84 28
rect 77 23 78 27
rect 82 23 84 27
rect 77 22 84 23
rect 54 18 62 22
rect 36 14 40 18
rect 34 12 40 14
rect 34 8 35 12
rect 39 8 40 12
rect 34 7 40 8
rect 56 12 62 18
rect 79 15 84 22
rect 86 20 94 28
rect 86 16 88 20
rect 92 16 94 20
rect 86 15 94 16
rect 56 8 57 12
rect 61 8 62 12
rect 56 7 62 8
<< pdiffusion >>
rect 7 62 12 70
rect 5 61 12 62
rect 5 57 6 61
rect 10 57 12 61
rect 5 54 12 57
rect 5 50 6 54
rect 10 50 12 54
rect 5 49 12 50
rect 7 42 12 49
rect 14 42 19 70
rect 21 69 31 70
rect 21 65 24 69
rect 28 65 31 69
rect 21 50 31 65
rect 33 50 38 70
rect 40 55 48 70
rect 40 51 42 55
rect 46 51 48 55
rect 40 50 48 51
rect 50 62 58 70
rect 50 58 52 62
rect 56 58 58 62
rect 50 50 58 58
rect 60 62 68 70
rect 60 58 62 62
rect 66 58 68 62
rect 60 55 68 58
rect 60 51 62 55
rect 66 51 68 55
rect 60 50 68 51
rect 70 50 75 70
rect 77 69 85 70
rect 77 65 79 69
rect 83 65 85 69
rect 77 62 85 65
rect 77 58 79 62
rect 83 58 85 62
rect 77 50 85 58
rect 21 42 26 50
rect 80 42 85 50
rect 87 63 92 70
rect 87 62 94 63
rect 87 58 89 62
rect 93 58 94 62
rect 87 55 94 58
rect 87 51 89 55
rect 93 51 94 55
rect 87 50 94 51
rect 87 42 92 50
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect -2 69 98 78
rect -2 68 24 69
rect 23 65 24 68
rect 28 68 79 69
rect 28 65 29 68
rect 78 65 79 68
rect 83 68 98 69
rect 83 65 84 68
rect 62 62 67 63
rect 6 61 10 62
rect 6 55 10 57
rect 2 54 10 55
rect 25 58 52 62
rect 56 58 57 62
rect 66 58 67 62
rect 78 62 84 65
rect 78 58 79 62
rect 83 58 84 62
rect 89 62 94 63
rect 93 58 94 62
rect 25 54 31 58
rect 62 55 67 58
rect 2 29 6 54
rect 10 50 31 54
rect 34 51 42 55
rect 46 51 62 55
rect 66 51 67 55
rect 89 55 94 58
rect 34 46 38 51
rect 22 42 38 46
rect 22 38 26 42
rect 42 38 46 47
rect 73 46 79 54
rect 93 51 94 55
rect 89 50 94 51
rect 55 42 56 46
rect 60 42 86 46
rect 82 38 86 42
rect 9 34 10 38
rect 14 34 26 38
rect 31 34 32 38
rect 36 34 72 38
rect 76 34 77 38
rect 22 29 26 34
rect 82 33 86 34
rect 2 25 13 29
rect 17 25 18 29
rect 22 25 23 29
rect 27 25 46 29
rect 50 25 51 29
rect 57 26 62 30
rect 66 26 71 30
rect 90 29 94 50
rect 78 27 94 29
rect 82 25 94 27
rect 78 21 82 23
rect 2 17 3 21
rect 7 17 29 21
rect 33 17 82 21
rect 88 20 92 21
rect 88 12 92 16
rect -2 8 35 12
rect 39 8 57 12
rect 61 8 98 12
rect -2 2 98 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
<< ntransistor >>
rect 9 16 11 30
rect 19 16 21 30
rect 42 18 44 30
rect 52 18 54 30
rect 84 15 86 28
<< ptransistor >>
rect 12 42 14 70
rect 19 42 21 70
rect 31 50 33 70
rect 38 50 40 70
rect 48 50 50 70
rect 58 50 60 70
rect 68 50 70 70
rect 75 50 77 70
rect 85 42 87 70
<< polycontact >>
rect 10 34 14 38
rect 56 42 60 46
rect 32 34 36 38
rect 72 34 76 38
rect 82 34 86 38
rect 29 17 33 21
rect 62 26 66 30
<< ndcontact >>
rect 3 17 7 21
rect 13 25 17 29
rect 23 25 27 29
rect 46 25 50 29
rect 78 23 82 27
rect 35 8 39 12
rect 88 16 92 20
rect 57 8 61 12
<< pdcontact >>
rect 6 57 10 61
rect 6 50 10 54
rect 24 65 28 69
rect 42 51 46 55
rect 52 58 56 62
rect 62 58 66 62
rect 62 51 66 55
rect 79 65 83 69
rect 79 58 83 62
rect 89 58 93 62
rect 89 51 93 55
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
rect 90 -2 94 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
rect 90 78 94 82
<< psubstratepdiff >>
rect 0 2 96 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 96 2
rect 0 -3 96 -2
<< nsubstratendiff >>
rect 0 82 96 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 96 82
rect 0 77 96 78
<< labels >>
rlabel ptransistor 13 53 13 53 6 an
rlabel polycontact 31 19 31 19 6 bn
rlabel metal1 4 40 4 40 6 z
rlabel metal1 12 52 12 52 6 z
rlabel metal1 17 36 17 36 6 an
rlabel metal1 20 52 20 52 6 z
rlabel metal1 28 56 28 56 6 z
rlabel metal1 48 6 48 6 6 vss
rlabel metal1 36 27 36 27 6 an
rlabel metal1 36 36 36 36 6 a1
rlabel metal1 44 40 44 40 6 a1
rlabel metal1 52 36 52 36 6 a1
rlabel metal1 36 60 36 60 6 z
rlabel metal1 44 60 44 60 6 z
rlabel metal1 52 60 52 60 6 z
rlabel metal1 48 74 48 74 6 vdd
rlabel metal1 60 28 60 28 6 a2
rlabel metal1 68 28 68 28 6 a2
rlabel metal1 60 36 60 36 6 a1
rlabel metal1 60 44 60 44 6 b
rlabel metal1 68 36 68 36 6 a1
rlabel metal1 68 44 68 44 6 b
rlabel metal1 76 48 76 48 6 b
rlabel metal1 50 53 50 53 6 an
rlabel metal1 64 57 64 57 6 an
rlabel metal1 80 23 80 23 6 bn
rlabel metal1 42 19 42 19 6 bn
rlabel polycontact 84 36 84 36 6 b
rlabel metal1 92 44 92 44 6 bn
<< end >>
