.subckt xaoi21v0x05 a1 a2 b vdd vss z
*   SPICE3 file   created from xaoi21v0x05.ext -      technology: scmos
m00 bn     b      vdd    vdd p w=16u  l=2.3636u ad=92p      pd=46u      as=86.7368p ps=32.8421u
m01 z      b      an     vdd p w=16u  l=2.3636u ad=65.7778p pd=24.8889u as=72p      ps=29.1429u
m02 w1     an     z      vdd p w=20u  l=2.3636u ad=50p      pd=25u      as=82.2222p ps=31.1111u
m03 vdd    bn     w1     vdd p w=20u  l=2.3636u ad=108.421p pd=41.0526u as=50p      ps=25u
m04 an     a2     vdd    vdd p w=20u  l=2.3636u ad=90p      pd=36.4286u as=108.421p ps=41.0526u
m05 vdd    a1     an     vdd p w=20u  l=2.3636u ad=108.421p pd=41.0526u as=90p      ps=36.4286u
m06 bn     b      vss    vss n w=10u  l=2.3636u ad=40p      pd=18u      as=117.5p   ps=47u
m07 z      an     bn     vss n w=10u  l=2.3636u ad=40p      pd=18u      as=40p      ps=18u
m08 an     bn     z      vss n w=10u  l=2.3636u ad=40p      pd=18u      as=40p      ps=18u
m09 w2     a2     an     vss n w=10u  l=2.3636u ad=25p      pd=15u      as=40p      ps=18u
m10 vss    a1     w2     vss n w=10u  l=2.3636u ad=117.5p   pd=47u      as=25p      ps=15u
C0  a2     bn     0.067f
C1  z      b      0.042f
C2  w1     vdd    0.005f
C3  a1     an     0.081f
C4  a2     b      0.018f
C5  a1     vdd    0.016f
C6  bn     an     0.188f
C7  w2     a1     0.009f
C8  vss    z      0.040f
C9  bn     vdd    0.052f
C10 an     b      0.090f
C11 vss    a2     0.011f
C12 b      vdd    0.036f
C13 vss    an     0.033f
C14 z      a2     0.025f
C15 a1     bn     0.034f
C16 z      an     0.428f
C17 vss    vdd    0.006f
C18 z      vdd    0.063f
C19 a1     b      0.012f
C20 a2     an     0.253f
C21 a2     vdd    0.050f
C22 bn     b      0.230f
C23 vss    a1     0.056f
C24 an     vdd    0.345f
C25 z      a1     0.020f
C26 vss    bn     0.153f
C27 z      bn     0.216f
C28 a1     a2     0.097f
C29 w1     an     0.018f
C30 vss    b      0.044f
C32 z      vss    0.011f
C33 a1     vss    0.021f
C34 a2     vss    0.020f
C35 bn     vss    0.049f
C36 an     vss    0.029f
C37 b      vss    0.042f
.ends
