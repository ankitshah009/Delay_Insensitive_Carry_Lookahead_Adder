.subckt nmx3_x4 cmd0 cmd1 i0 i1 i2 nq vdd vss
*   SPICE3 file   created from nmx3_x4.ext -      technology: scmos
m00 w1     i2     w2     vdd p w=20u  l=2.3636u ad=100p     pd=30u      as=120p     ps=38.6667u
m01 w3     cmd1   w1     vdd p w=20u  l=2.3636u ad=136p     pd=44u      as=100p     ps=30u
m02 w4     w5     w3     vdd p w=20u  l=2.3636u ad=60p      pd=26u      as=136p     ps=44u
m03 w2     i1     w4     vdd p w=20u  l=2.3636u ad=120p     pd=38.6667u as=60p      ps=26u
m04 vdd    w6     w2     vdd p w=20u  l=2.3636u ad=131.429p pd=39.5238u as=120p     ps=38.6667u
m05 w7     cmd0   vdd    vdd p w=20u  l=2.3636u ad=60p      pd=26u      as=131.429p ps=39.5238u
m06 w3     i0     w7     vdd p w=20u  l=2.3636u ad=136p     pd=44u      as=60p      ps=26u
m07 w5     cmd1   vdd    vdd p w=14u  l=2.3636u ad=112p     pd=44u      as=92p      ps=27.6667u
m08 w5     cmd1   vss    vss n w=8u   l=2.3636u ad=64p      pd=32u      as=59.7333p ps=21.3333u
m09 vdd    cmd0   w6     vdd p w=14u  l=2.3636u ad=92p      pd=27.6667u as=112p     ps=44u
m10 nq     w8     vdd    vdd p w=40u  l=2.3636u ad=200p     pd=50u      as=262.857p ps=79.0476u
m11 vdd    w8     nq     vdd p w=40u  l=2.3636u ad=262.857p pd=79.0476u as=200p     ps=50u
m12 w8     w3     vdd    vdd p w=20u  l=2.3636u ad=160p     pd=56u      as=131.429p ps=39.5238u
m13 w9     i2     w10    vss n w=12u  l=2.3636u ad=60p      pd=22u      as=80p      ps=30.6667u
m14 w3     w5     w9     vss n w=12u  l=2.3636u ad=100p     pd=37.3333u as=60p      ps=22u
m15 w11    cmd1   w3     vss n w=12u  l=2.3636u ad=36p      pd=18u      as=100p     ps=37.3333u
m16 w10    i1     w11    vss n w=12u  l=2.3636u ad=80p      pd=30.6667u as=36p      ps=18u
m17 vss    cmd0   w6     vss n w=8u   l=2.3636u ad=59.7333p pd=21.3333u as=64p      ps=32u
m18 vss    cmd0   w10    vss n w=12u  l=2.3636u ad=89.6p    pd=32u      as=80p      ps=30.6667u
m19 w12    w6     vss    vss n w=12u  l=2.3636u ad=36p      pd=18u      as=89.6p    ps=32u
m20 w3     i0     w12    vss n w=12u  l=2.3636u ad=100p     pd=37.3333u as=36p      ps=18u
m21 nq     w8     vss    vss n w=20u  l=2.3636u ad=118p     pd=36u      as=149.333p ps=53.3333u
m22 vss    w8     nq     vss n w=20u  l=2.3636u ad=149.333p pd=53.3333u as=118p     ps=36u
m23 w8     w3     vss    vss n w=10u  l=2.3636u ad=80p      pd=36u      as=74.6667p ps=26.6667u
C0  vss    w3     0.465f
C1  vdd    i0     0.026f
C2  vss    i2     0.010f
C3  w3     i1     0.133f
C4  w11    w10    0.011f
C5  i1     i2     0.075f
C6  w5     cmd1   0.502f
C7  nq     vdd    0.200f
C8  w8     cmd0   0.065f
C9  vdd    w6     0.028f
C10 w3     cmd1   0.075f
C11 w2     i1     0.025f
C12 w11    vss    0.006f
C13 cmd1   i2     0.197f
C14 nq     i0     0.029f
C15 vss    w8     0.039f
C16 w4     w2     0.014f
C17 w7     vdd    0.014f
C18 vdd    w5     0.048f
C19 w2     cmd1   0.136f
C20 i0     w6     0.340f
C21 w10    vss    0.434f
C22 w10    i1     0.025f
C23 vss    cmd0   0.017f
C24 nq     w6     0.075f
C25 w1     w2     0.024f
C26 w3     vdd    0.346f
C27 cmd0   i1     0.081f
C28 vdd    i2     0.010f
C29 i0     w5     0.016f
C30 w2     vdd    0.452f
C31 vss    i1     0.017f
C32 w3     i0     0.208f
C33 w10    cmd1   0.006f
C34 w6     w5     0.041f
C35 cmd0   cmd1   0.030f
C36 nq     w3     0.532f
C37 vdd    w8     0.107f
C38 w3     w6     0.515f
C39 vss    cmd1   0.053f
C40 i1     cmd1   0.143f
C41 w6     i2     0.022f
C42 w8     i0     0.026f
C43 vdd    cmd0   0.018f
C44 w3     w5     0.194f
C45 w12    vss    0.011f
C46 w9     w10    0.019f
C47 w5     i2     0.238f
C48 nq     w8     0.084f
C49 i0     cmd0   0.341f
C50 vdd    i1     0.018f
C51 w2     w5     0.079f
C52 w8     w6     0.038f
C53 w3     i2     0.018f
C54 w9     vss    0.010f
C55 w3     w2     0.234f
C56 w4     vdd    0.014f
C57 vss    i0     0.021f
C58 nq     cmd0   0.005f
C59 w10    w6     0.030f
C60 w2     i2     0.013f
C61 vdd    cmd1   0.118f
C62 cmd0   w6     0.333f
C63 i0     i1     0.030f
C64 nq     vss    0.032f
C65 vss    w6     0.091f
C66 w1     vdd    0.023f
C67 w3     w8     0.506f
C68 w10    w5     0.180f
C69 w6     i1     0.129f
C70 cmd0   w5     0.027f
C71 i0     cmd1   0.008f
C72 w10    w3     0.162f
C73 w3     cmd0   0.270f
C74 vss    w5     0.047f
C75 w10    i2     0.017f
C76 w6     cmd1   0.044f
C77 i1     w5     0.198f
C78 cmd0   i2     0.014f
C79 nq     vss    0.015f
C81 w3     vss    0.109f
C83 w8     vss    0.062f
C84 i0     vss    0.051f
C85 cmd0   vss    0.067f
C86 w6     vss    0.059f
C87 i1     vss    0.040f
C88 w5     vss    0.059f
C89 cmd1   vss    0.073f
C90 i2     vss    0.037f
.ends
