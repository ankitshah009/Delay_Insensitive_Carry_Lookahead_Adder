magic
tech scmos
timestamp 1179385899
<< checkpaint >>
rect -22 -22 46 94
<< ab >>
rect 0 0 24 72
<< pwell >>
rect -4 -4 28 32
<< nwell >>
rect -4 32 28 76
<< polysilicon >>
rect 9 66 11 70
rect 9 35 11 39
rect 9 34 15 35
rect 9 30 10 34
rect 14 30 15 34
rect 9 29 15 30
rect 9 26 11 29
rect 9 9 11 14
<< ndiffusion >>
rect 2 25 9 26
rect 2 21 3 25
rect 7 21 9 25
rect 2 20 9 21
rect 4 14 9 20
rect 11 19 19 26
rect 11 15 13 19
rect 17 15 19 19
rect 11 14 19 15
<< pdiffusion >>
rect 4 52 9 66
rect 2 51 9 52
rect 2 47 3 51
rect 7 47 9 51
rect 2 44 9 47
rect 2 40 3 44
rect 7 40 9 44
rect 2 39 9 40
rect 11 65 19 66
rect 11 61 13 65
rect 17 61 19 65
rect 11 58 19 61
rect 11 54 13 58
rect 17 54 19 58
rect 11 39 19 54
<< metal1 >>
rect -2 65 26 72
rect -2 64 13 65
rect 12 61 13 64
rect 17 64 26 65
rect 17 61 18 64
rect 12 58 18 61
rect 12 54 13 58
rect 17 54 18 58
rect 2 47 3 51
rect 7 47 14 51
rect 2 45 14 47
rect 2 44 7 45
rect 2 40 3 44
rect 2 39 7 40
rect 2 25 6 39
rect 18 35 22 43
rect 10 34 22 35
rect 14 30 22 34
rect 10 29 22 30
rect 2 21 3 25
rect 7 21 8 25
rect 2 20 8 21
rect 13 19 17 20
rect 13 8 17 15
rect -2 0 26 8
<< ntransistor >>
rect 9 14 11 26
<< ptransistor >>
rect 9 39 11 66
<< polycontact >>
rect 10 30 14 34
<< ndcontact >>
rect 3 21 7 25
rect 13 15 17 19
<< pdcontact >>
rect 3 47 7 51
rect 3 40 7 44
rect 13 61 17 65
rect 13 54 17 58
<< labels >>
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 4 12 4 6 vss
rlabel polycontact 12 32 12 32 6 a
rlabel metal1 12 48 12 48 6 z
rlabel metal1 12 68 12 68 6 vdd
rlabel metal1 20 36 20 36 6 a
<< end >>
