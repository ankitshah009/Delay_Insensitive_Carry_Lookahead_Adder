magic
tech scmos
timestamp 1185038990
<< checkpaint >>
rect -22 -24 92 124
<< ab >>
rect 0 0 70 100
<< pwell >>
rect -2 -4 72 49
<< nwell >>
rect -2 49 72 104
<< polysilicon >>
rect 35 95 37 98
rect 47 95 49 98
rect 11 85 13 88
rect 23 85 25 88
rect 11 43 13 65
rect 23 43 25 65
rect 57 82 63 83
rect 57 78 58 82
rect 62 78 63 82
rect 57 77 63 78
rect 57 75 59 77
rect 35 43 37 55
rect 47 43 49 55
rect 7 42 13 43
rect 7 38 8 42
rect 12 38 13 42
rect 7 37 13 38
rect 17 42 25 43
rect 17 38 18 42
rect 22 38 25 42
rect 17 37 25 38
rect 33 42 53 43
rect 33 38 48 42
rect 52 38 53 42
rect 33 37 53 38
rect 11 35 13 37
rect 21 35 23 37
rect 33 25 35 37
rect 45 25 47 37
rect 57 25 59 55
rect 11 12 13 15
rect 21 12 23 15
rect 57 12 59 15
rect 33 2 35 5
rect 45 2 47 5
<< ndiffusion >>
rect 3 22 11 35
rect 3 18 4 22
rect 8 18 11 22
rect 3 15 11 18
rect 13 15 21 35
rect 23 25 31 35
rect 23 15 33 25
rect 25 12 33 15
rect 25 8 26 12
rect 30 8 33 12
rect 25 5 33 8
rect 35 22 45 25
rect 35 18 38 22
rect 42 18 45 22
rect 35 5 45 18
rect 47 15 57 25
rect 59 22 67 25
rect 59 18 62 22
rect 66 18 67 22
rect 59 15 67 18
rect 47 12 55 15
rect 47 8 50 12
rect 54 8 55 12
rect 47 5 55 8
<< pdiffusion >>
rect 3 92 9 93
rect 3 88 4 92
rect 8 88 9 92
rect 27 92 35 95
rect 27 88 28 92
rect 32 88 35 92
rect 3 85 9 88
rect 27 85 35 88
rect 3 82 11 85
rect 3 78 4 82
rect 8 78 11 82
rect 3 65 11 78
rect 13 82 23 85
rect 13 78 16 82
rect 20 78 23 82
rect 13 65 23 78
rect 25 65 35 85
rect 27 55 35 65
rect 37 72 47 95
rect 37 68 40 72
rect 44 68 47 72
rect 37 62 47 68
rect 37 58 40 62
rect 44 58 47 62
rect 37 55 47 58
rect 49 92 57 95
rect 49 88 52 92
rect 56 88 57 92
rect 49 85 57 88
rect 49 75 55 85
rect 49 55 57 75
rect 59 72 67 75
rect 59 68 62 72
rect 66 68 67 72
rect 59 62 67 68
rect 59 58 62 62
rect 66 58 67 62
rect 59 55 67 58
<< metal1 >>
rect -2 92 72 101
rect -2 88 4 92
rect 8 88 28 92
rect 32 88 52 92
rect 56 88 72 92
rect -2 87 72 88
rect 3 82 9 87
rect 3 78 4 82
rect 8 78 9 82
rect 3 77 9 78
rect 15 82 21 83
rect 57 82 63 83
rect 15 78 16 82
rect 20 78 58 82
rect 62 78 63 82
rect 15 77 21 78
rect 7 42 13 72
rect 7 38 8 42
rect 12 38 13 42
rect 7 28 13 38
rect 17 42 23 72
rect 17 38 18 42
rect 22 38 23 42
rect 17 28 23 38
rect 3 22 9 23
rect 28 22 32 78
rect 57 77 63 78
rect 3 18 4 22
rect 8 18 32 22
rect 37 72 45 73
rect 37 68 40 72
rect 44 68 45 72
rect 37 67 45 68
rect 61 72 67 73
rect 61 68 62 72
rect 66 68 67 72
rect 61 67 67 68
rect 37 63 43 67
rect 62 63 66 67
rect 37 62 45 63
rect 37 58 40 62
rect 44 58 45 62
rect 37 57 45 58
rect 61 62 67 63
rect 61 58 62 62
rect 66 58 67 62
rect 61 57 67 58
rect 37 22 43 57
rect 47 42 53 43
rect 62 42 66 57
rect 47 38 48 42
rect 52 38 66 42
rect 47 37 53 38
rect 62 23 66 38
rect 37 18 38 22
rect 42 18 43 22
rect 3 17 9 18
rect 37 17 43 18
rect 61 22 67 23
rect 61 18 62 22
rect 66 18 67 22
rect 61 17 67 18
rect -2 12 72 13
rect -2 8 26 12
rect 30 8 50 12
rect 54 8 72 12
rect -2 4 4 8
rect 8 4 14 8
rect 18 4 72 8
rect -2 -1 72 4
<< ntransistor >>
rect 11 15 13 35
rect 21 15 23 35
rect 33 5 35 25
rect 45 5 47 25
rect 57 15 59 25
<< ptransistor >>
rect 11 65 13 85
rect 23 65 25 85
rect 35 55 37 95
rect 47 55 49 95
rect 57 55 59 75
<< polycontact >>
rect 58 78 62 82
rect 8 38 12 42
rect 18 38 22 42
rect 48 38 52 42
<< ndcontact >>
rect 4 18 8 22
rect 26 8 30 12
rect 38 18 42 22
rect 62 18 66 22
rect 50 8 54 12
<< pdcontact >>
rect 4 88 8 92
rect 28 88 32 92
rect 4 78 8 82
rect 16 78 20 82
rect 40 68 44 72
rect 40 58 44 62
rect 52 88 56 92
rect 62 68 66 72
rect 62 58 66 62
<< psubstratepcontact >>
rect 4 4 8 8
rect 14 4 18 8
<< psubstratepdiff >>
rect 3 8 19 9
rect 3 4 4 8
rect 8 4 14 8
rect 18 4 19 8
rect 3 3 19 4
<< labels >>
rlabel metal1 10 50 10 50 6 i0
rlabel metal1 10 50 10 50 6 i0
rlabel metal1 20 50 20 50 6 i1
rlabel metal1 20 50 20 50 6 i1
rlabel metal1 35 6 35 6 6 vss
rlabel metal1 35 6 35 6 6 vss
rlabel metal1 40 45 40 45 6 nq
rlabel metal1 40 45 40 45 6 nq
rlabel metal1 35 94 35 94 6 vdd
rlabel metal1 35 94 35 94 6 vdd
<< end >>
