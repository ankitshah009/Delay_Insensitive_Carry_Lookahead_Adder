magic
tech scmos
timestamp 1179387197
<< checkpaint >>
rect -22 -22 62 94
<< ab >>
rect 0 0 40 72
<< pwell >>
rect -4 -4 44 32
<< nwell >>
rect -4 32 44 76
<< polysilicon >>
rect 9 59 11 64
rect 19 59 25 60
rect 19 55 20 59
rect 24 55 25 59
rect 19 54 25 55
rect 22 51 24 54
rect 29 51 31 56
rect 9 37 11 41
rect 9 36 15 37
rect 9 32 10 36
rect 14 32 15 36
rect 22 33 24 41
rect 9 31 15 32
rect 19 31 24 33
rect 29 35 31 41
rect 29 34 35 35
rect 9 26 11 31
rect 19 26 21 31
rect 29 30 30 34
rect 34 30 35 34
rect 29 29 35 30
rect 29 26 31 29
rect 9 12 11 17
rect 19 15 21 20
rect 29 15 31 20
<< ndiffusion >>
rect 2 25 9 26
rect 2 21 3 25
rect 7 21 9 25
rect 2 20 9 21
rect 4 17 9 20
rect 11 20 19 26
rect 21 25 29 26
rect 21 21 23 25
rect 27 21 29 25
rect 21 20 29 21
rect 31 25 38 26
rect 31 21 33 25
rect 37 21 38 25
rect 31 20 38 21
rect 11 17 17 20
rect 13 13 17 17
rect 13 12 19 13
rect 13 8 14 12
rect 18 8 19 12
rect 13 7 19 8
<< pdiffusion >>
rect 13 68 19 69
rect 13 64 14 68
rect 18 64 19 68
rect 13 62 19 64
rect 13 59 17 62
rect 4 54 9 59
rect 2 53 9 54
rect 2 49 3 53
rect 7 49 9 53
rect 2 46 9 49
rect 2 42 3 46
rect 7 42 9 46
rect 2 41 9 42
rect 11 51 17 59
rect 11 41 22 51
rect 24 41 29 51
rect 31 50 38 51
rect 31 46 33 50
rect 37 46 38 50
rect 31 45 38 46
rect 31 41 36 45
<< metal1 >>
rect -2 68 42 72
rect -2 64 14 68
rect 18 64 24 68
rect 28 64 32 68
rect 36 64 42 68
rect 2 54 6 59
rect 10 55 20 59
rect 24 55 25 59
rect 2 53 7 54
rect 2 49 3 53
rect 2 46 7 49
rect 2 42 3 46
rect 10 53 25 55
rect 10 45 14 53
rect 18 46 33 50
rect 37 46 38 50
rect 2 41 7 42
rect 2 27 6 41
rect 18 37 22 46
rect 10 36 22 37
rect 14 32 22 36
rect 34 35 38 43
rect 10 31 22 32
rect 2 25 14 27
rect 2 21 3 25
rect 7 21 14 25
rect 18 25 22 31
rect 26 34 38 35
rect 26 30 30 34
rect 34 30 38 34
rect 26 29 38 30
rect 18 21 23 25
rect 27 21 28 25
rect 32 21 33 25
rect 37 21 38 25
rect 14 12 18 13
rect 32 8 38 21
rect -2 4 24 8
rect 28 4 32 8
rect 36 4 42 8
rect -2 0 42 4
<< ntransistor >>
rect 9 17 11 26
rect 19 20 21 26
rect 29 20 31 26
<< ptransistor >>
rect 9 41 11 59
rect 22 41 24 51
rect 29 41 31 51
<< polycontact >>
rect 20 55 24 59
rect 10 32 14 36
rect 30 30 34 34
<< ndcontact >>
rect 3 21 7 25
rect 23 21 27 25
rect 33 21 37 25
rect 14 8 18 12
<< pdcontact >>
rect 14 64 18 68
rect 3 49 7 53
rect 3 42 7 46
rect 33 46 37 50
<< psubstratepcontact >>
rect 24 4 28 8
rect 32 4 36 8
<< nsubstratencontact >>
rect 24 64 28 68
rect 32 64 36 68
<< psubstratepdiff >>
rect 23 8 37 9
rect 23 4 24 8
rect 28 4 32 8
rect 36 4 37 8
rect 23 3 37 4
<< nsubstratendiff >>
rect 23 68 37 69
rect 23 64 24 68
rect 28 64 32 68
rect 36 64 37 68
rect 23 63 37 64
<< labels >>
rlabel polycontact 12 34 12 34 6 zn
rlabel metal1 4 40 4 40 6 z
rlabel metal1 12 24 12 24 6 z
rlabel metal1 12 52 12 52 6 a
rlabel metal1 20 4 20 4 6 vss
rlabel metal1 23 23 23 23 6 zn
rlabel metal1 28 32 28 32 6 b
rlabel metal1 16 34 16 34 6 zn
rlabel metal1 20 56 20 56 6 a
rlabel metal1 20 68 20 68 6 vdd
rlabel metal1 36 36 36 36 6 b
rlabel metal1 28 48 28 48 6 zn
<< end >>
