magic
tech scmos
timestamp 1179387081
<< checkpaint >>
rect -22 -22 78 94
<< ab >>
rect 0 0 56 72
<< pwell >>
rect -4 -4 60 32
<< nwell >>
rect -4 32 60 76
<< polysilicon >>
rect 13 66 15 70
rect 21 66 23 70
rect 31 66 33 70
rect 39 66 41 70
rect 13 36 15 39
rect 21 36 23 39
rect 9 35 15 36
rect 9 31 10 35
rect 14 31 15 35
rect 9 30 15 31
rect 19 35 25 36
rect 31 35 33 39
rect 39 36 41 39
rect 39 35 48 36
rect 19 31 20 35
rect 24 31 25 35
rect 19 30 25 31
rect 29 34 35 35
rect 29 30 30 34
rect 34 30 35 34
rect 39 31 43 35
rect 47 31 48 35
rect 39 30 48 31
rect 9 26 11 30
rect 19 26 21 30
rect 29 29 35 30
rect 29 23 31 29
rect 41 23 43 30
rect 9 7 11 12
rect 19 7 21 12
rect 29 7 31 12
rect 41 7 43 12
<< ndiffusion >>
rect 4 18 9 26
rect 2 17 9 18
rect 2 13 3 17
rect 7 13 9 17
rect 2 12 9 13
rect 11 25 19 26
rect 11 21 13 25
rect 17 21 19 25
rect 11 12 19 21
rect 21 23 26 26
rect 21 17 29 23
rect 21 13 23 17
rect 27 13 29 17
rect 21 12 29 13
rect 31 12 41 23
rect 43 18 48 23
rect 43 17 50 18
rect 43 13 45 17
rect 49 13 50 17
rect 43 12 50 13
rect 33 8 39 12
rect 33 4 34 8
rect 38 4 39 8
rect 33 3 39 4
<< pdiffusion >>
rect 5 65 13 66
rect 5 61 7 65
rect 11 61 13 65
rect 5 39 13 61
rect 15 39 21 66
rect 23 58 31 66
rect 23 54 25 58
rect 29 54 31 58
rect 23 39 31 54
rect 33 39 39 66
rect 41 65 48 66
rect 41 61 43 65
rect 47 61 48 65
rect 41 58 48 61
rect 41 54 43 58
rect 47 54 48 58
rect 41 39 48 54
<< metal1 >>
rect -2 65 58 72
rect -2 64 7 65
rect 6 61 7 64
rect 11 64 43 65
rect 11 61 12 64
rect 42 61 43 64
rect 47 64 58 65
rect 47 61 48 64
rect 2 54 25 58
rect 29 54 30 58
rect 2 25 6 54
rect 34 50 38 59
rect 42 58 48 61
rect 42 54 43 58
rect 47 54 48 58
rect 10 46 23 50
rect 34 46 47 50
rect 10 35 14 46
rect 10 29 14 31
rect 18 38 39 42
rect 18 35 24 38
rect 18 31 20 35
rect 43 35 47 46
rect 18 29 24 31
rect 29 30 30 34
rect 34 30 39 34
rect 43 30 47 31
rect 33 26 39 30
rect 2 21 13 25
rect 17 21 18 25
rect 33 22 47 26
rect 2 13 3 17
rect 7 13 23 17
rect 27 13 45 17
rect 49 13 50 17
rect -2 4 34 8
rect 38 4 58 8
rect -2 0 58 4
<< ntransistor >>
rect 9 12 11 26
rect 19 12 21 26
rect 29 12 31 23
rect 41 12 43 23
<< ptransistor >>
rect 13 39 15 66
rect 21 39 23 66
rect 31 39 33 66
rect 39 39 41 66
<< polycontact >>
rect 10 31 14 35
rect 20 31 24 35
rect 30 30 34 34
rect 43 31 47 35
<< ndcontact >>
rect 3 13 7 17
rect 13 21 17 25
rect 23 13 27 17
rect 45 13 49 17
rect 34 4 38 8
<< pdcontact >>
rect 7 61 11 65
rect 25 54 29 58
rect 43 61 47 65
rect 43 54 47 58
<< labels >>
rlabel metal1 4 36 4 36 6 z
rlabel metal1 20 32 20 32 6 b2
rlabel metal1 12 36 12 36 6 b1
rlabel metal1 20 48 20 48 6 b1
rlabel metal1 20 56 20 56 6 z
rlabel metal1 12 56 12 56 6 z
rlabel metal1 28 4 28 4 6 vss
rlabel metal1 36 28 36 28 6 a2
rlabel metal1 36 40 36 40 6 b2
rlabel metal1 28 40 28 40 6 b2
rlabel metal1 36 56 36 56 6 a1
rlabel metal1 28 68 28 68 6 vdd
rlabel ndcontact 26 15 26 15 6 n3
rlabel metal1 44 24 44 24 6 a2
rlabel metal1 44 48 44 48 6 a1
<< end >>
