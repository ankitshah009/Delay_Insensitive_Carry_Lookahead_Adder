magic
tech scmos
timestamp 1179386791
<< checkpaint >>
rect -22 -25 54 105
<< ab >>
rect 0 0 32 80
<< pwell >>
rect -4 -7 36 36
<< nwell >>
rect -4 36 36 87
<< polysilicon >>
rect 12 61 14 65
rect 19 61 21 66
rect 12 43 14 46
rect 9 42 15 43
rect 9 38 10 42
rect 14 38 15 42
rect 9 37 15 38
rect 19 40 21 46
rect 19 39 25 40
rect 10 26 12 37
rect 19 35 20 39
rect 24 35 25 39
rect 19 34 25 35
rect 20 26 22 34
rect 10 15 12 19
rect 20 15 22 19
<< ndiffusion >>
rect 2 24 10 26
rect 2 20 3 24
rect 7 20 10 24
rect 2 19 10 20
rect 12 25 20 26
rect 12 21 14 25
rect 18 21 20 25
rect 12 19 20 21
rect 22 24 30 26
rect 22 20 25 24
rect 29 20 30 24
rect 22 19 30 20
<< pdiffusion >>
rect 5 60 12 61
rect 5 56 6 60
rect 10 56 12 60
rect 5 55 12 56
rect 7 46 12 55
rect 14 46 19 61
rect 21 60 30 61
rect 21 56 25 60
rect 29 56 30 60
rect 21 46 30 56
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect -2 68 34 78
rect 2 33 6 63
rect 25 60 29 68
rect 10 56 11 60
rect 25 55 29 56
rect 18 47 22 55
rect 10 43 22 47
rect 10 42 14 43
rect 26 39 30 47
rect 10 37 14 38
rect 18 35 20 39
rect 24 35 30 39
rect 18 33 30 35
rect 2 29 14 33
rect 3 24 7 25
rect 10 21 14 29
rect 18 21 19 25
rect 25 24 29 25
rect 3 12 7 20
rect 25 12 29 20
rect -2 2 34 12
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
<< ntransistor >>
rect 10 19 12 26
rect 20 19 22 26
<< ptransistor >>
rect 12 46 14 61
rect 19 46 21 61
<< polycontact >>
rect 10 38 14 42
rect 20 35 24 39
<< ndcontact >>
rect 3 20 7 24
rect 14 21 18 25
rect 25 20 29 24
<< pdcontact >>
rect 6 56 10 60
rect 25 56 29 60
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
<< psubstratepdiff >>
rect 0 2 32 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 32 2
rect 0 -3 32 -2
<< nsubstratendiff >>
rect 0 82 32 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 32 82
rect 0 77 32 78
<< labels >>
rlabel metal1 4 48 4 48 6 z
rlabel metal1 12 28 12 28 6 z
rlabel metal1 12 44 12 44 6 b
rlabel metal1 16 6 16 6 6 vss
rlabel metal1 20 36 20 36 6 a
rlabel metal1 20 52 20 52 6 b
rlabel metal1 16 74 16 74 6 vdd
rlabel metal1 28 40 28 40 6 a
<< end >>
