.subckt nao22_x1 i0 i1 i2 nq vdd vss
*   SPICE3 file   created from nao22_x1.ext -      technology: scmos
m00 w1     i0     vdd    vdd p w=40u  l=2.3636u ad=200p     pd=50u      as=320p     ps=96u
m01 nq     i1     w1     vdd p w=40u  l=2.3636u ad=200p     pd=50u      as=200p     ps=50u
m02 vdd    i2     nq     vdd p w=40u  l=2.3636u ad=320p     pd=96u      as=200p     ps=50u
m03 nq     i0     w2     vss n w=20u  l=2.3636u ad=124p     pd=38u      as=120p     ps=38.6667u
m04 w2     i1     nq     vss n w=20u  l=2.3636u ad=120p     pd=38.6667u as=124p     ps=38u
m05 vss    i2     w2     vss n w=20u  l=2.3636u ad=160p     pd=56u      as=120p     ps=38.6667u
C0  w2     i2     0.039f
C1  vss    vdd    0.015f
C2  w2     i0     0.018f
C3  w1     vdd    0.023f
C4  nq     i2     0.417f
C5  vss    i1     0.013f
C6  w1     i1     0.054f
C7  vdd    i2     0.203f
C8  nq     i0     0.098f
C9  vdd    i0     0.105f
C10 i2     i1     0.157f
C11 w2     nq     0.138f
C12 i1     i0     0.416f
C13 nq     vdd    0.119f
C14 vss    i2     0.134f
C15 w2     i1     0.017f
C16 vss    i0     0.013f
C17 nq     i1     0.393f
C18 vdd    i1     0.073f
C19 w1     i0     0.014f
C20 w2     vss    0.254f
C21 i2     i0     0.084f
C22 vss    nq     0.082f
C24 nq     vss    0.023f
C26 i2     vss    0.040f
C27 i1     vss    0.032f
C28 i0     vss    0.026f
.ends
