magic
tech scmos
timestamp 1179386097
<< checkpaint >>
rect -22 -25 86 105
<< ab >>
rect 0 0 64 80
<< pwell >>
rect -4 -7 68 36
<< nwell >>
rect -4 36 68 87
<< polysilicon >>
rect 20 72 55 74
rect 10 54 12 59
rect 20 54 22 72
rect 53 63 55 72
rect 30 62 36 63
rect 30 58 31 62
rect 35 58 36 62
rect 30 57 36 58
rect 30 54 32 57
rect 40 54 42 59
rect 53 46 55 57
rect 50 45 56 46
rect 10 39 12 42
rect 2 38 12 39
rect 20 38 22 42
rect 2 34 3 38
rect 7 34 12 38
rect 30 34 32 42
rect 2 33 12 34
rect 10 23 12 33
rect 20 32 32 34
rect 40 39 42 42
rect 50 41 51 45
rect 55 41 56 45
rect 50 40 56 41
rect 40 38 46 39
rect 40 34 41 38
rect 45 34 46 38
rect 40 33 46 34
rect 20 23 22 32
rect 30 23 32 28
rect 40 23 42 33
rect 53 27 55 40
rect 53 18 55 21
rect 10 12 12 17
rect 20 12 22 17
rect 30 9 32 17
rect 40 13 42 17
rect 51 15 55 18
rect 51 9 53 15
rect 30 7 53 9
<< ndiffusion >>
rect 44 23 53 27
rect 2 22 10 23
rect 2 18 3 22
rect 7 18 10 22
rect 2 17 10 18
rect 12 22 20 23
rect 12 18 14 22
rect 18 18 20 22
rect 12 17 20 18
rect 22 22 30 23
rect 22 18 24 22
rect 28 18 30 22
rect 22 17 30 18
rect 32 22 40 23
rect 32 18 34 22
rect 38 18 40 22
rect 32 17 40 18
rect 42 22 53 23
rect 42 18 44 22
rect 48 21 53 22
rect 55 26 62 27
rect 55 22 57 26
rect 61 22 62 26
rect 55 21 62 22
rect 48 18 49 21
rect 42 17 49 18
<< pdiffusion >>
rect 2 63 8 64
rect 2 59 3 63
rect 7 59 8 63
rect 2 54 8 59
rect 44 69 50 70
rect 44 65 45 69
rect 49 65 50 69
rect 44 63 50 65
rect 44 57 53 63
rect 55 62 62 63
rect 55 58 57 62
rect 61 58 62 62
rect 55 57 62 58
rect 44 54 50 57
rect 2 42 10 54
rect 12 47 20 54
rect 12 43 14 47
rect 18 43 20 47
rect 12 42 20 43
rect 22 47 30 54
rect 22 43 24 47
rect 28 43 30 47
rect 22 42 30 43
rect 32 47 40 54
rect 32 43 34 47
rect 38 43 40 47
rect 32 42 40 43
rect 42 49 50 54
rect 42 42 48 49
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect -2 69 66 78
rect -2 68 45 69
rect 3 63 7 68
rect 44 65 45 68
rect 49 68 66 69
rect 49 65 50 68
rect 3 58 7 59
rect 30 58 31 62
rect 35 58 57 62
rect 61 58 62 62
rect 2 50 15 54
rect 2 39 6 50
rect 26 48 30 55
rect 41 50 54 54
rect 24 47 30 48
rect 13 43 14 47
rect 18 43 20 47
rect 2 38 7 39
rect 2 34 3 38
rect 2 33 7 34
rect 3 22 7 23
rect 16 22 20 43
rect 28 43 30 47
rect 24 42 30 43
rect 26 23 30 42
rect 13 18 14 22
rect 18 18 20 22
rect 24 22 30 23
rect 28 18 30 22
rect 33 43 34 47
rect 38 43 39 47
rect 50 46 54 50
rect 50 45 55 46
rect 33 22 37 43
rect 50 41 51 45
rect 50 40 55 41
rect 41 38 46 39
rect 45 34 46 38
rect 41 33 46 34
rect 42 31 46 33
rect 42 25 54 31
rect 58 27 62 58
rect 57 26 62 27
rect 61 22 62 26
rect 33 18 34 22
rect 38 18 39 22
rect 43 18 44 22
rect 48 18 49 22
rect 57 21 62 22
rect 3 12 7 18
rect 24 17 30 18
rect 43 12 49 18
rect -2 2 66 12
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
<< ntransistor >>
rect 10 17 12 23
rect 20 17 22 23
rect 30 17 32 23
rect 40 17 42 23
rect 53 21 55 27
<< ptransistor >>
rect 53 57 55 63
rect 10 42 12 54
rect 20 42 22 54
rect 30 42 32 54
rect 40 42 42 54
<< polycontact >>
rect 31 58 35 62
rect 3 34 7 38
rect 51 41 55 45
rect 41 34 45 38
<< ndcontact >>
rect 3 18 7 22
rect 14 18 18 22
rect 24 18 28 22
rect 34 18 38 22
rect 44 18 48 22
rect 57 22 61 26
<< pdcontact >>
rect 3 59 7 63
rect 45 65 49 69
rect 57 58 61 62
rect 14 43 18 47
rect 24 43 28 47
rect 34 43 38 47
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
<< psubstratepdiff >>
rect 0 2 64 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 64 2
rect 0 -3 64 -2
<< nsubstratendiff >>
rect 0 82 64 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 64 82
rect 0 77 64 78
<< labels >>
rlabel polycontact 33 60 33 60 6 sn
rlabel metal1 4 40 4 40 6 a0
rlabel metal1 18 32 18 32 6 a0n
rlabel pdcontact 16 45 16 45 6 a0n
rlabel metal1 12 52 12 52 6 a0
rlabel metal1 32 6 32 6 6 vss
rlabel metal1 35 32 35 32 6 a1n
rlabel metal1 28 36 28 36 6 z
rlabel metal1 32 74 32 74 6 vdd
rlabel metal1 44 32 44 32 6 a1
rlabel pdcontact 36 45 36 45 6 a1n
rlabel metal1 44 52 44 52 6 s
rlabel metal1 52 28 52 28 6 a1
rlabel polycontact 52 44 52 44 6 s
rlabel metal1 60 41 60 41 6 sn
rlabel metal1 46 60 46 60 6 sn
<< end >>
