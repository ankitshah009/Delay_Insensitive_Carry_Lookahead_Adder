magic
tech scmos
timestamp 1179384990
<< checkpaint >>
rect -22 -25 78 105
<< ab >>
rect 0 0 56 80
<< pwell >>
rect -4 -7 60 36
<< nwell >>
rect -4 36 60 87
<< polysilicon >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 67 31 72
rect 39 67 41 72
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 39 39 41 42
rect 9 38 22 39
rect 9 34 15 38
rect 19 34 22 38
rect 9 33 22 34
rect 28 38 34 39
rect 28 34 29 38
rect 33 34 34 38
rect 28 33 34 34
rect 10 30 12 33
rect 20 30 22 33
rect 32 30 34 33
rect 39 38 47 39
rect 39 34 42 38
rect 46 34 47 38
rect 39 33 47 34
rect 39 30 41 33
rect 10 11 12 16
rect 20 11 22 16
rect 32 6 34 10
rect 39 6 41 10
<< ndiffusion >>
rect 2 16 10 30
rect 12 22 20 30
rect 12 18 14 22
rect 18 18 20 22
rect 12 16 20 18
rect 22 16 32 30
rect 2 12 8 16
rect 2 8 3 12
rect 7 8 8 12
rect 24 15 32 16
rect 24 11 25 15
rect 29 11 32 15
rect 24 10 32 11
rect 34 10 39 30
rect 41 23 46 30
rect 41 22 48 23
rect 41 18 43 22
rect 47 18 48 22
rect 41 17 48 18
rect 41 10 46 17
rect 2 7 8 8
<< pdiffusion >>
rect 2 69 9 70
rect 2 65 3 69
rect 7 65 9 69
rect 2 62 9 65
rect 2 58 3 62
rect 7 58 9 62
rect 2 42 9 58
rect 11 62 19 70
rect 11 58 13 62
rect 17 58 19 62
rect 11 55 19 58
rect 11 51 13 55
rect 17 51 19 55
rect 11 42 19 51
rect 21 67 27 70
rect 21 66 29 67
rect 21 62 23 66
rect 27 62 29 66
rect 21 42 29 62
rect 31 62 39 67
rect 31 58 33 62
rect 37 58 39 62
rect 31 55 39 58
rect 31 51 33 55
rect 37 51 39 55
rect 31 42 39 51
rect 41 66 48 67
rect 41 62 43 66
rect 47 62 48 66
rect 41 58 48 62
rect 41 54 43 58
rect 47 54 48 58
rect 41 42 48 54
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect -2 69 58 78
rect -2 68 3 69
rect 2 65 3 68
rect 7 68 58 69
rect 7 65 8 68
rect 2 62 8 65
rect 23 66 27 68
rect 2 58 3 62
rect 7 58 8 62
rect 13 62 17 63
rect 43 66 47 68
rect 23 61 27 62
rect 33 62 37 63
rect 13 55 17 58
rect 2 51 13 55
rect 33 55 37 58
rect 2 50 17 51
rect 23 51 33 54
rect 43 58 47 62
rect 43 53 47 54
rect 23 50 37 51
rect 2 22 6 50
rect 23 46 27 50
rect 15 42 27 46
rect 33 42 47 46
rect 15 38 19 42
rect 41 38 47 42
rect 25 34 29 38
rect 15 30 19 34
rect 33 30 37 38
rect 41 34 42 38
rect 46 34 47 38
rect 15 26 28 30
rect 33 26 47 30
rect 24 22 28 26
rect 2 18 14 22
rect 18 18 19 22
rect 24 18 43 22
rect 47 18 48 22
rect 2 17 19 18
rect 24 12 25 15
rect -2 8 3 12
rect 7 11 25 12
rect 29 12 30 15
rect 29 11 58 12
rect 7 8 58 11
rect -2 2 58 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
<< ntransistor >>
rect 10 16 12 30
rect 20 16 22 30
rect 32 10 34 30
rect 39 10 41 30
<< ptransistor >>
rect 9 42 11 70
rect 19 42 21 70
rect 29 42 31 67
rect 39 42 41 67
<< polycontact >>
rect 15 34 19 38
rect 29 34 33 38
rect 42 34 46 38
<< ndcontact >>
rect 14 18 18 22
rect 3 8 7 12
rect 25 11 29 15
rect 43 18 47 22
<< pdcontact >>
rect 3 65 7 69
rect 3 58 7 62
rect 13 58 17 62
rect 13 51 17 55
rect 23 62 27 66
rect 33 58 37 62
rect 33 51 37 55
rect 43 62 47 66
rect 43 54 47 58
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
<< psubstratepdiff >>
rect 0 2 56 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 56 2
rect 0 -3 56 -2
<< nsubstratendiff >>
rect 0 82 56 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 56 82
rect 0 77 56 78
<< labels >>
rlabel polysilicon 15 36 15 36 6 zn
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 20 12 20 6 z
rlabel polycontact 17 36 17 36 6 zn
rlabel metal1 12 52 12 52 6 z
rlabel metal1 28 6 28 6 6 vss
rlabel metal1 28 36 28 36 6 a
rlabel metal1 36 28 36 28 6 a
rlabel metal1 36 44 36 44 6 b
rlabel metal1 35 56 35 56 6 zn
rlabel metal1 28 74 28 74 6 vdd
rlabel metal1 36 20 36 20 6 zn
rlabel metal1 44 28 44 28 6 a
rlabel metal1 44 40 44 40 6 b
<< end >>
