magic
tech scmos
timestamp 1179385026
<< checkpaint >>
rect -22 -25 62 105
<< ab >>
rect 0 0 40 80
<< pwell >>
rect -4 -7 44 36
<< nwell >>
rect -4 36 44 87
<< polysilicon >>
rect 9 60 11 65
rect 19 56 21 61
rect 29 56 31 61
rect 9 39 11 42
rect 19 39 21 50
rect 29 47 31 50
rect 29 46 35 47
rect 29 42 30 46
rect 34 42 35 46
rect 29 41 35 42
rect 9 38 15 39
rect 9 34 10 38
rect 14 34 15 38
rect 9 33 15 34
rect 19 38 25 39
rect 19 34 20 38
rect 24 34 25 38
rect 19 33 25 34
rect 9 28 11 33
rect 22 23 24 33
rect 29 23 31 41
rect 9 15 11 19
rect 22 12 24 17
rect 29 12 31 17
<< ndiffusion >>
rect 4 25 9 28
rect 2 24 9 25
rect 2 20 3 24
rect 7 20 9 24
rect 2 19 9 20
rect 11 23 20 28
rect 11 19 22 23
rect 13 17 22 19
rect 24 17 29 23
rect 31 22 38 23
rect 31 18 33 22
rect 37 18 38 22
rect 31 17 38 18
rect 13 12 20 17
rect 13 8 14 12
rect 18 8 20 12
rect 13 7 20 8
<< pdiffusion >>
rect 13 68 19 69
rect 13 64 14 68
rect 18 64 19 68
rect 13 63 19 64
rect 32 68 38 69
rect 32 64 33 68
rect 37 64 38 68
rect 32 63 38 64
rect 13 60 17 63
rect 4 55 9 60
rect 2 54 9 55
rect 2 50 3 54
rect 7 50 9 54
rect 2 47 9 50
rect 2 43 3 47
rect 7 43 9 47
rect 2 42 9 43
rect 11 56 17 60
rect 33 56 38 63
rect 11 50 19 56
rect 21 55 29 56
rect 21 51 23 55
rect 27 51 29 55
rect 21 50 29 51
rect 31 50 38 56
rect 11 42 17 50
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect -2 68 42 78
rect 14 63 18 64
rect 33 63 37 64
rect 2 54 7 55
rect 2 50 3 54
rect 2 47 7 50
rect 2 43 3 47
rect 2 42 7 43
rect 10 51 23 55
rect 27 51 28 55
rect 2 25 6 42
rect 10 38 14 51
rect 25 42 30 46
rect 34 42 38 55
rect 17 34 20 38
rect 24 34 31 38
rect 10 30 14 34
rect 10 26 22 30
rect 25 26 31 34
rect 2 24 7 25
rect 2 20 3 24
rect 7 20 14 23
rect 2 17 14 20
rect 18 22 22 26
rect 18 18 33 22
rect 37 18 38 22
rect -2 8 14 12
rect 18 8 42 12
rect -2 2 42 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
<< ntransistor >>
rect 9 19 11 28
rect 22 17 24 23
rect 29 17 31 23
<< ptransistor >>
rect 9 42 11 60
rect 19 50 21 56
rect 29 50 31 56
<< polycontact >>
rect 30 42 34 46
rect 10 34 14 38
rect 20 34 24 38
<< ndcontact >>
rect 3 20 7 24
rect 33 18 37 22
rect 14 8 18 12
<< pdcontact >>
rect 14 64 18 68
rect 33 64 37 68
rect 3 50 7 54
rect 3 43 7 47
rect 23 51 27 55
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
<< psubstratepdiff >>
rect 0 2 40 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 40 2
rect 0 -3 40 -2
<< nsubstratendiff >>
rect 0 82 40 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 40 82
rect 0 77 40 78
<< labels >>
rlabel polycontact 12 36 12 36 6 zn
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 20 12 20 6 z
rlabel metal1 12 40 12 40 6 zn
rlabel metal1 20 6 20 6 6 vss
rlabel metal1 20 36 20 36 6 a
rlabel metal1 28 32 28 32 6 a
rlabel metal1 28 44 28 44 6 b
rlabel metal1 19 53 19 53 6 zn
rlabel metal1 20 74 20 74 6 vdd
rlabel metal1 28 20 28 20 6 zn
rlabel metal1 36 52 36 52 6 b
<< end >>
