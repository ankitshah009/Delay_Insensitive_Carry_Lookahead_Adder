magic
tech scmos
timestamp 1179387643
<< checkpaint >>
rect -22 -22 134 94
<< ab >>
rect 0 0 112 72
<< pwell >>
rect -4 -4 116 32
<< nwell >>
rect -4 32 116 76
<< polysilicon >>
rect 9 66 11 70
rect 19 66 21 70
rect 61 66 63 70
rect 71 66 73 70
rect 29 59 31 64
rect 39 59 41 64
rect 48 43 54 44
rect 48 39 49 43
rect 53 39 54 43
rect 48 38 54 39
rect 81 59 83 64
rect 91 59 93 64
rect 9 35 11 38
rect 19 35 21 38
rect 29 35 31 38
rect 39 35 41 38
rect 48 35 50 38
rect 9 34 25 35
rect 9 33 20 34
rect 16 30 20 33
rect 24 30 25 34
rect 29 33 50 35
rect 61 35 63 38
rect 71 35 73 38
rect 81 35 83 38
rect 91 35 93 38
rect 61 34 73 35
rect 61 33 66 34
rect 16 29 25 30
rect 9 24 11 29
rect 16 27 28 29
rect 16 24 18 27
rect 26 24 28 27
rect 33 24 35 33
rect 65 30 66 33
rect 70 33 73 34
rect 78 34 103 35
rect 78 33 98 34
rect 70 30 71 33
rect 65 29 71 30
rect 78 29 80 33
rect 97 30 98 33
rect 102 30 103 34
rect 97 29 103 30
rect 65 24 67 29
rect 75 27 80 29
rect 75 24 77 27
rect 85 26 91 27
rect 9 4 11 12
rect 16 8 18 12
rect 26 8 28 12
rect 33 4 35 12
rect 9 2 35 4
rect 85 22 86 26
rect 90 23 91 26
rect 90 22 97 23
rect 85 21 97 22
rect 85 18 87 21
rect 95 18 97 21
rect 65 2 67 6
rect 75 2 77 6
rect 85 4 87 9
rect 95 4 97 9
<< ndiffusion >>
rect 2 17 9 24
rect 2 13 3 17
rect 7 13 9 17
rect 2 12 9 13
rect 11 12 16 24
rect 18 23 26 24
rect 18 19 20 23
rect 24 19 26 23
rect 18 12 26 19
rect 28 12 33 24
rect 35 12 44 24
rect 37 8 44 12
rect 37 4 38 8
rect 42 4 44 8
rect 37 3 44 4
rect 60 19 65 24
rect 58 18 65 19
rect 58 14 59 18
rect 63 14 65 18
rect 58 13 65 14
rect 60 6 65 13
rect 67 23 75 24
rect 67 19 69 23
rect 73 19 75 23
rect 67 6 75 19
rect 77 18 83 24
rect 77 14 85 18
rect 77 10 79 14
rect 83 10 85 14
rect 77 9 85 10
rect 87 17 95 18
rect 87 13 89 17
rect 93 13 95 17
rect 87 9 95 13
rect 97 9 105 18
rect 77 6 83 9
rect 99 8 105 9
rect 99 4 100 8
rect 104 4 105 8
rect 99 3 105 4
<< pdiffusion >>
rect 4 59 9 66
rect 2 58 9 59
rect 2 54 3 58
rect 7 54 9 58
rect 2 51 9 54
rect 2 47 3 51
rect 7 47 9 51
rect 2 46 9 47
rect 4 38 9 46
rect 11 50 19 66
rect 11 46 13 50
rect 17 46 19 50
rect 11 43 19 46
rect 11 39 13 43
rect 17 39 19 43
rect 11 38 19 39
rect 21 59 26 66
rect 54 65 61 66
rect 54 61 55 65
rect 59 61 61 65
rect 21 58 29 59
rect 21 54 23 58
rect 27 54 29 58
rect 21 38 29 54
rect 31 43 39 59
rect 31 39 33 43
rect 37 39 39 43
rect 31 38 39 39
rect 41 58 48 59
rect 41 54 43 58
rect 47 54 48 58
rect 41 53 48 54
rect 54 58 61 61
rect 54 54 55 58
rect 59 54 61 58
rect 54 53 61 54
rect 41 38 46 53
rect 56 38 61 53
rect 63 57 71 66
rect 63 53 65 57
rect 69 53 71 57
rect 63 50 71 53
rect 63 46 65 50
rect 69 46 71 50
rect 63 38 71 46
rect 73 59 79 66
rect 73 58 81 59
rect 73 54 75 58
rect 79 54 81 58
rect 73 38 81 54
rect 83 43 91 59
rect 83 39 85 43
rect 89 39 91 43
rect 83 38 91 39
rect 93 58 100 59
rect 93 54 95 58
rect 99 54 100 58
rect 93 38 100 54
<< metal1 >>
rect -2 68 114 72
rect -2 65 104 68
rect -2 64 55 65
rect 54 61 55 64
rect 59 64 104 65
rect 108 64 114 68
rect 59 61 60 64
rect 54 58 60 61
rect 74 58 80 64
rect 2 54 3 58
rect 7 54 23 58
rect 27 54 43 58
rect 47 54 48 58
rect 54 54 55 58
rect 59 54 60 58
rect 65 57 69 58
rect 2 51 7 54
rect 2 47 3 51
rect 74 54 75 58
rect 79 54 80 58
rect 94 58 100 64
rect 94 54 95 58
rect 99 54 100 58
rect 65 50 69 53
rect 2 46 7 47
rect 12 46 13 50
rect 17 46 65 50
rect 69 46 110 50
rect 2 26 6 46
rect 12 43 17 46
rect 49 43 53 46
rect 12 39 13 43
rect 12 38 17 39
rect 32 39 33 43
rect 37 39 38 43
rect 32 34 38 39
rect 84 42 85 43
rect 49 38 53 39
rect 57 39 85 42
rect 89 39 90 43
rect 57 38 90 39
rect 57 34 61 38
rect 97 34 103 42
rect 19 30 20 34
rect 24 30 61 34
rect 65 30 66 34
rect 70 30 82 34
rect 89 30 98 34
rect 102 30 103 34
rect 57 26 61 30
rect 78 26 82 30
rect 2 23 24 26
rect 2 22 20 23
rect 57 23 73 26
rect 57 22 69 23
rect 20 18 24 19
rect 78 22 86 26
rect 90 22 91 26
rect 69 18 73 19
rect 3 17 7 18
rect 20 14 59 18
rect 63 14 64 18
rect 106 17 110 46
rect 79 14 83 15
rect 3 8 7 13
rect 88 13 89 17
rect 93 13 110 17
rect 79 8 83 10
rect -2 4 38 8
rect 42 4 49 8
rect 53 4 100 8
rect 104 4 114 8
rect -2 0 114 4
<< ntransistor >>
rect 9 12 11 24
rect 16 12 18 24
rect 26 12 28 24
rect 33 12 35 24
rect 65 6 67 24
rect 75 6 77 24
rect 85 9 87 18
rect 95 9 97 18
<< ptransistor >>
rect 9 38 11 66
rect 19 38 21 66
rect 29 38 31 59
rect 39 38 41 59
rect 61 38 63 66
rect 71 38 73 66
rect 81 38 83 59
rect 91 38 93 59
<< polycontact >>
rect 49 39 53 43
rect 20 30 24 34
rect 66 30 70 34
rect 98 30 102 34
rect 86 22 90 26
<< ndcontact >>
rect 3 13 7 17
rect 20 19 24 23
rect 38 4 42 8
rect 59 14 63 18
rect 69 19 73 23
rect 79 10 83 14
rect 89 13 93 17
rect 100 4 104 8
<< pdcontact >>
rect 3 54 7 58
rect 3 47 7 51
rect 13 46 17 50
rect 13 39 17 43
rect 55 61 59 65
rect 23 54 27 58
rect 33 39 37 43
rect 43 54 47 58
rect 55 54 59 58
rect 65 53 69 57
rect 65 46 69 50
rect 75 54 79 58
rect 85 39 89 43
rect 95 54 99 58
<< psubstratepcontact >>
rect 49 4 53 8
<< nsubstratencontact >>
rect 104 64 108 68
<< psubstratepdiff >>
rect 48 8 54 24
rect 48 4 49 8
rect 53 4 54 8
rect 48 3 54 4
<< nsubstratendiff >>
rect 103 68 109 69
rect 103 64 104 68
rect 108 64 109 68
rect 103 63 109 64
<< labels >>
rlabel polycontact 51 41 51 41 6 bn
rlabel metal1 12 24 12 24 6 z
rlabel metal1 4 40 4 40 6 z
rlabel metal1 14 44 14 44 6 bn
rlabel metal1 12 56 12 56 6 z
rlabel metal1 36 16 36 16 6 z
rlabel metal1 28 16 28 16 6 z
rlabel metal1 20 24 20 24 6 z
rlabel metal1 35 36 35 36 6 an
rlabel metal1 36 56 36 56 6 z
rlabel metal1 28 56 28 56 6 z
rlabel metal1 20 56 20 56 6 z
rlabel metal1 56 4 56 4 6 vss
rlabel ndcontact 60 16 60 16 6 z
rlabel metal1 52 16 52 16 6 z
rlabel metal1 44 16 44 16 6 z
rlabel metal1 40 32 40 32 6 an
rlabel metal1 51 44 51 44 6 bn
rlabel pdcontact 44 56 44 56 6 z
rlabel metal1 56 68 56 68 6 vdd
rlabel ndcontact 71 22 71 22 6 an
rlabel metal1 84 24 84 24 6 b
rlabel metal1 76 32 76 32 6 b
rlabel polycontact 68 32 68 32 6 b
rlabel pdcontact 87 40 87 40 6 an
rlabel metal1 67 52 67 52 6 bn
rlabel metal1 99 15 99 15 6 bn
rlabel metal1 92 32 92 32 6 a
rlabel metal1 100 36 100 36 6 a
rlabel metal1 61 48 61 48 6 bn
<< end >>
