magic
tech scmos
timestamp 1179385815
<< checkpaint >>
rect -22 -25 46 105
<< ab >>
rect 0 0 24 80
<< pwell >>
rect -4 -7 28 36
<< nwell >>
rect -4 36 28 87
<< polysilicon >>
rect 9 60 11 65
rect 9 39 11 42
rect 9 38 16 39
rect 9 34 11 38
rect 15 34 16 38
rect 9 33 16 34
rect 9 30 11 33
rect 9 16 11 21
<< ndiffusion >>
rect 2 29 9 30
rect 2 25 3 29
rect 7 25 9 29
rect 2 24 9 25
rect 4 21 9 24
rect 11 26 19 30
rect 11 22 13 26
rect 17 22 19 26
rect 11 21 19 22
<< pdiffusion >>
rect 13 62 20 63
rect 13 60 14 62
rect 4 55 9 60
rect 2 54 9 55
rect 2 50 3 54
rect 7 50 9 54
rect 2 47 9 50
rect 2 43 3 47
rect 7 43 9 47
rect 2 42 9 43
rect 11 58 14 60
rect 18 58 20 62
rect 11 42 20 58
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect -2 68 26 78
rect 13 62 19 68
rect 13 58 14 62
rect 18 58 19 62
rect 2 54 14 55
rect 2 50 3 54
rect 7 50 14 54
rect 2 49 14 50
rect 2 47 7 49
rect 2 43 3 47
rect 2 42 7 43
rect 2 30 6 42
rect 18 39 22 55
rect 10 38 22 39
rect 10 34 11 38
rect 15 34 22 38
rect 10 33 22 34
rect 2 29 7 30
rect 2 25 3 29
rect 2 24 7 25
rect 13 26 17 27
rect 2 17 6 24
rect 13 12 17 22
rect -2 2 26 12
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
<< ntransistor >>
rect 9 21 11 30
<< ptransistor >>
rect 9 42 11 60
<< polycontact >>
rect 11 34 15 38
<< ndcontact >>
rect 3 25 7 29
rect 13 22 17 26
<< pdcontact >>
rect 3 50 7 54
rect 3 43 7 47
rect 14 58 18 62
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
<< psubstratepdiff >>
rect 0 2 24 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 24 2
rect 0 -3 24 -2
<< nsubstratendiff >>
rect 0 82 24 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 24 82
rect 0 77 24 78
<< labels >>
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 6 12 6 6 vss
rlabel polycontact 12 36 12 36 6 a
rlabel metal1 12 52 12 52 6 z
rlabel metal1 12 74 12 74 6 vdd
rlabel metal1 20 44 20 44 6 a
<< end >>
