magic
tech scmos
timestamp 1185094723
<< checkpaint >>
rect -22 -22 92 122
<< ab >>
rect 0 0 70 100
<< pwell >>
rect -4 -4 74 48
<< nwell >>
rect -4 48 74 104
<< polysilicon >>
rect 15 94 17 98
rect 23 94 25 98
rect 35 94 37 98
rect 43 94 45 98
rect 57 80 59 85
rect 15 53 17 56
rect 8 52 17 53
rect 8 48 9 52
rect 13 50 17 52
rect 13 48 19 50
rect 8 47 19 48
rect 7 42 13 43
rect 7 38 8 42
rect 12 38 13 42
rect 7 37 13 38
rect 11 31 13 37
rect 17 37 19 47
rect 23 43 25 56
rect 35 53 37 56
rect 29 52 37 53
rect 29 48 30 52
rect 34 48 37 52
rect 29 47 37 48
rect 23 42 33 43
rect 23 41 28 42
rect 27 38 28 41
rect 32 38 33 42
rect 27 37 33 38
rect 43 41 45 56
rect 57 53 59 56
rect 51 52 59 53
rect 51 48 52 52
rect 56 48 59 52
rect 51 47 59 48
rect 43 40 52 41
rect 43 37 47 40
rect 17 34 21 37
rect 19 31 21 34
rect 31 31 33 37
rect 39 36 47 37
rect 51 36 52 40
rect 39 35 52 36
rect 39 31 41 35
rect 57 31 59 47
rect 57 14 59 19
rect 11 9 13 14
rect 19 9 21 14
rect 31 9 33 14
rect 39 9 41 14
<< ndiffusion >>
rect 3 14 11 31
rect 13 14 19 31
rect 21 22 31 31
rect 21 18 24 22
rect 28 18 31 22
rect 21 14 31 18
rect 33 14 39 31
rect 41 30 57 31
rect 41 26 48 30
rect 52 26 57 30
rect 41 22 57 26
rect 41 18 48 22
rect 52 19 57 22
rect 59 30 67 31
rect 59 26 62 30
rect 66 26 67 30
rect 59 25 67 26
rect 59 19 64 25
rect 52 18 55 19
rect 41 14 55 18
rect 3 11 9 14
rect 3 7 4 11
rect 8 7 9 11
rect 3 6 9 7
<< pdiffusion >>
rect 6 92 15 94
rect 6 88 8 92
rect 12 88 15 92
rect 6 82 15 88
rect 6 78 8 82
rect 12 78 15 82
rect 6 56 15 78
rect 17 56 23 94
rect 25 62 35 94
rect 25 58 28 62
rect 32 58 35 62
rect 25 56 35 58
rect 37 56 43 94
rect 45 92 55 94
rect 45 88 48 92
rect 52 88 55 92
rect 45 82 55 88
rect 45 78 48 82
rect 52 80 55 82
rect 52 78 57 80
rect 45 56 57 78
rect 59 70 64 80
rect 59 69 67 70
rect 59 65 62 69
rect 66 65 67 69
rect 59 61 67 65
rect 59 57 62 61
rect 66 57 67 61
rect 59 56 67 57
<< metal1 >>
rect -2 96 72 100
rect -2 92 62 96
rect 66 92 72 96
rect -2 88 8 92
rect 12 88 48 92
rect 52 88 72 92
rect 8 82 12 88
rect 8 77 12 78
rect 48 82 52 88
rect 48 77 52 78
rect 7 68 53 72
rect 7 52 13 68
rect 7 48 9 52
rect 7 47 13 48
rect 18 53 22 63
rect 28 62 42 63
rect 32 58 42 62
rect 28 57 42 58
rect 18 52 34 53
rect 18 48 30 52
rect 18 47 34 48
rect 18 43 22 47
rect 7 42 22 43
rect 7 38 8 42
rect 12 38 22 42
rect 7 37 22 38
rect 27 42 33 43
rect 27 38 28 42
rect 32 38 33 42
rect 27 32 33 38
rect 7 28 33 32
rect 7 18 13 28
rect 38 22 42 57
rect 47 53 53 68
rect 62 69 66 70
rect 62 61 66 65
rect 47 52 57 53
rect 47 48 52 52
rect 56 48 57 52
rect 47 47 57 48
rect 62 40 66 57
rect 46 36 47 40
rect 51 36 66 40
rect 23 18 24 22
rect 28 18 42 22
rect 23 17 42 18
rect 48 30 52 31
rect 48 22 52 26
rect 62 30 66 36
rect 62 25 66 26
rect 48 12 52 18
rect -2 11 72 12
rect -2 7 4 11
rect 8 8 72 11
rect 8 7 62 8
rect -2 4 62 7
rect 66 4 72 8
rect -2 0 72 4
<< ntransistor >>
rect 11 14 13 31
rect 19 14 21 31
rect 31 14 33 31
rect 39 14 41 31
rect 57 19 59 31
<< ptransistor >>
rect 15 56 17 94
rect 23 56 25 94
rect 35 56 37 94
rect 43 56 45 94
rect 57 56 59 80
<< polycontact >>
rect 9 48 13 52
rect 8 38 12 42
rect 30 48 34 52
rect 28 38 32 42
rect 52 48 56 52
rect 47 36 51 40
<< ndcontact >>
rect 24 18 28 22
rect 48 26 52 30
rect 48 18 52 22
rect 62 26 66 30
rect 4 7 8 11
<< pdcontact >>
rect 8 88 12 92
rect 8 78 12 82
rect 28 58 32 62
rect 48 88 52 92
rect 48 78 52 82
rect 62 65 66 69
rect 62 57 66 61
<< psubstratepcontact >>
rect 62 4 66 8
<< nsubstratencontact >>
rect 62 92 66 96
<< psubstratepdiff >>
rect 61 8 67 9
rect 61 4 62 8
rect 66 4 67 8
rect 61 3 67 4
<< nsubstratendiff >>
rect 61 96 67 97
rect 61 92 62 96
rect 66 92 67 96
rect 61 91 67 92
<< labels >>
rlabel polysilicon 47 38 47 38 6 sn
rlabel metal1 10 25 10 25 6 a0
rlabel metal1 20 30 20 30 6 a0
rlabel polycontact 10 40 10 40 6 a1
rlabel metal1 20 50 20 50 6 a1
rlabel metal1 10 60 10 60 6 s
rlabel metal1 20 70 20 70 6 s
rlabel metal1 35 6 35 6 6 vss
rlabel metal1 30 20 30 20 6 z
rlabel metal1 30 35 30 35 6 a0
rlabel metal1 30 50 30 50 6 a1
rlabel pdcontact 30 60 30 60 6 z
rlabel metal1 30 70 30 70 6 s
rlabel metal1 35 94 35 94 6 vdd
rlabel metal1 40 40 40 40 6 z
rlabel metal1 50 60 50 60 6 s
rlabel metal1 40 70 40 70 6 s
rlabel metal1 56 38 56 38 6 sn
rlabel metal1 64 47 64 47 6 sn
<< end >>
