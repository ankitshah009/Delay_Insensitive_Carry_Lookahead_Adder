magic
tech scmos
timestamp 1179387535
<< checkpaint >>
rect -22 -22 94 94
<< ab >>
rect 0 0 72 72
<< pwell >>
rect -4 -4 76 32
<< nwell >>
rect -4 32 76 76
<< polysilicon >>
rect 9 50 11 55
rect 41 68 63 70
rect 21 58 27 59
rect 21 54 22 58
rect 26 54 27 58
rect 21 53 27 54
rect 31 58 37 59
rect 31 54 32 58
rect 36 54 37 58
rect 31 53 37 54
rect 21 50 23 53
rect 31 50 33 53
rect 41 50 43 68
rect 61 59 63 68
rect 51 50 53 55
rect 9 34 11 38
rect 9 33 15 34
rect 9 29 10 33
rect 14 29 15 33
rect 21 31 23 38
rect 31 35 33 38
rect 31 33 37 35
rect 41 34 43 38
rect 51 35 53 38
rect 61 35 63 47
rect 48 34 54 35
rect 9 28 15 29
rect 19 28 23 31
rect 35 30 37 33
rect 48 30 49 34
rect 53 30 54 34
rect 9 25 11 28
rect 19 25 21 28
rect 29 25 31 29
rect 35 28 41 30
rect 48 29 54 30
rect 58 34 64 35
rect 58 30 59 34
rect 63 30 64 34
rect 58 29 64 30
rect 39 25 41 28
rect 50 26 52 29
rect 9 14 11 19
rect 19 14 21 19
rect 29 4 31 19
rect 39 14 41 19
rect 50 15 52 20
rect 61 19 63 29
rect 61 4 63 13
rect 29 2 63 4
<< ndiffusion >>
rect 43 25 50 26
rect 2 24 9 25
rect 2 20 3 24
rect 7 20 9 24
rect 2 19 9 20
rect 11 19 19 25
rect 21 24 29 25
rect 21 20 23 24
rect 27 20 29 24
rect 21 19 29 20
rect 31 24 39 25
rect 31 20 33 24
rect 37 20 39 24
rect 31 19 39 20
rect 41 21 44 25
rect 48 21 50 25
rect 41 20 50 21
rect 52 20 59 26
rect 41 19 46 20
rect 13 9 17 19
rect 11 8 17 9
rect 11 4 12 8
rect 16 4 17 8
rect 11 3 17 4
rect 54 19 59 20
rect 54 13 61 19
rect 63 18 70 19
rect 63 14 65 18
rect 69 14 70 18
rect 63 13 70 14
rect 54 12 59 13
rect 53 11 59 12
rect 53 7 54 11
rect 58 7 59 11
rect 53 6 59 7
<< pdiffusion >>
rect 13 68 19 69
rect 13 64 14 68
rect 18 64 19 68
rect 13 50 19 64
rect 53 65 59 66
rect 53 61 54 65
rect 58 61 59 65
rect 53 59 59 61
rect 53 57 61 59
rect 55 50 61 57
rect 4 44 9 50
rect 2 43 9 44
rect 2 39 3 43
rect 7 39 9 43
rect 2 38 9 39
rect 11 38 21 50
rect 23 49 31 50
rect 23 45 25 49
rect 29 45 31 49
rect 23 38 31 45
rect 33 43 41 50
rect 33 39 35 43
rect 39 39 41 43
rect 33 38 41 39
rect 43 43 51 50
rect 43 39 45 43
rect 49 39 51 43
rect 43 38 51 39
rect 53 47 61 50
rect 63 58 70 59
rect 63 54 65 58
rect 69 54 70 58
rect 63 53 70 54
rect 63 47 68 53
rect 53 38 59 47
<< metal1 >>
rect -2 68 74 72
rect -2 64 4 68
rect 8 64 14 68
rect 18 64 29 68
rect 33 65 74 68
rect 33 64 54 65
rect 53 61 54 64
rect 58 64 74 65
rect 58 61 59 64
rect 9 54 22 58
rect 26 54 27 58
rect 31 54 32 58
rect 36 54 65 58
rect 69 54 70 58
rect 18 45 22 54
rect 25 49 56 51
rect 29 47 56 49
rect 2 39 3 43
rect 7 39 14 43
rect 2 37 14 39
rect 2 25 6 37
rect 9 29 10 33
rect 14 29 16 33
rect 2 24 7 25
rect 2 20 3 24
rect 2 19 7 20
rect 12 17 16 29
rect 25 24 29 45
rect 22 20 23 24
rect 27 20 29 24
rect 33 43 39 44
rect 33 39 35 43
rect 33 38 39 39
rect 42 43 49 44
rect 42 39 45 43
rect 42 38 49 39
rect 33 24 37 38
rect 42 25 46 38
rect 52 35 56 47
rect 49 34 56 35
rect 53 30 56 34
rect 49 29 56 30
rect 59 34 63 35
rect 59 26 63 30
rect 42 21 44 25
rect 48 21 49 25
rect 57 22 63 26
rect 33 17 37 20
rect 57 18 61 22
rect 66 19 70 54
rect 12 13 37 17
rect 49 14 61 18
rect 65 18 70 19
rect 69 14 70 18
rect 65 13 70 14
rect 53 8 54 11
rect -2 4 12 8
rect 16 4 22 8
rect 26 7 54 8
rect 58 8 59 11
rect 58 7 74 8
rect 26 4 74 7
rect -2 0 74 4
<< ntransistor >>
rect 9 19 11 25
rect 19 19 21 25
rect 29 19 31 25
rect 39 19 41 25
rect 50 20 52 26
rect 61 13 63 19
<< ptransistor >>
rect 9 38 11 50
rect 21 38 23 50
rect 31 38 33 50
rect 41 38 43 50
rect 51 38 53 50
rect 61 47 63 59
<< polycontact >>
rect 22 54 26 58
rect 32 54 36 58
rect 10 29 14 33
rect 49 30 53 34
rect 59 30 63 34
<< ndcontact >>
rect 3 20 7 24
rect 23 20 27 24
rect 33 20 37 24
rect 44 21 48 25
rect 12 4 16 8
rect 65 14 69 18
rect 54 7 58 11
<< pdcontact >>
rect 14 64 18 68
rect 54 61 58 65
rect 3 39 7 43
rect 25 45 29 49
rect 35 39 39 43
rect 45 39 49 43
rect 65 54 69 58
<< psubstratepcontact >>
rect 22 4 26 8
<< nsubstratencontact >>
rect 4 64 8 68
rect 29 64 33 68
<< psubstratepdiff >>
rect 21 8 27 9
rect 21 4 22 8
rect 26 4 27 8
rect 21 3 27 4
<< nsubstratendiff >>
rect 3 68 9 69
rect 3 64 4 68
rect 8 64 9 68
rect 3 63 9 64
rect 28 68 34 69
rect 28 64 29 68
rect 33 64 34 68
rect 28 63 34 64
<< labels >>
rlabel polycontact 12 31 12 31 6 zn
rlabel polycontact 34 56 34 56 6 bn
rlabel polycontact 51 32 51 32 6 an
rlabel polycontact 12 31 12 31 6 zn
rlabel metal1 4 32 4 32 6 z
rlabel metal1 12 40 12 40 6 z
rlabel metal1 12 56 12 56 6 a
rlabel metal1 27 35 27 35 6 an
rlabel metal1 20 52 20 52 6 a
rlabel metal1 36 4 36 4 6 vss
rlabel metal1 52 16 52 16 6 b
rlabel metal1 45 41 45 41 6 ai
rlabel metal1 44 32 44 32 6 ai
rlabel metal1 35 28 35 28 6 zn
rlabel metal1 36 68 36 68 6 vdd
rlabel metal1 60 24 60 24 6 b
rlabel metal1 54 40 54 40 6 an
rlabel metal1 50 56 50 56 6 bn
rlabel metal1 68 35 68 35 6 bn
<< end >>
