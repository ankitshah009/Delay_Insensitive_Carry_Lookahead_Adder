magic
tech scmos
timestamp 1183911780
<< checkpaint >>
rect -22 -22 102 94
<< ab >>
rect 0 0 80 72
<< pwell >>
rect -4 -4 84 32
<< nwell >>
rect -4 32 84 76
<< polysilicon >>
rect 42 68 71 70
rect 9 56 11 61
rect 35 60 37 65
rect 42 60 44 68
rect 52 60 54 64
rect 59 60 61 64
rect 69 60 71 68
rect 19 50 21 55
rect 35 51 37 54
rect 31 50 37 51
rect 31 46 32 50
rect 36 46 37 50
rect 31 45 37 46
rect 9 35 11 38
rect 19 35 21 38
rect 9 34 31 35
rect 9 33 26 34
rect 10 16 12 33
rect 24 30 26 33
rect 30 30 31 34
rect 24 29 31 30
rect 24 26 26 29
rect 35 20 37 45
rect 42 35 44 54
rect 52 45 54 48
rect 48 44 54 45
rect 48 40 49 44
rect 53 40 54 44
rect 59 43 61 48
rect 48 39 54 40
rect 58 42 64 43
rect 58 38 59 42
rect 63 38 64 42
rect 58 37 64 38
rect 42 33 54 35
rect 41 28 47 29
rect 41 24 42 28
rect 46 24 47 28
rect 41 23 47 24
rect 42 20 44 23
rect 52 20 54 33
rect 59 20 61 37
rect 69 33 71 48
rect 65 32 71 33
rect 65 28 66 32
rect 70 28 71 32
rect 65 27 71 28
rect 69 24 71 27
rect 24 15 26 20
rect 35 9 37 14
rect 42 9 44 14
rect 52 9 54 14
rect 59 9 61 14
rect 69 13 71 18
rect 10 2 12 7
<< ndiffusion >>
rect 2 17 8 18
rect 2 13 3 17
rect 7 16 8 17
rect 17 25 24 26
rect 17 21 18 25
rect 22 21 24 25
rect 17 20 24 21
rect 26 25 33 26
rect 26 21 28 25
rect 32 21 33 25
rect 26 20 33 21
rect 63 20 69 24
rect 7 13 10 16
rect 2 12 10 13
rect 5 7 10 12
rect 12 12 19 16
rect 28 14 35 20
rect 37 14 42 20
rect 44 19 52 20
rect 44 15 46 19
rect 50 15 52 19
rect 44 14 52 15
rect 54 14 59 20
rect 61 18 69 20
rect 71 23 78 24
rect 71 19 73 23
rect 77 19 78 23
rect 71 18 78 19
rect 61 14 67 18
rect 12 8 14 12
rect 18 8 19 12
rect 63 11 67 14
rect 12 7 19 8
rect 63 8 69 11
rect 63 4 64 8
rect 68 4 69 8
rect 63 3 69 4
<< pdiffusion >>
rect 28 59 35 60
rect 4 51 9 56
rect 2 50 9 51
rect 2 46 3 50
rect 7 46 9 50
rect 2 43 9 46
rect 2 39 3 43
rect 7 39 9 43
rect 2 38 9 39
rect 11 50 17 56
rect 28 55 29 59
rect 33 55 35 59
rect 28 54 35 55
rect 37 54 42 60
rect 44 59 52 60
rect 44 55 46 59
rect 50 55 52 59
rect 44 54 52 55
rect 11 49 19 50
rect 11 45 13 49
rect 17 45 19 49
rect 11 38 19 45
rect 21 49 28 50
rect 21 45 23 49
rect 27 45 28 49
rect 21 44 28 45
rect 21 38 26 44
rect 47 48 52 54
rect 54 48 59 60
rect 61 59 69 60
rect 61 55 63 59
rect 67 55 69 59
rect 61 48 69 55
rect 71 54 76 60
rect 71 53 78 54
rect 71 49 73 53
rect 77 49 78 53
rect 71 48 78 49
<< metal1 >>
rect -2 68 82 72
rect -2 64 4 68
rect 8 64 12 68
rect 16 64 82 68
rect 2 50 7 51
rect 2 46 3 50
rect 2 43 7 46
rect 12 49 18 64
rect 29 59 33 64
rect 63 59 67 64
rect 29 54 33 55
rect 41 55 46 59
rect 50 55 51 59
rect 12 45 13 49
rect 17 45 18 49
rect 23 49 32 50
rect 27 46 32 49
rect 36 46 37 50
rect 2 39 3 43
rect 23 42 27 45
rect 41 42 45 55
rect 63 54 67 55
rect 73 53 77 54
rect 2 38 7 39
rect 18 38 27 42
rect 35 38 45 42
rect 49 49 73 50
rect 77 49 78 50
rect 49 46 78 49
rect 49 44 53 46
rect 2 27 6 38
rect 2 21 14 27
rect 18 25 22 38
rect 35 34 39 38
rect 49 34 53 40
rect 25 30 26 34
rect 30 30 39 34
rect 2 17 8 21
rect 18 20 22 21
rect 28 25 32 26
rect 2 13 3 17
rect 7 13 8 17
rect 14 12 18 13
rect 28 8 32 21
rect 35 19 39 30
rect 42 30 53 34
rect 58 42 63 43
rect 58 38 59 42
rect 58 37 63 38
rect 42 28 46 30
rect 58 26 62 37
rect 42 23 46 24
rect 49 22 62 26
rect 66 32 70 33
rect 35 15 46 19
rect 50 15 51 19
rect 66 18 70 28
rect 74 24 78 46
rect 73 23 78 24
rect 77 19 78 23
rect 73 18 78 19
rect 57 14 70 18
rect -2 4 24 8
rect 28 4 64 8
rect 68 4 82 8
rect -2 0 82 4
<< ntransistor >>
rect 24 20 26 26
rect 10 7 12 16
rect 35 14 37 20
rect 42 14 44 20
rect 52 14 54 20
rect 59 14 61 20
rect 69 18 71 24
<< ptransistor >>
rect 9 38 11 56
rect 35 54 37 60
rect 42 54 44 60
rect 19 38 21 50
rect 52 48 54 60
rect 59 48 61 60
rect 69 48 71 60
<< polycontact >>
rect 32 46 36 50
rect 26 30 30 34
rect 49 40 53 44
rect 59 38 63 42
rect 42 24 46 28
rect 66 28 70 32
<< ndcontact >>
rect 3 13 7 17
rect 18 21 22 25
rect 28 21 32 25
rect 46 15 50 19
rect 73 19 77 23
rect 14 8 18 12
rect 64 4 68 8
<< pdcontact >>
rect 3 46 7 50
rect 3 39 7 43
rect 29 55 33 59
rect 46 55 50 59
rect 13 45 17 49
rect 23 45 27 49
rect 63 55 67 59
rect 73 49 77 53
<< psubstratepcontact >>
rect 24 4 28 8
<< nsubstratencontact >>
rect 4 64 8 68
rect 12 64 16 68
<< psubstratepdiff >>
rect 23 8 29 9
rect 23 4 24 8
rect 28 4 29 8
rect 23 3 29 4
<< nsubstratendiff >>
rect 3 68 17 69
rect 3 64 4 68
rect 8 64 12 68
rect 16 64 17 68
rect 3 63 17 64
<< labels >>
rlabel polycontact 44 26 44 26 6 en
rlabel polycontact 27 32 27 32 6 n1
rlabel polycontact 34 48 34 48 6 n2
rlabel polycontact 51 42 51 42 6 en
rlabel metal1 4 32 4 32 6 z
rlabel metal1 12 24 12 24 6 z
rlabel metal1 32 32 32 32 6 n1
rlabel metal1 25 44 25 44 6 n2
rlabel metal1 20 31 20 31 6 n2
rlabel metal1 30 48 30 48 6 n2
rlabel metal1 40 4 40 4 6 vss
rlabel metal1 43 17 43 17 6 n1
rlabel metal1 44 28 44 28 6 en
rlabel metal1 52 24 52 24 6 d
rlabel metal1 51 40 51 40 6 en
rlabel metal1 46 57 46 57 6 n1
rlabel metal1 40 68 40 68 6 vdd
rlabel metal1 60 16 60 16 6 e
rlabel metal1 68 24 68 24 6 e
rlabel metal1 60 36 60 36 6 d
rlabel metal1 76 34 76 34 6 en
rlabel pdcontact 75 50 75 50 6 en
<< end >>
