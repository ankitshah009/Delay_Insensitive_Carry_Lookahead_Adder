magic
tech scmos
timestamp 1179387100
<< checkpaint >>
rect -22 -25 94 105
<< ab >>
rect 0 0 72 80
<< pwell >>
rect -4 -7 76 36
<< nwell >>
rect -4 36 76 87
<< polysilicon >>
rect 11 67 13 72
rect 18 67 20 72
rect 28 67 30 72
rect 35 67 37 72
rect 47 66 49 71
rect 57 66 59 71
rect 11 48 13 51
rect 3 47 13 48
rect 3 43 4 47
rect 8 46 13 47
rect 8 43 9 46
rect 3 42 9 43
rect 18 41 20 51
rect 28 47 30 51
rect 35 48 37 51
rect 47 48 49 53
rect 57 50 59 53
rect 57 49 64 50
rect 35 47 53 48
rect 13 39 20 41
rect 25 46 31 47
rect 25 42 26 46
rect 30 42 31 46
rect 25 41 31 42
rect 35 46 48 47
rect 13 38 15 39
rect 9 37 15 38
rect 9 33 10 37
rect 14 33 15 37
rect 25 35 27 41
rect 35 35 37 46
rect 47 43 48 46
rect 52 43 53 47
rect 57 45 59 49
rect 63 45 64 49
rect 57 44 64 45
rect 47 42 53 43
rect 51 39 53 42
rect 9 32 15 33
rect 13 29 15 32
rect 23 32 27 35
rect 33 32 37 35
rect 41 37 47 38
rect 51 37 56 39
rect 41 33 42 37
rect 46 33 47 37
rect 41 32 47 33
rect 23 29 25 32
rect 33 29 35 32
rect 43 29 45 32
rect 54 29 56 37
rect 61 29 63 44
rect 13 17 15 22
rect 23 17 25 22
rect 33 17 35 22
rect 43 17 45 22
rect 54 13 56 18
rect 61 13 63 18
<< ndiffusion >>
rect 4 22 13 29
rect 15 27 23 29
rect 15 23 17 27
rect 21 23 23 27
rect 15 22 23 23
rect 25 28 33 29
rect 25 24 27 28
rect 31 24 33 28
rect 25 22 33 24
rect 35 27 43 29
rect 35 23 37 27
rect 41 23 43 27
rect 35 22 43 23
rect 45 23 54 29
rect 45 22 48 23
rect 4 12 11 22
rect 47 19 48 22
rect 52 19 54 23
rect 47 18 54 19
rect 56 18 61 29
rect 63 28 70 29
rect 63 24 65 28
rect 69 24 70 28
rect 63 23 70 24
rect 63 18 68 23
rect 4 8 6 12
rect 10 8 11 12
rect 4 7 11 8
<< pdiffusion >>
rect 39 72 45 73
rect 39 68 40 72
rect 44 68 45 72
rect 61 72 68 73
rect 39 67 45 68
rect 2 66 11 67
rect 2 62 3 66
rect 7 62 11 66
rect 2 59 11 62
rect 2 55 3 59
rect 7 55 11 59
rect 2 51 11 55
rect 13 51 18 67
rect 20 56 28 67
rect 20 52 22 56
rect 26 52 28 56
rect 20 51 28 52
rect 30 51 35 67
rect 37 66 45 67
rect 61 68 62 72
rect 66 68 68 72
rect 61 66 68 68
rect 37 53 47 66
rect 49 63 57 66
rect 49 59 51 63
rect 55 59 57 63
rect 49 53 57 59
rect 59 53 68 66
rect 37 51 45 53
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect -2 72 74 78
rect -2 68 40 72
rect 44 68 62 72
rect 66 68 74 72
rect 3 66 7 68
rect 3 59 7 62
rect 3 54 7 55
rect 10 59 51 63
rect 55 59 70 63
rect 10 47 14 59
rect 3 43 4 47
rect 8 43 14 47
rect 10 37 14 39
rect 18 37 22 56
rect 26 52 27 56
rect 33 50 63 54
rect 33 47 38 50
rect 59 49 63 50
rect 26 46 38 47
rect 30 42 38 46
rect 26 41 38 42
rect 47 43 48 47
rect 52 46 53 47
rect 52 43 55 46
rect 59 44 63 45
rect 47 41 55 43
rect 51 38 55 41
rect 18 33 32 37
rect 41 33 42 37
rect 46 33 48 37
rect 51 34 63 38
rect 10 31 14 33
rect 2 25 14 31
rect 26 28 32 33
rect 44 30 48 33
rect 66 30 70 59
rect 44 28 70 30
rect 17 27 21 28
rect 2 17 6 25
rect 26 24 27 28
rect 31 24 32 28
rect 37 27 41 28
rect 17 21 21 23
rect 44 26 65 28
rect 64 24 65 26
rect 69 24 70 28
rect 37 21 41 23
rect 17 17 41 21
rect 47 19 48 23
rect 52 19 53 23
rect 47 12 53 19
rect -2 8 6 12
rect 10 8 74 12
rect -2 2 74 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
<< ntransistor >>
rect 13 22 15 29
rect 23 22 25 29
rect 33 22 35 29
rect 43 22 45 29
rect 54 18 56 29
rect 61 18 63 29
<< ptransistor >>
rect 11 51 13 67
rect 18 51 20 67
rect 28 51 30 67
rect 35 51 37 67
rect 47 53 49 66
rect 57 53 59 66
<< polycontact >>
rect 4 43 8 47
rect 26 42 30 46
rect 10 33 14 37
rect 48 43 52 47
rect 59 45 63 49
rect 42 33 46 37
<< ndcontact >>
rect 17 23 21 27
rect 27 24 31 28
rect 37 23 41 27
rect 48 19 52 23
rect 65 24 69 28
rect 6 8 10 12
<< pdcontact >>
rect 40 68 44 72
rect 3 62 7 66
rect 3 55 7 59
rect 22 52 26 56
rect 62 68 66 72
rect 51 59 55 63
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
<< psubstratepdiff >>
rect 0 2 72 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 72 2
rect 0 -3 72 -2
<< nsubstratendiff >>
rect 0 82 72 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 72 82
rect 0 77 72 78
<< labels >>
rlabel polycontact 6 45 6 45 6 b
rlabel metal1 4 24 4 24 6 a3
rlabel metal1 19 22 19 22 6 n4
rlabel metal1 12 32 12 32 6 a3
rlabel metal1 8 45 8 45 6 b
rlabel metal1 20 44 20 44 6 z
rlabel metal1 36 6 36 6 6 vss
rlabel metal1 28 28 28 28 6 z
rlabel metal1 39 22 39 22 6 n4
rlabel polycontact 28 44 28 44 6 b2
rlabel metal1 36 48 36 48 6 b2
rlabel metal1 36 74 36 74 6 vdd
rlabel metal1 52 44 52 44 6 b1
rlabel metal1 52 52 52 52 6 b2
rlabel metal1 44 52 44 52 6 b2
rlabel metal1 60 36 60 36 6 b1
rlabel metal1 60 52 60 52 6 b2
rlabel metal1 68 43 68 43 6 b
rlabel metal1 40 61 40 61 6 b
<< end >>
