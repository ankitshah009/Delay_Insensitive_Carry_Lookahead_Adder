.subckt iv1v0x8 a vdd vss z
*   SPICE3 file   created from iv1v0x8.ext -      technology: scmos
m00 z      a      vdd    vdd p w=28u  l=2.3636u ad=176p     pd=50u      as=196p     ps=70u
m01 vdd    a      z      vdd p w=28u  l=2.3636u ad=196p     pd=70u      as=176p     ps=50u
m02 z      a      vdd    vdd p w=28u  l=2.3636u ad=176p     pd=50u      as=196p     ps=70u
m03 vdd    a      z      vdd p w=28u  l=2.3636u ad=196p     pd=70u      as=176p     ps=50u
m04 z      a      vss    vss n w=20u  l=2.3636u ad=136p     pd=42u      as=140p     ps=54u
m05 vss    a      z      vss n w=20u  l=2.3636u ad=140p     pd=54u      as=136p     ps=42u
m06 z      a      vss    vss n w=20u  l=2.3636u ad=136p     pd=42u      as=140p     ps=54u
m07 vss    a      z      vss n w=20u  l=2.3636u ad=140p     pd=54u      as=136p     ps=42u
C0  vss    a      0.136f
C1  z      vdd    0.246f
C2  vss    z      0.274f
C3  z      a      0.434f
C4  vss    vdd    0.013f
C5  a      vdd    0.428f
C7  z      vss    0.010f
C8  a      vss    0.186f
.ends
