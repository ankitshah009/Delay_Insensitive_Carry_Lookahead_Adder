magic
tech scmos
timestamp 1180600808
<< checkpaint >>
rect -22 -22 132 122
<< ab >>
rect 0 0 110 100
<< pwell >>
rect -4 -4 114 48
<< nwell >>
rect -4 48 114 104
<< polysilicon >>
rect 35 94 37 98
rect 47 94 49 98
rect 57 94 59 98
rect 81 94 83 98
rect 93 94 95 98
rect 11 84 13 88
rect 23 85 25 89
rect 11 43 13 55
rect 23 53 25 56
rect 35 53 37 56
rect 21 51 25 53
rect 33 51 37 53
rect 21 43 23 51
rect 33 43 35 51
rect 7 42 13 43
rect 7 38 8 42
rect 12 38 13 42
rect 7 37 13 38
rect 17 42 23 43
rect 17 38 18 42
rect 22 38 23 42
rect 17 37 23 38
rect 27 42 35 43
rect 27 38 28 42
rect 32 38 35 42
rect 47 43 49 55
rect 57 43 59 55
rect 81 53 83 56
rect 93 53 95 56
rect 75 52 95 53
rect 75 48 76 52
rect 80 48 95 52
rect 75 47 95 48
rect 47 42 53 43
rect 47 39 48 42
rect 27 37 35 38
rect 11 34 13 37
rect 21 34 23 37
rect 33 34 35 37
rect 45 38 48 39
rect 52 38 53 42
rect 45 37 53 38
rect 57 42 63 43
rect 57 38 58 42
rect 62 38 63 42
rect 57 37 63 38
rect 45 34 47 37
rect 57 34 59 37
rect 81 35 83 47
rect 93 35 95 47
rect 33 18 35 22
rect 45 18 47 22
rect 11 12 13 16
rect 21 13 23 17
rect 57 18 59 22
rect 81 11 83 15
rect 93 11 95 15
<< ndiffusion >>
rect 3 16 11 34
rect 13 17 21 34
rect 23 22 33 34
rect 35 22 45 34
rect 47 22 57 34
rect 59 22 67 34
rect 23 18 26 22
rect 30 18 31 22
rect 37 18 38 22
rect 42 18 43 22
rect 23 17 31 18
rect 37 17 43 18
rect 13 16 18 17
rect 3 12 9 16
rect 49 12 55 22
rect 61 18 62 22
rect 66 18 67 22
rect 61 17 67 18
rect 73 32 81 35
rect 73 28 74 32
rect 78 28 81 32
rect 73 22 81 28
rect 73 18 74 22
rect 78 18 81 22
rect 73 15 81 18
rect 83 32 93 35
rect 83 28 86 32
rect 90 28 93 32
rect 83 22 93 28
rect 83 18 86 22
rect 90 18 93 22
rect 83 15 93 18
rect 95 32 103 35
rect 95 28 98 32
rect 102 28 103 32
rect 95 22 103 28
rect 95 18 98 22
rect 102 18 103 22
rect 95 15 103 18
rect 3 8 4 12
rect 8 8 9 12
rect 3 7 9 8
rect 49 8 50 12
rect 54 8 55 12
rect 49 7 55 8
<< pdiffusion >>
rect 15 92 21 93
rect 15 88 16 92
rect 20 88 21 92
rect 15 85 21 88
rect 28 85 35 94
rect 15 84 23 85
rect 3 82 11 84
rect 3 78 4 82
rect 8 78 11 82
rect 3 55 11 78
rect 13 56 23 84
rect 25 82 35 85
rect 25 78 28 82
rect 32 78 35 82
rect 25 56 35 78
rect 37 72 47 94
rect 37 68 40 72
rect 44 68 47 72
rect 37 56 47 68
rect 13 55 18 56
rect 42 55 47 56
rect 49 55 57 94
rect 59 82 67 94
rect 59 78 62 82
rect 66 78 67 82
rect 59 55 67 78
rect 73 92 81 94
rect 73 88 74 92
rect 78 88 81 92
rect 73 82 81 88
rect 73 78 74 82
rect 78 78 81 82
rect 73 56 81 78
rect 83 82 93 94
rect 83 78 86 82
rect 90 78 93 82
rect 83 72 93 78
rect 83 68 86 72
rect 90 68 93 72
rect 83 62 93 68
rect 83 58 86 62
rect 90 58 93 62
rect 83 56 93 58
rect 95 92 103 94
rect 95 88 98 92
rect 102 88 103 92
rect 95 82 103 88
rect 95 78 98 82
rect 102 78 103 82
rect 95 72 103 78
rect 95 68 98 72
rect 102 68 103 72
rect 95 62 103 68
rect 95 58 98 62
rect 102 58 103 62
rect 95 56 103 58
<< metal1 >>
rect -2 92 112 100
rect -2 88 16 92
rect 20 88 74 92
rect 78 88 98 92
rect 102 88 112 92
rect 74 82 78 88
rect 88 82 92 83
rect 3 78 4 82
rect 8 78 28 82
rect 32 78 62 82
rect 66 78 67 82
rect 85 78 86 82
rect 90 78 92 82
rect 74 77 78 78
rect 8 42 12 73
rect 8 17 12 38
rect 18 42 22 73
rect 18 27 22 38
rect 28 42 32 73
rect 88 72 92 78
rect 28 37 32 38
rect 38 68 40 72
rect 44 68 80 72
rect 85 68 86 72
rect 90 68 92 72
rect 38 32 42 68
rect 28 28 42 32
rect 48 42 52 63
rect 28 22 32 28
rect 48 27 52 38
rect 58 42 62 63
rect 76 52 80 68
rect 88 62 92 68
rect 85 58 86 62
rect 90 58 92 62
rect 76 47 80 48
rect 58 27 62 38
rect 74 32 78 33
rect 88 32 92 58
rect 98 82 102 88
rect 98 72 102 78
rect 98 62 102 68
rect 98 57 102 58
rect 85 28 86 32
rect 90 28 92 32
rect 74 22 78 28
rect 88 22 92 28
rect 25 18 26 22
rect 30 18 32 22
rect 37 18 38 22
rect 42 18 62 22
rect 66 18 67 22
rect 85 18 86 22
rect 90 18 92 22
rect 74 12 78 18
rect 88 17 92 18
rect 98 32 102 33
rect 98 22 102 28
rect 98 12 102 18
rect -2 8 4 12
rect 8 10 50 12
rect 8 8 22 10
rect -2 6 22 8
rect 26 6 30 10
rect 34 6 38 10
rect 42 8 50 10
rect 54 8 112 12
rect 42 6 62 8
rect -2 4 62 6
rect 66 4 74 8
rect 78 4 86 8
rect 90 4 98 8
rect 102 4 112 8
rect -2 0 112 4
<< ntransistor >>
rect 11 16 13 34
rect 21 17 23 34
rect 33 22 35 34
rect 45 22 47 34
rect 57 22 59 34
rect 81 15 83 35
rect 93 15 95 35
<< ptransistor >>
rect 11 55 13 84
rect 23 56 25 85
rect 35 56 37 94
rect 47 55 49 94
rect 57 55 59 94
rect 81 56 83 94
rect 93 56 95 94
<< polycontact >>
rect 8 38 12 42
rect 18 38 22 42
rect 28 38 32 42
rect 76 48 80 52
rect 48 38 52 42
rect 58 38 62 42
<< ndcontact >>
rect 26 18 30 22
rect 38 18 42 22
rect 62 18 66 22
rect 74 28 78 32
rect 74 18 78 22
rect 86 28 90 32
rect 86 18 90 22
rect 98 28 102 32
rect 98 18 102 22
rect 4 8 8 12
rect 50 8 54 12
<< pdcontact >>
rect 16 88 20 92
rect 4 78 8 82
rect 28 78 32 82
rect 40 68 44 72
rect 62 78 66 82
rect 74 88 78 92
rect 74 78 78 82
rect 86 78 90 82
rect 86 68 90 72
rect 86 58 90 62
rect 98 88 102 92
rect 98 78 102 82
rect 98 68 102 72
rect 98 58 102 62
<< psubstratepcontact >>
rect 22 6 26 10
rect 30 6 34 10
rect 38 6 42 10
rect 62 4 66 8
rect 74 4 78 8
rect 86 4 90 8
rect 98 4 102 8
<< psubstratepdiff >>
rect 21 10 43 11
rect 21 6 22 10
rect 26 6 30 10
rect 34 6 38 10
rect 42 6 43 10
rect 61 8 103 9
rect 21 5 43 6
rect 61 4 62 8
rect 66 4 74 8
rect 78 4 86 8
rect 90 4 98 8
rect 102 4 103 8
rect 61 3 103 4
<< labels >>
rlabel metal1 10 45 10 45 6 i0
rlabel metal1 20 50 20 50 6 i1
rlabel metal1 30 55 30 55 6 i4
rlabel metal1 55 6 55 6 6 vss
rlabel metal1 60 45 60 45 6 i3
rlabel metal1 50 45 50 45 6 i2
rlabel metal1 55 94 55 94 6 vdd
rlabel metal1 90 50 90 50 6 q
<< end >>
