magic
tech scmos
timestamp 1179387191
<< checkpaint >>
rect -22 -25 126 105
<< ab >>
rect 0 0 104 80
<< pwell >>
rect -4 -7 108 36
<< nwell >>
rect -4 36 108 87
<< polysilicon >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 66 31 71
rect 39 66 41 71
rect 49 66 51 71
rect 56 66 58 71
rect 66 66 68 71
rect 73 66 75 71
rect 83 60 85 65
rect 90 60 92 65
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 39 39 41 42
rect 49 39 51 42
rect 9 38 41 39
rect 9 37 32 38
rect 9 30 11 37
rect 19 30 21 37
rect 29 34 32 37
rect 36 37 41 38
rect 45 38 51 39
rect 36 34 37 37
rect 29 33 37 34
rect 45 34 46 38
rect 50 34 51 38
rect 45 33 51 34
rect 56 39 58 42
rect 66 39 68 42
rect 56 38 68 39
rect 56 34 63 38
rect 67 34 68 38
rect 56 33 68 34
rect 73 39 75 42
rect 83 39 85 42
rect 90 39 92 42
rect 73 37 85 39
rect 89 38 95 39
rect 29 30 31 33
rect 9 13 11 18
rect 46 28 48 33
rect 56 28 58 33
rect 73 31 75 37
rect 89 34 90 38
rect 94 34 95 38
rect 89 33 95 34
rect 72 30 78 31
rect 72 26 73 30
rect 77 26 78 30
rect 72 25 78 26
rect 19 6 21 10
rect 29 6 31 10
rect 46 6 48 10
rect 56 6 58 10
<< ndiffusion >>
rect 2 29 9 30
rect 2 25 3 29
rect 7 25 9 29
rect 2 24 9 25
rect 4 18 9 24
rect 11 23 19 30
rect 11 19 13 23
rect 17 19 19 23
rect 11 18 19 19
rect 13 10 19 18
rect 21 29 29 30
rect 21 25 23 29
rect 27 25 29 29
rect 21 22 29 25
rect 21 18 23 22
rect 27 18 29 22
rect 21 10 29 18
rect 31 28 44 30
rect 31 16 46 28
rect 31 12 33 16
rect 37 12 46 16
rect 31 10 46 12
rect 48 21 56 28
rect 48 17 50 21
rect 54 17 56 21
rect 48 10 56 17
rect 58 22 65 28
rect 58 18 60 22
rect 64 18 65 22
rect 58 15 65 18
rect 58 11 60 15
rect 64 11 65 15
rect 58 10 65 11
<< pdiffusion >>
rect 2 69 9 70
rect 2 65 3 69
rect 7 65 9 69
rect 2 62 9 65
rect 2 58 3 62
rect 7 58 9 62
rect 2 42 9 58
rect 11 62 19 70
rect 11 58 13 62
rect 17 58 19 62
rect 11 55 19 58
rect 11 51 13 55
rect 17 51 19 55
rect 11 42 19 51
rect 21 66 27 70
rect 21 65 29 66
rect 21 61 23 65
rect 27 61 29 65
rect 21 42 29 61
rect 31 62 39 66
rect 31 58 33 62
rect 37 58 39 62
rect 31 55 39 58
rect 31 51 33 55
rect 37 51 39 55
rect 31 42 39 51
rect 41 65 49 66
rect 41 61 43 65
rect 47 61 49 65
rect 41 57 49 61
rect 41 53 43 57
rect 47 53 49 57
rect 41 42 49 53
rect 51 42 56 66
rect 58 56 66 66
rect 58 52 60 56
rect 64 52 66 56
rect 58 48 66 52
rect 58 44 60 48
rect 64 44 66 48
rect 58 42 66 44
rect 68 42 73 66
rect 75 60 81 66
rect 75 59 83 60
rect 75 55 77 59
rect 81 55 83 59
rect 75 42 83 55
rect 85 42 90 60
rect 92 55 97 60
rect 92 54 99 55
rect 92 50 94 54
rect 98 50 99 54
rect 92 47 99 50
rect 92 43 94 47
rect 98 43 99 47
rect 92 42 99 43
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect -2 69 106 78
rect -2 68 3 69
rect 2 65 3 68
rect 7 68 106 69
rect 7 65 8 68
rect 2 62 8 65
rect 23 65 27 68
rect 2 58 3 62
rect 7 58 8 62
rect 13 62 17 63
rect 43 65 47 68
rect 23 60 27 61
rect 33 62 39 63
rect 13 55 17 58
rect 9 51 13 54
rect 37 58 39 62
rect 33 55 39 58
rect 17 51 33 54
rect 37 51 39 55
rect 43 57 47 61
rect 77 59 81 68
rect 43 52 47 53
rect 60 56 64 57
rect 77 54 81 55
rect 94 54 98 55
rect 9 50 39 51
rect 18 39 22 50
rect 60 48 64 52
rect 2 38 22 39
rect 37 44 60 46
rect 94 47 98 50
rect 64 44 94 46
rect 37 43 94 44
rect 37 42 98 43
rect 37 38 41 42
rect 2 34 27 38
rect 31 34 32 38
rect 36 34 41 38
rect 45 34 46 38
rect 50 34 55 38
rect 62 34 63 38
rect 67 34 90 38
rect 94 34 95 38
rect 2 29 7 34
rect 2 25 3 29
rect 2 24 7 25
rect 23 29 27 34
rect 13 23 17 24
rect 13 12 17 19
rect 23 22 27 25
rect 37 26 41 34
rect 49 30 55 34
rect 49 26 73 30
rect 77 26 78 30
rect 89 26 95 34
rect 37 22 45 26
rect 23 17 27 18
rect 41 21 45 22
rect 41 17 50 21
rect 54 17 55 21
rect 59 18 60 22
rect 64 18 65 22
rect 33 16 37 17
rect 59 15 65 18
rect 74 17 78 26
rect 59 12 60 15
rect -2 11 60 12
rect 64 12 65 15
rect 64 11 106 12
rect -2 2 106 11
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
<< ntransistor >>
rect 9 18 11 30
rect 19 10 21 30
rect 29 10 31 30
rect 46 10 48 28
rect 56 10 58 28
<< ptransistor >>
rect 9 42 11 70
rect 19 42 21 70
rect 29 42 31 66
rect 39 42 41 66
rect 49 42 51 66
rect 56 42 58 66
rect 66 42 68 66
rect 73 42 75 66
rect 83 42 85 60
rect 90 42 92 60
<< polycontact >>
rect 32 34 36 38
rect 46 34 50 38
rect 63 34 67 38
rect 90 34 94 38
rect 73 26 77 30
<< ndcontact >>
rect 3 25 7 29
rect 13 19 17 23
rect 23 25 27 29
rect 23 18 27 22
rect 33 12 37 16
rect 50 17 54 21
rect 60 18 64 22
rect 60 11 64 15
<< pdcontact >>
rect 3 65 7 69
rect 3 58 7 62
rect 13 58 17 62
rect 13 51 17 55
rect 23 61 27 65
rect 33 58 37 62
rect 33 51 37 55
rect 43 61 47 65
rect 43 53 47 57
rect 60 52 64 56
rect 60 44 64 48
rect 77 55 81 59
rect 94 50 98 54
rect 94 43 98 47
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
rect 90 -2 94 2
rect 98 -2 102 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
rect 90 78 94 82
rect 98 78 102 82
<< psubstratepdiff >>
rect 0 2 104 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 104 2
rect 0 -3 104 -2
<< nsubstratendiff >>
rect 0 82 104 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 104 82
rect 0 77 104 78
<< labels >>
rlabel polycontact 33 36 33 36 6 zn
rlabel metal1 4 32 4 32 6 z
rlabel metal1 12 36 12 36 6 z
rlabel metal1 12 52 12 52 6 z
rlabel metal1 20 44 20 44 6 z
rlabel metal1 28 52 28 52 6 z
rlabel metal1 36 56 36 56 6 z
rlabel metal1 52 6 52 6 6 vss
rlabel metal1 48 19 48 19 6 zn
rlabel metal1 60 28 60 28 6 a
rlabel metal1 52 32 52 32 6 a
rlabel metal1 36 36 36 36 6 zn
rlabel metal1 52 74 52 74 6 vdd
rlabel metal1 68 28 68 28 6 a
rlabel metal1 76 20 76 20 6 a
rlabel metal1 68 36 68 36 6 b
rlabel metal1 76 36 76 36 6 b
rlabel metal1 62 49 62 49 6 zn
rlabel metal1 92 32 92 32 6 b
rlabel metal1 84 36 84 36 6 b
rlabel metal1 96 48 96 48 6 zn
<< end >>
