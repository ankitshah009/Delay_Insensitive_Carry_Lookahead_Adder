magic
tech scmos
timestamp 1179386226
<< checkpaint >>
rect -22 -25 62 105
<< ab >>
rect 0 0 40 80
<< pwell >>
rect -4 -7 44 36
<< nwell >>
rect -4 36 44 87
<< polysilicon >>
rect 10 63 16 64
rect 10 59 11 63
rect 15 59 16 63
rect 10 58 16 59
rect 10 56 12 58
rect 9 53 12 56
rect 29 55 31 60
rect 9 50 11 53
rect 19 50 21 54
rect 9 30 11 42
rect 19 39 21 42
rect 16 38 23 39
rect 16 34 18 38
rect 22 34 23 38
rect 16 33 23 34
rect 16 30 18 33
rect 29 31 31 45
rect 28 30 34 31
rect 9 18 11 23
rect 16 18 18 23
rect 28 26 29 30
rect 33 26 34 30
rect 28 25 34 26
rect 28 22 30 25
rect 28 11 30 16
<< ndiffusion >>
rect 2 29 9 30
rect 2 25 3 29
rect 7 25 9 29
rect 2 23 9 25
rect 11 23 16 30
rect 18 23 26 30
rect 20 22 26 23
rect 20 16 28 22
rect 30 21 37 22
rect 30 17 32 21
rect 36 17 37 21
rect 30 16 37 17
rect 20 12 26 16
rect 20 8 21 12
rect 25 8 26 12
rect 20 7 26 8
<< pdiffusion >>
rect 2 72 8 73
rect 2 68 3 72
rect 7 68 8 72
rect 2 58 8 68
rect 21 61 27 62
rect 2 50 7 58
rect 21 57 22 61
rect 26 57 27 61
rect 21 56 27 57
rect 23 55 27 56
rect 23 50 29 55
rect 2 42 9 50
rect 11 47 19 50
rect 11 43 13 47
rect 17 43 19 47
rect 11 42 19 43
rect 21 45 29 50
rect 31 54 38 55
rect 31 50 33 54
rect 37 50 38 54
rect 31 49 38 50
rect 31 45 36 49
rect 21 42 27 45
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect -2 72 42 78
rect -2 68 3 72
rect 7 68 42 72
rect 2 59 11 63
rect 15 59 16 63
rect 2 57 16 59
rect 21 61 27 68
rect 21 57 22 61
rect 26 57 27 61
rect 2 41 6 57
rect 26 50 33 54
rect 37 50 38 54
rect 10 43 13 47
rect 17 43 23 47
rect 10 42 23 43
rect 10 31 14 42
rect 26 39 30 50
rect 2 29 14 31
rect 2 25 3 29
rect 7 25 14 29
rect 18 38 30 39
rect 22 35 30 38
rect 18 21 22 34
rect 34 31 38 47
rect 26 30 38 31
rect 26 26 29 30
rect 33 26 38 30
rect 26 25 38 26
rect 18 17 32 21
rect 36 17 37 21
rect -2 8 21 12
rect 25 8 42 12
rect -2 2 42 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
<< ntransistor >>
rect 9 23 11 30
rect 16 23 18 30
rect 28 16 30 22
<< ptransistor >>
rect 9 42 11 50
rect 19 42 21 50
rect 29 45 31 55
<< polycontact >>
rect 11 59 15 63
rect 18 34 22 38
rect 29 26 33 30
<< ndcontact >>
rect 3 25 7 29
rect 32 17 36 21
rect 21 8 25 12
<< pdcontact >>
rect 3 68 7 72
rect 22 57 26 61
rect 13 43 17 47
rect 33 50 37 54
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
<< psubstratepdiff >>
rect 0 2 40 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 40 2
rect 0 -3 40 -2
<< nsubstratendiff >>
rect 0 82 40 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 40 82
rect 0 77 40 78
<< labels >>
rlabel ptransistor 20 43 20 43 6 an
rlabel ndcontact 4 28 4 28 6 z
rlabel metal1 4 52 4 52 6 b
rlabel metal1 12 36 12 36 6 z
rlabel polycontact 12 60 12 60 6 b
rlabel metal1 20 6 20 6 6 vss
rlabel metal1 20 28 20 28 6 an
rlabel metal1 28 28 28 28 6 a
rlabel metal1 20 44 20 44 6 z
rlabel metal1 20 74 20 74 6 vdd
rlabel metal1 27 19 27 19 6 an
rlabel metal1 36 36 36 36 6 a
rlabel metal1 32 52 32 52 6 an
<< end >>
