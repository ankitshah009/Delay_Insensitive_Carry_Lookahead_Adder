magic
tech scmos
timestamp 1179387207
<< checkpaint >>
rect -22 -25 78 105
<< ab >>
rect 0 0 56 80
<< pwell >>
rect -4 -7 60 36
<< nwell >>
rect -4 36 60 87
<< polysilicon >>
rect 32 70 34 74
rect 39 70 41 74
rect 9 61 11 65
rect 19 61 21 67
rect 9 44 11 47
rect 19 44 21 47
rect 9 43 24 44
rect 9 42 19 43
rect 18 39 19 42
rect 23 39 24 43
rect 48 42 54 43
rect 32 39 34 42
rect 39 39 41 42
rect 48 39 49 42
rect 18 38 24 39
rect 29 38 35 39
rect 9 30 11 35
rect 19 30 21 38
rect 29 34 30 38
rect 34 34 35 38
rect 29 33 35 34
rect 39 38 49 39
rect 53 38 54 42
rect 39 37 54 38
rect 29 25 31 33
rect 39 25 41 37
rect 9 8 11 16
rect 19 12 21 16
rect 29 12 31 17
rect 39 8 41 17
rect 9 6 41 8
<< ndiffusion >>
rect 2 29 9 30
rect 2 25 3 29
rect 7 25 9 29
rect 2 22 9 25
rect 2 18 3 22
rect 7 18 9 22
rect 2 16 9 18
rect 11 29 19 30
rect 11 25 13 29
rect 17 25 19 29
rect 11 22 19 25
rect 11 18 13 22
rect 17 18 19 22
rect 11 16 19 18
rect 21 25 27 30
rect 21 22 29 25
rect 21 18 23 22
rect 27 18 29 22
rect 21 17 29 18
rect 31 24 39 25
rect 31 20 33 24
rect 37 20 39 24
rect 31 17 39 20
rect 41 22 48 25
rect 41 18 43 22
rect 47 18 48 22
rect 41 17 48 18
rect 21 16 27 17
<< pdiffusion >>
rect 23 69 32 70
rect 23 65 24 69
rect 28 65 32 69
rect 23 62 32 65
rect 23 61 24 62
rect 2 60 9 61
rect 2 56 3 60
rect 7 56 9 60
rect 2 53 9 56
rect 2 49 3 53
rect 7 49 9 53
rect 2 47 9 49
rect 11 60 19 61
rect 11 56 13 60
rect 17 56 19 60
rect 11 53 19 56
rect 11 49 13 53
rect 17 49 19 53
rect 11 47 19 49
rect 21 58 24 61
rect 28 58 32 62
rect 21 47 32 58
rect 26 42 32 47
rect 34 42 39 70
rect 41 63 46 70
rect 41 62 48 63
rect 41 58 43 62
rect 47 58 48 62
rect 41 55 48 58
rect 41 51 43 55
rect 47 51 48 55
rect 41 50 48 51
rect 41 42 46 50
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect -2 69 58 78
rect -2 68 24 69
rect 2 60 7 68
rect 23 65 24 68
rect 28 68 58 69
rect 28 65 29 68
rect 23 62 29 65
rect 2 56 3 60
rect 2 53 7 56
rect 13 60 17 61
rect 23 58 24 62
rect 28 58 29 62
rect 43 62 47 63
rect 13 55 17 56
rect 43 55 47 58
rect 2 49 3 53
rect 2 48 7 49
rect 10 53 22 55
rect 10 49 13 53
rect 17 49 22 53
rect 30 51 43 54
rect 30 50 47 51
rect 2 30 6 48
rect 10 30 14 49
rect 30 46 34 50
rect 50 46 54 55
rect 21 43 34 46
rect 18 39 19 43
rect 23 42 34 43
rect 41 42 54 46
rect 23 39 25 42
rect 21 30 25 39
rect 53 41 54 42
rect 29 34 30 38
rect 34 34 46 38
rect 49 37 53 38
rect 2 29 7 30
rect 2 25 3 29
rect 10 29 17 30
rect 10 25 13 29
rect 21 26 37 30
rect 2 22 7 25
rect 2 18 3 22
rect 2 17 7 18
rect 13 22 17 25
rect 33 24 37 26
rect 42 25 46 34
rect 13 17 17 18
rect 22 18 23 22
rect 27 18 28 22
rect 33 18 37 20
rect 42 18 43 22
rect 47 18 48 22
rect 22 12 28 18
rect 42 12 48 18
rect -2 2 58 12
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
<< ntransistor >>
rect 9 16 11 30
rect 19 16 21 30
rect 29 17 31 25
rect 39 17 41 25
<< ptransistor >>
rect 9 47 11 61
rect 19 47 21 61
rect 32 42 34 70
rect 39 42 41 70
<< polycontact >>
rect 19 39 23 43
rect 30 34 34 38
rect 49 38 53 42
<< ndcontact >>
rect 3 25 7 29
rect 3 18 7 22
rect 13 25 17 29
rect 13 18 17 22
rect 23 18 27 22
rect 33 20 37 24
rect 43 18 47 22
<< pdcontact >>
rect 24 65 28 69
rect 3 56 7 60
rect 3 49 7 53
rect 13 56 17 60
rect 13 49 17 53
rect 24 58 28 62
rect 43 58 47 62
rect 43 51 47 55
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
<< psubstratepdiff >>
rect 0 2 56 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 56 2
rect 0 -3 56 -2
<< nsubstratendiff >>
rect 0 82 56 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 56 82
rect 0 77 56 78
<< labels >>
rlabel polysilicon 20 39 20 39 6 zn
rlabel polycontact 21 41 21 41 6 zn
rlabel metal1 12 40 12 40 6 z
rlabel metal1 20 52 20 52 6 z
rlabel metal1 28 6 28 6 6 vss
rlabel metal1 35 24 35 24 6 zn
rlabel metal1 36 36 36 36 6 a
rlabel metal1 28 74 28 74 6 vdd
rlabel metal1 44 28 44 28 6 a
rlabel metal1 44 44 44 44 6 b
rlabel metal1 52 48 52 48 6 b
rlabel metal1 45 56 45 56 6 zn
<< end >>
