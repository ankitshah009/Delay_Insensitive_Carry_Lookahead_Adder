magic
tech scmos
timestamp 1179386930
<< checkpaint >>
rect -22 -22 102 94
<< ab >>
rect 0 0 80 72
<< pwell >>
rect -4 -4 84 32
<< nwell >>
rect -4 32 84 76
<< polysilicon >>
rect 13 64 15 69
rect 20 64 22 69
rect 27 64 29 69
rect 34 64 36 69
rect 44 57 46 61
rect 51 57 53 61
rect 58 57 60 61
rect 65 57 67 61
rect 13 36 15 39
rect 2 35 15 36
rect 2 31 3 35
rect 7 34 15 35
rect 7 31 11 34
rect 2 30 11 31
rect 9 18 11 30
rect 20 29 22 39
rect 27 36 29 39
rect 34 36 36 39
rect 44 36 46 39
rect 27 33 30 36
rect 34 34 46 36
rect 17 28 23 29
rect 17 24 18 28
rect 22 24 23 28
rect 17 23 23 24
rect 28 27 30 33
rect 28 26 34 27
rect 19 18 21 23
rect 28 22 29 26
rect 33 22 34 26
rect 28 21 34 22
rect 31 18 33 21
rect 41 18 43 34
rect 51 27 53 39
rect 58 30 60 39
rect 65 36 67 39
rect 65 35 73 36
rect 65 34 68 35
rect 67 31 68 34
rect 72 31 73 35
rect 67 30 73 31
rect 47 26 53 27
rect 47 22 48 26
rect 52 22 53 26
rect 57 29 63 30
rect 57 25 58 29
rect 62 25 63 29
rect 57 24 63 25
rect 47 21 53 22
rect 57 18 63 19
rect 57 14 58 18
rect 62 14 63 18
rect 57 13 63 14
rect 9 7 11 12
rect 19 7 21 12
rect 31 7 33 12
rect 41 9 43 12
rect 57 9 59 13
rect 41 7 59 9
<< ndiffusion >>
rect 2 17 9 18
rect 2 13 3 17
rect 7 13 9 17
rect 2 12 9 13
rect 11 17 19 18
rect 11 13 13 17
rect 17 13 19 17
rect 11 12 19 13
rect 21 12 31 18
rect 33 17 41 18
rect 33 13 35 17
rect 39 13 41 17
rect 33 12 41 13
rect 43 17 50 18
rect 43 13 45 17
rect 49 13 50 17
rect 43 12 50 13
rect 23 8 29 12
rect 23 4 24 8
rect 28 4 29 8
rect 23 3 29 4
<< pdiffusion >>
rect 4 68 11 69
rect 4 64 6 68
rect 10 64 11 68
rect 4 39 13 64
rect 15 39 20 64
rect 22 39 27 64
rect 29 39 34 64
rect 36 57 41 64
rect 36 50 44 57
rect 36 46 38 50
rect 42 46 44 50
rect 36 39 44 46
rect 46 39 51 57
rect 53 39 58 57
rect 60 39 65 57
rect 67 56 74 57
rect 67 52 69 56
rect 73 52 74 56
rect 67 49 74 52
rect 67 45 69 49
rect 73 45 74 49
rect 67 39 74 45
<< metal1 >>
rect -2 68 82 72
rect -2 64 6 68
rect 10 64 46 68
rect 50 64 68 68
rect 72 64 82 68
rect 2 54 62 58
rect 2 36 6 54
rect 10 46 38 50
rect 42 46 43 50
rect 2 35 7 36
rect 2 31 3 35
rect 2 30 7 31
rect 10 18 14 46
rect 58 42 62 54
rect 68 56 74 64
rect 68 52 69 56
rect 73 52 74 56
rect 68 49 74 52
rect 68 45 69 49
rect 73 45 74 49
rect 18 38 53 42
rect 58 38 73 42
rect 18 28 22 38
rect 49 34 53 38
rect 67 35 73 38
rect 33 26 39 34
rect 49 30 62 34
rect 67 31 68 35
rect 72 31 73 35
rect 58 29 62 30
rect 18 23 22 24
rect 28 22 29 26
rect 33 22 48 26
rect 52 22 53 26
rect 58 24 62 25
rect 66 19 70 27
rect 58 18 70 19
rect 3 17 7 18
rect 10 17 40 18
rect 10 13 13 17
rect 17 13 35 17
rect 39 13 40 17
rect 45 17 49 18
rect 62 14 70 18
rect 58 13 70 14
rect 3 8 7 13
rect 45 8 49 13
rect -2 4 24 8
rect 28 4 68 8
rect 72 4 82 8
rect -2 0 82 4
<< ntransistor >>
rect 9 12 11 18
rect 19 12 21 18
rect 31 12 33 18
rect 41 12 43 18
<< ptransistor >>
rect 13 39 15 64
rect 20 39 22 64
rect 27 39 29 64
rect 34 39 36 64
rect 44 39 46 57
rect 51 39 53 57
rect 58 39 60 57
rect 65 39 67 57
<< polycontact >>
rect 3 31 7 35
rect 18 24 22 28
rect 29 22 33 26
rect 68 31 72 35
rect 48 22 52 26
rect 58 25 62 29
rect 58 14 62 18
<< ndcontact >>
rect 3 13 7 17
rect 13 13 17 17
rect 35 13 39 17
rect 45 13 49 17
rect 24 4 28 8
<< pdcontact >>
rect 6 64 10 68
rect 38 46 42 50
rect 69 52 73 56
rect 69 45 73 49
<< psubstratepcontact >>
rect 68 4 72 8
<< nsubstratencontact >>
rect 46 64 50 68
rect 68 64 72 68
<< psubstratepdiff >>
rect 67 8 73 24
rect 67 4 68 8
rect 72 4 73 8
rect 67 3 73 4
<< nsubstratendiff >>
rect 45 68 73 69
rect 45 64 46 68
rect 50 64 68 68
rect 72 64 73 68
rect 45 63 73 64
<< labels >>
rlabel metal1 4 44 4 44 6 a
rlabel metal1 28 16 28 16 6 z
rlabel metal1 20 16 20 16 6 z
rlabel metal1 20 32 20 32 6 b
rlabel metal1 12 28 12 28 6 z
rlabel metal1 28 40 28 40 6 b
rlabel metal1 28 48 28 48 6 z
rlabel metal1 20 48 20 48 6 z
rlabel metal1 28 56 28 56 6 a
rlabel metal1 20 56 20 56 6 a
rlabel metal1 12 56 12 56 6 a
rlabel metal1 40 4 40 4 6 vss
rlabel ndcontact 36 16 36 16 6 z
rlabel metal1 44 24 44 24 6 c
rlabel metal1 36 28 36 28 6 c
rlabel metal1 44 40 44 40 6 b
rlabel metal1 36 40 36 40 6 b
rlabel metal1 36 48 36 48 6 z
rlabel metal1 44 56 44 56 6 a
rlabel metal1 36 56 36 56 6 a
rlabel metal1 40 68 40 68 6 vdd
rlabel polycontact 60 16 60 16 6 d
rlabel metal1 52 32 52 32 6 b
rlabel metal1 60 48 60 48 6 a
rlabel metal1 52 56 52 56 6 a
rlabel metal1 68 20 68 20 6 d
rlabel metal1 68 40 68 40 6 a
<< end >>
