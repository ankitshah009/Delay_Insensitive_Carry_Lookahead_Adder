magic
tech scmos
timestamp 1179386616
<< checkpaint >>
rect -22 -25 166 105
<< ab >>
rect 0 0 144 80
<< pwell >>
rect -4 -7 148 36
<< nwell >>
rect -4 36 148 87
<< polysilicon >>
rect 20 69 22 74
rect 30 69 32 74
rect 40 69 42 74
rect 50 69 52 74
rect 70 69 72 74
rect 80 69 82 74
rect 100 69 102 74
rect 110 69 112 74
rect 120 69 122 74
rect 20 39 22 42
rect 30 39 32 42
rect 40 39 42 42
rect 10 38 42 39
rect 10 34 11 38
rect 15 34 18 38
rect 22 34 42 38
rect 10 33 42 34
rect 10 30 12 33
rect 20 30 22 33
rect 30 30 32 33
rect 40 30 42 33
rect 50 39 52 42
rect 70 39 72 42
rect 80 39 82 42
rect 100 39 102 42
rect 110 39 112 42
rect 120 39 122 42
rect 50 38 92 39
rect 50 34 51 38
rect 55 34 58 38
rect 62 34 92 38
rect 50 33 92 34
rect 50 30 52 33
rect 60 30 62 33
rect 70 30 72 33
rect 80 30 82 33
rect 90 30 92 33
rect 100 38 132 39
rect 100 34 119 38
rect 123 34 127 38
rect 131 34 132 38
rect 100 33 132 34
rect 100 30 102 33
rect 110 30 112 33
rect 120 30 122 33
rect 130 30 132 33
rect 80 15 82 20
rect 90 15 92 20
rect 10 6 12 10
rect 20 6 22 10
rect 30 6 32 10
rect 40 6 42 10
rect 50 6 52 10
rect 60 6 62 10
rect 70 6 72 10
rect 100 6 102 10
rect 110 6 112 10
rect 120 6 122 10
rect 130 6 132 10
<< ndiffusion >>
rect 3 29 10 30
rect 3 25 4 29
rect 8 25 10 29
rect 3 22 10 25
rect 3 18 4 22
rect 8 18 10 22
rect 3 17 10 18
rect 5 10 10 17
rect 12 22 20 30
rect 12 18 14 22
rect 18 18 20 22
rect 12 15 20 18
rect 12 11 14 15
rect 18 11 20 15
rect 12 10 20 11
rect 22 29 30 30
rect 22 25 24 29
rect 28 25 30 29
rect 22 22 30 25
rect 22 18 24 22
rect 28 18 30 22
rect 22 10 30 18
rect 32 15 40 30
rect 32 11 34 15
rect 38 11 40 15
rect 32 10 40 11
rect 42 22 50 30
rect 42 18 44 22
rect 48 18 50 22
rect 42 10 50 18
rect 52 29 60 30
rect 52 25 54 29
rect 58 25 60 29
rect 52 10 60 25
rect 62 22 70 30
rect 62 18 64 22
rect 68 18 70 22
rect 62 10 70 18
rect 72 29 80 30
rect 72 25 74 29
rect 78 25 80 29
rect 72 20 80 25
rect 82 25 90 30
rect 82 21 84 25
rect 88 21 90 25
rect 82 20 90 21
rect 92 29 100 30
rect 92 25 94 29
rect 98 25 100 29
rect 92 20 100 25
rect 72 10 77 20
rect 95 10 100 20
rect 102 29 110 30
rect 102 25 104 29
rect 108 25 110 29
rect 102 10 110 25
rect 112 21 120 30
rect 112 17 114 21
rect 118 17 120 21
rect 112 10 120 17
rect 122 29 130 30
rect 122 25 124 29
rect 128 25 130 29
rect 122 10 130 25
rect 132 29 139 30
rect 132 25 134 29
rect 138 25 139 29
rect 132 22 139 25
rect 132 18 134 22
rect 138 18 139 22
rect 132 17 139 18
rect 132 10 137 17
<< pdiffusion >>
rect 13 68 20 69
rect 13 64 14 68
rect 18 64 20 68
rect 13 61 20 64
rect 13 57 14 61
rect 18 57 20 61
rect 13 42 20 57
rect 22 54 30 69
rect 22 50 24 54
rect 28 50 30 54
rect 22 47 30 50
rect 22 43 24 47
rect 28 43 30 47
rect 22 42 30 43
rect 32 68 40 69
rect 32 64 34 68
rect 38 64 40 68
rect 32 61 40 64
rect 32 57 34 61
rect 38 57 40 61
rect 32 42 40 57
rect 42 54 50 69
rect 42 50 44 54
rect 48 50 50 54
rect 42 47 50 50
rect 42 43 44 47
rect 48 43 50 47
rect 42 42 50 43
rect 52 68 70 69
rect 52 64 54 68
rect 58 64 64 68
rect 68 64 70 68
rect 52 61 70 64
rect 52 57 54 61
rect 58 57 64 61
rect 68 57 70 61
rect 52 42 70 57
rect 72 54 80 69
rect 72 50 74 54
rect 78 50 80 54
rect 72 47 80 50
rect 72 43 74 47
rect 78 43 80 47
rect 72 42 80 43
rect 82 68 89 69
rect 82 64 84 68
rect 88 64 89 68
rect 82 61 89 64
rect 82 57 84 61
rect 88 57 89 61
rect 82 42 89 57
rect 95 55 100 69
rect 93 54 100 55
rect 93 50 94 54
rect 98 50 100 54
rect 93 47 100 50
rect 93 43 94 47
rect 98 43 100 47
rect 93 42 100 43
rect 102 68 110 69
rect 102 64 104 68
rect 108 64 110 68
rect 102 61 110 64
rect 102 57 104 61
rect 108 57 110 61
rect 102 42 110 57
rect 112 54 120 69
rect 112 50 114 54
rect 118 50 120 54
rect 112 47 120 50
rect 112 43 114 47
rect 118 43 120 47
rect 112 42 120 43
rect 122 68 130 69
rect 122 64 124 68
rect 128 64 130 68
rect 122 61 130 64
rect 122 57 124 61
rect 128 57 130 61
rect 122 42 130 57
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect 118 78 122 82
rect 126 78 130 82
rect 134 78 138 82
rect 142 78 146 82
rect -2 68 146 78
rect 14 61 18 64
rect 14 56 18 57
rect 34 61 38 64
rect 34 56 38 57
rect 54 61 58 64
rect 54 56 58 57
rect 64 61 68 64
rect 64 56 68 57
rect 2 38 6 55
rect 24 54 28 55
rect 24 47 28 50
rect 44 54 48 55
rect 44 47 48 50
rect 28 43 44 46
rect 74 54 78 63
rect 84 61 88 64
rect 84 56 88 57
rect 104 61 108 64
rect 104 56 108 57
rect 124 61 128 64
rect 124 56 128 57
rect 74 47 78 50
rect 48 43 74 46
rect 94 54 98 55
rect 94 47 98 50
rect 78 43 94 46
rect 114 54 118 55
rect 114 47 118 50
rect 98 43 114 46
rect 24 42 118 43
rect 2 34 11 38
rect 15 34 18 38
rect 22 34 23 38
rect 2 33 23 34
rect 41 34 51 38
rect 55 34 58 38
rect 62 34 63 38
rect 4 29 28 30
rect 8 26 24 29
rect 4 22 8 25
rect 41 26 47 34
rect 75 30 98 34
rect 106 30 110 42
rect 129 38 135 46
rect 118 34 119 38
rect 123 34 127 38
rect 131 34 135 38
rect 75 29 79 30
rect 53 25 54 29
rect 58 25 74 29
rect 78 25 79 29
rect 94 29 98 30
rect 84 25 88 26
rect 24 22 28 25
rect 4 17 8 18
rect 13 18 14 22
rect 18 18 19 22
rect 28 18 44 22
rect 48 18 64 22
rect 68 21 84 22
rect 68 18 88 21
rect 103 29 129 30
rect 103 25 104 29
rect 108 25 124 29
rect 128 25 129 29
rect 134 29 138 30
rect 94 21 98 25
rect 134 22 138 25
rect 13 15 19 18
rect 94 17 114 21
rect 118 18 134 21
rect 118 17 138 18
rect 13 12 14 15
rect -2 11 14 12
rect 18 12 19 15
rect 33 12 34 15
rect 18 11 34 12
rect 38 12 39 15
rect 38 11 146 12
rect -2 2 146 11
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 122 2
rect 126 -2 130 2
rect 134 -2 138 2
rect 142 -2 146 2
<< ntransistor >>
rect 10 10 12 30
rect 20 10 22 30
rect 30 10 32 30
rect 40 10 42 30
rect 50 10 52 30
rect 60 10 62 30
rect 70 10 72 30
rect 80 20 82 30
rect 90 20 92 30
rect 100 10 102 30
rect 110 10 112 30
rect 120 10 122 30
rect 130 10 132 30
<< ptransistor >>
rect 20 42 22 69
rect 30 42 32 69
rect 40 42 42 69
rect 50 42 52 69
rect 70 42 72 69
rect 80 42 82 69
rect 100 42 102 69
rect 110 42 112 69
rect 120 42 122 69
<< polycontact >>
rect 11 34 15 38
rect 18 34 22 38
rect 51 34 55 38
rect 58 34 62 38
rect 119 34 123 38
rect 127 34 131 38
<< ndcontact >>
rect 4 25 8 29
rect 4 18 8 22
rect 14 18 18 22
rect 14 11 18 15
rect 24 25 28 29
rect 24 18 28 22
rect 34 11 38 15
rect 44 18 48 22
rect 54 25 58 29
rect 64 18 68 22
rect 74 25 78 29
rect 84 21 88 25
rect 94 25 98 29
rect 104 25 108 29
rect 114 17 118 21
rect 124 25 128 29
rect 134 25 138 29
rect 134 18 138 22
<< pdcontact >>
rect 14 64 18 68
rect 14 57 18 61
rect 24 50 28 54
rect 24 43 28 47
rect 34 64 38 68
rect 34 57 38 61
rect 44 50 48 54
rect 44 43 48 47
rect 54 64 58 68
rect 64 64 68 68
rect 54 57 58 61
rect 64 57 68 61
rect 74 50 78 54
rect 74 43 78 47
rect 84 64 88 68
rect 84 57 88 61
rect 94 50 98 54
rect 94 43 98 47
rect 104 64 108 68
rect 104 57 108 61
rect 114 50 118 54
rect 114 43 118 47
rect 124 64 128 68
rect 124 57 128 61
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
rect 90 -2 94 2
rect 98 -2 102 2
rect 106 -2 110 2
rect 114 -2 118 2
rect 122 -2 126 2
rect 130 -2 134 2
rect 138 -2 142 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
rect 90 78 94 82
rect 98 78 102 82
rect 106 78 110 82
rect 114 78 118 82
rect 122 78 126 82
rect 130 78 134 82
rect 138 78 142 82
<< psubstratepdiff >>
rect 0 2 144 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 122 2
rect 126 -2 130 2
rect 134 -2 138 2
rect 142 -2 144 2
rect 0 -3 144 -2
<< nsubstratendiff >>
rect 0 82 144 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect 118 78 122 82
rect 126 78 130 82
rect 134 78 138 82
rect 142 78 144 82
rect 0 77 144 78
<< labels >>
rlabel metal1 6 23 6 23 6 n1
rlabel metal1 4 44 4 44 6 a
rlabel polycontact 12 36 12 36 6 a
rlabel polycontact 20 36 20 36 6 a
rlabel metal1 26 24 26 24 6 n1
rlabel metal1 44 32 44 32 6 b
rlabel metal1 28 44 28 44 6 z
rlabel metal1 44 44 44 44 6 z
rlabel metal1 52 44 52 44 6 z
rlabel polycontact 52 36 52 36 6 b
rlabel metal1 36 44 36 44 6 z
rlabel metal1 72 6 72 6 6 vss
rlabel metal1 66 27 66 27 6 n2
rlabel metal1 60 44 60 44 6 z
rlabel polycontact 60 36 60 36 6 b
rlabel metal1 84 44 84 44 6 z
rlabel metal1 68 44 68 44 6 z
rlabel pdcontact 76 52 76 52 6 z
rlabel metal1 72 74 72 74 6 vdd
rlabel metal1 56 20 56 20 6 n1
rlabel metal1 96 25 96 25 6 n2
rlabel metal1 92 44 92 44 6 z
rlabel metal1 100 44 100 44 6 z
rlabel metal1 108 36 108 36 6 z
rlabel metal1 116 28 116 28 6 z
rlabel ndcontact 116 19 116 19 6 n2
rlabel metal1 136 23 136 23 6 n2
rlabel metal1 124 28 124 28 6 z
rlabel metal1 132 40 132 40 6 c
rlabel metal1 124 36 124 36 6 c
rlabel pdcontact 116 52 116 52 6 z
<< end >>
