.subckt oai21v0x1 a1 a2 b vdd vss z
*   SPICE3 file   created from oai21v0x1.ext -      technology: scmos
m00 vdd    vdd    w1     vdd p w=28u  l=2.3636u ad=182.667p pd=56.6667u as=196p     ps=70u
m01 w2     a1     vdd    vdd p w=28u  l=2.3636u ad=196p     pd=70u      as=182.667p ps=56.6667u
m02 z      a2     w2     vdd p w=28u  l=2.3636u ad=176p     pd=50u      as=196p     ps=70u
m03 vdd    b      z      vdd p w=28u  l=2.3636u ad=182.667p pd=56.6667u as=176p     ps=50u
m04 vss    vdd    w3     vss n w=20u  l=2.3636u ad=137.333p pd=46u      as=140p     ps=54u
m05 w4     a1     vss    vss n w=20u  l=2.3636u ad=137.333p pd=46u      as=137.333p ps=46u
m06 w4     a2     vss    vss n w=20u  l=2.3636u ad=137.333p pd=46u      as=137.333p ps=46u
m07 z      b      w4     vss n w=20u  l=2.3636u ad=140p     pd=54u      as=137.333p ps=46u
C0  b      a1     0.040f
C1  z      a2     0.174f
C2  vss    w2     0.004f
C3  a2     a1     0.141f
C4  z      vdd    0.021f
C5  w4     z      0.163f
C6  vss    b      0.010f
C7  a1     vdd    0.075f
C8  w2     b      0.004f
C9  vss    a2     0.023f
C10 w4     a1     0.011f
C11 w2     a2     0.027f
C12 vss    vdd    0.010f
C13 w4     vss    0.240f
C14 w2     vdd    0.093f
C15 b      a2     0.110f
C16 w4     w2     0.025f
C17 z      a1     0.033f
C18 b      vdd    0.067f
C19 a2     vdd    0.031f
C20 w4     a2     0.023f
C21 vss    z      0.033f
C22 vss    a1     0.011f
C23 w2     z      0.010f
C24 w2     a1     0.027f
C25 b      z      0.254f
C26 w4     vss    0.002f
C28 w2     vss    0.004f
C29 b      vss    0.044f
C30 z      vss    0.006f
C31 a2     vss    0.045f
C32 a1     vss    0.045f
.ends
