magic
tech scmos
timestamp 1179385993
<< checkpaint >>
rect -22 -25 46 105
<< ab >>
rect 0 0 24 80
<< pwell >>
rect -4 -7 28 36
<< nwell >>
rect -4 36 28 87
<< polysilicon >>
rect 9 62 11 66
rect 9 41 11 44
rect 9 40 22 41
rect 9 36 17 40
rect 21 36 22 40
rect 9 35 22 36
rect 9 30 11 35
rect 9 18 11 23
<< ndiffusion >>
rect 2 29 9 30
rect 2 25 3 29
rect 7 25 9 29
rect 2 23 9 25
rect 11 23 20 30
rect 13 22 20 23
rect 13 18 14 22
rect 18 18 20 22
rect 13 17 20 18
<< pdiffusion >>
rect 13 72 20 73
rect 13 68 14 72
rect 18 68 20 72
rect 13 62 20 68
rect 4 50 9 62
rect 2 49 9 50
rect 2 45 3 49
rect 7 45 9 49
rect 2 44 9 45
rect 11 44 20 62
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect -2 72 26 78
rect -2 68 14 72
rect 18 68 26 72
rect 2 57 22 63
rect 2 49 7 50
rect 2 45 3 49
rect 2 31 7 45
rect 18 41 22 57
rect 16 40 22 41
rect 16 36 17 40
rect 21 36 22 40
rect 16 35 22 36
rect 2 29 22 31
rect 2 25 3 29
rect 7 25 22 29
rect 13 18 14 22
rect 18 18 19 22
rect 13 12 19 18
rect -2 2 26 12
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
<< ntransistor >>
rect 9 23 11 30
<< ptransistor >>
rect 9 44 11 62
<< polycontact >>
rect 17 36 21 40
<< ndcontact >>
rect 3 25 7 29
rect 14 18 18 22
<< pdcontact >>
rect 14 68 18 72
rect 3 45 7 49
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
<< psubstratepdiff >>
rect 0 2 24 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 24 2
rect 0 -3 24 -2
<< nsubstratendiff >>
rect 0 82 24 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 24 82
rect 0 77 24 78
<< labels >>
rlabel metal1 4 36 4 36 6 z
rlabel metal1 4 60 4 60 6 a
rlabel metal1 12 6 12 6 6 vss
rlabel metal1 12 28 12 28 6 z
rlabel metal1 12 60 12 60 6 a
rlabel metal1 12 74 12 74 6 vdd
rlabel metal1 20 28 20 28 6 z
rlabel metal1 20 52 20 52 6 a
<< end >>
