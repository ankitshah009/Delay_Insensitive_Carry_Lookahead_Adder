magic
tech scmos
timestamp 1179386171
<< checkpaint >>
rect -22 -25 78 105
<< ab >>
rect 0 0 56 80
<< pwell >>
rect -4 -7 60 36
<< nwell >>
rect -4 36 60 87
<< polysilicon >>
rect 9 63 11 68
rect 22 63 24 68
rect 32 63 34 68
rect 44 61 46 65
rect 9 37 11 51
rect 22 47 24 51
rect 16 46 24 47
rect 16 42 17 46
rect 21 42 24 46
rect 16 41 24 42
rect 9 36 15 37
rect 9 32 10 36
rect 14 32 15 36
rect 9 31 15 32
rect 22 31 24 41
rect 32 40 34 51
rect 44 46 46 49
rect 41 45 47 46
rect 41 41 42 45
rect 46 41 47 45
rect 41 40 47 41
rect 32 38 37 40
rect 35 36 37 38
rect 35 35 41 36
rect 35 31 36 35
rect 40 31 41 35
rect 9 26 11 31
rect 22 29 30 31
rect 28 26 30 29
rect 35 30 41 31
rect 35 26 37 30
rect 45 26 47 40
rect 9 15 11 20
rect 28 11 30 16
rect 35 11 37 16
rect 45 15 47 20
<< ndiffusion >>
rect 2 25 9 26
rect 2 21 3 25
rect 7 21 9 25
rect 2 20 9 21
rect 11 20 17 26
rect 23 24 28 26
rect 13 14 17 20
rect 21 23 28 24
rect 21 19 22 23
rect 26 19 28 23
rect 21 18 28 19
rect 23 16 28 18
rect 30 16 35 26
rect 37 25 45 26
rect 37 21 39 25
rect 43 21 45 25
rect 37 20 45 21
rect 47 25 54 26
rect 47 21 49 25
rect 53 21 54 25
rect 47 20 54 21
rect 37 16 43 20
rect 13 12 19 14
rect 13 8 14 12
rect 18 8 19 12
rect 13 7 19 8
<< pdiffusion >>
rect 4 57 9 63
rect 2 56 9 57
rect 2 52 3 56
rect 7 52 9 56
rect 2 51 9 52
rect 11 62 22 63
rect 11 58 15 62
rect 19 58 22 62
rect 11 51 22 58
rect 24 57 32 63
rect 24 53 26 57
rect 30 53 32 57
rect 24 51 32 53
rect 34 62 42 63
rect 34 58 36 62
rect 40 61 42 62
rect 40 58 44 61
rect 34 51 44 58
rect 36 49 44 51
rect 46 55 51 61
rect 46 54 53 55
rect 46 50 48 54
rect 52 50 53 54
rect 46 49 53 50
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect -2 68 58 78
rect 15 62 19 68
rect 15 57 19 58
rect 26 57 30 63
rect 35 62 41 68
rect 35 58 36 62
rect 40 58 41 62
rect 3 56 7 57
rect 3 46 7 52
rect 2 42 17 46
rect 21 42 22 46
rect 2 26 6 42
rect 10 36 22 39
rect 14 33 22 36
rect 2 25 7 26
rect 2 21 3 25
rect 2 20 7 21
rect 10 17 14 32
rect 18 19 22 23
rect 26 19 30 53
rect 34 47 38 55
rect 47 50 48 54
rect 52 50 54 54
rect 34 45 47 47
rect 34 41 42 45
rect 46 41 47 45
rect 50 35 54 50
rect 35 31 36 35
rect 40 31 54 35
rect 50 26 54 31
rect 18 17 30 19
rect 39 25 43 26
rect 39 12 43 21
rect 49 25 54 26
rect 53 21 54 25
rect 49 20 54 21
rect -2 8 14 12
rect 18 8 58 12
rect -2 2 58 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
<< ntransistor >>
rect 9 20 11 26
rect 28 16 30 26
rect 35 16 37 26
rect 45 20 47 26
<< ptransistor >>
rect 9 51 11 63
rect 22 51 24 63
rect 32 51 34 63
rect 44 49 46 61
<< polycontact >>
rect 17 42 21 46
rect 10 32 14 36
rect 42 41 46 45
rect 36 31 40 35
<< ndcontact >>
rect 3 21 7 25
rect 22 19 26 23
rect 39 21 43 25
rect 49 21 53 25
rect 14 8 18 12
<< pdcontact >>
rect 3 52 7 56
rect 15 58 19 62
rect 26 53 30 57
rect 36 58 40 62
rect 48 50 52 54
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
<< psubstratepdiff >>
rect 0 2 56 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 56 2
rect 0 -3 56 -2
<< nsubstratendiff >>
rect 0 82 56 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 56 82
rect 0 77 56 78
<< labels >>
rlabel polycontact 20 44 20 44 6 bn
rlabel polycontact 38 33 38 33 6 an
rlabel metal1 5 49 5 49 6 bn
rlabel metal1 4 33 4 33 6 bn
rlabel metal1 20 20 20 20 6 z
rlabel metal1 12 28 12 28 6 b
rlabel metal1 20 36 20 36 6 b
rlabel metal1 12 44 12 44 6 bn
rlabel metal1 28 6 28 6 6 vss
rlabel metal1 28 40 28 40 6 z
rlabel metal1 36 48 36 48 6 a
rlabel metal1 28 74 28 74 6 vdd
rlabel metal1 44 33 44 33 6 an
rlabel polycontact 44 44 44 44 6 a
rlabel metal1 52 37 52 37 6 an
rlabel pdcontact 50 52 50 52 6 an
<< end >>
