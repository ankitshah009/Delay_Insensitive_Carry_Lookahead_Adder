magic
tech scmos
timestamp 1179385864
<< checkpaint >>
rect -22 -25 46 105
<< ab >>
rect 0 0 24 80
<< pwell >>
rect -4 -7 28 36
<< nwell >>
rect -4 36 28 87
<< polysilicon >>
rect 9 62 15 63
rect 9 58 10 62
rect 14 58 15 62
rect 9 57 15 58
rect 9 54 11 57
rect 9 30 11 42
rect 9 17 11 22
<< ndiffusion >>
rect 2 29 9 30
rect 2 25 3 29
rect 7 25 9 29
rect 2 24 9 25
rect 4 22 9 24
rect 11 27 18 30
rect 11 23 13 27
rect 17 23 18 27
rect 11 22 18 23
<< pdiffusion >>
rect 2 72 8 73
rect 2 68 3 72
rect 7 68 8 72
rect 2 65 8 68
rect 2 54 7 65
rect 2 42 9 54
rect 11 48 16 54
rect 11 47 18 48
rect 11 43 13 47
rect 17 43 18 47
rect 11 42 18 43
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect -2 72 26 78
rect -2 68 3 72
rect 7 68 26 72
rect 2 62 14 63
rect 2 58 10 62
rect 2 57 14 58
rect 2 49 6 57
rect 10 43 13 47
rect 17 43 18 47
rect 10 39 14 43
rect 2 33 14 39
rect 2 29 8 33
rect 2 25 3 29
rect 7 25 8 29
rect 13 27 17 28
rect 13 12 17 23
rect -2 2 26 12
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
<< ntransistor >>
rect 9 22 11 30
<< ptransistor >>
rect 9 42 11 54
<< polycontact >>
rect 10 58 14 62
<< ndcontact >>
rect 3 25 7 29
rect 13 23 17 27
<< pdcontact >>
rect 3 68 7 72
rect 13 43 17 47
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
<< psubstratepdiff >>
rect 0 2 24 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 24 2
rect 0 -3 24 -2
<< nsubstratendiff >>
rect 0 82 24 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 24 82
rect 0 77 24 78
<< labels >>
rlabel metal1 4 32 4 32 6 z
rlabel metal1 4 56 4 56 6 a
rlabel metal1 12 6 12 6 6 vss
rlabel metal1 12 40 12 40 6 z
rlabel polycontact 12 60 12 60 6 a
rlabel metal1 12 74 12 74 6 vdd
<< end >>
