magic
tech scmos
timestamp 1185039028
<< checkpaint >>
rect -22 -24 62 124
<< ab >>
rect 0 0 40 100
<< pwell >>
rect -2 -4 42 49
<< nwell >>
rect -2 49 42 104
<< polysilicon >>
rect 19 95 21 98
rect 27 95 29 98
rect 19 53 21 55
rect 17 52 23 53
rect 17 49 18 52
rect 13 48 18 49
rect 22 48 23 52
rect 13 47 23 48
rect 13 25 15 47
rect 27 43 29 55
rect 27 42 33 43
rect 27 41 28 42
rect 25 38 28 41
rect 32 38 33 42
rect 25 37 33 38
rect 25 25 27 37
rect 13 12 15 15
rect 25 12 27 15
<< ndiffusion >>
rect 5 15 13 25
rect 15 22 25 25
rect 15 18 18 22
rect 22 18 25 22
rect 15 15 25 18
rect 27 15 35 25
rect 5 12 11 15
rect 29 12 35 15
rect 5 8 6 12
rect 10 8 11 12
rect 5 7 11 8
rect 29 8 30 12
rect 34 8 35 12
rect 29 7 35 8
<< pdiffusion >>
rect 15 85 19 95
rect 7 82 19 85
rect 7 78 8 82
rect 12 78 19 82
rect 7 72 19 78
rect 7 68 8 72
rect 12 68 19 72
rect 7 62 19 68
rect 7 58 8 62
rect 12 58 19 62
rect 7 55 19 58
rect 21 55 27 95
rect 29 92 37 95
rect 29 88 32 92
rect 36 88 37 92
rect 29 55 37 88
<< metal1 >>
rect -2 92 42 101
rect -2 88 32 92
rect 36 88 42 92
rect -2 87 42 88
rect 7 82 13 83
rect 7 78 8 82
rect 12 78 13 82
rect 7 72 13 78
rect 7 68 8 72
rect 12 68 13 72
rect 7 62 13 68
rect 7 58 8 62
rect 12 58 13 62
rect 7 23 13 58
rect 17 52 23 82
rect 17 48 18 52
rect 22 48 23 52
rect 17 28 23 48
rect 27 42 33 82
rect 27 38 28 42
rect 32 38 33 42
rect 7 22 23 23
rect 7 18 18 22
rect 22 18 23 22
rect 27 18 33 38
rect 8 17 23 18
rect -2 12 42 13
rect -2 8 6 12
rect 10 8 30 12
rect 34 8 42 12
rect -2 -1 42 8
<< ntransistor >>
rect 13 15 15 25
rect 25 15 27 25
<< ptransistor >>
rect 19 55 21 95
rect 27 55 29 95
<< polycontact >>
rect 18 48 22 52
rect 28 38 32 42
<< ndcontact >>
rect 18 18 22 22
rect 6 8 10 12
rect 30 8 34 12
<< pdcontact >>
rect 8 78 12 82
rect 8 68 12 72
rect 8 58 12 62
rect 32 88 36 92
<< labels >>
rlabel metal1 10 50 10 50 6 nq
rlabel metal1 10 50 10 50 6 nq
rlabel metal1 20 6 20 6 6 vss
rlabel metal1 20 6 20 6 6 vss
rlabel metal1 30 50 30 50 6 i0
rlabel metal1 30 50 30 50 6 i0
rlabel metal1 20 55 20 55 6 i1
rlabel metal1 20 55 20 55 6 i1
rlabel metal1 20 94 20 94 6 vdd
rlabel metal1 20 94 20 94 6 vdd
<< end >>
