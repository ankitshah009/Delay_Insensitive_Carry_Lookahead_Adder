magic
tech scmos
timestamp 1179386817
<< checkpaint >>
rect -22 -25 86 105
<< ab >>
rect 0 0 64 80
<< pwell >>
rect -4 -7 68 36
<< nwell >>
rect -4 36 68 87
<< polysilicon >>
rect 12 70 14 74
rect 19 70 21 74
rect 29 70 31 74
rect 36 70 38 74
rect 46 70 48 74
rect 53 70 55 74
rect 12 39 14 42
rect 19 39 21 42
rect 29 39 31 42
rect 9 38 15 39
rect 9 34 10 38
rect 14 34 15 38
rect 19 38 31 39
rect 19 37 23 38
rect 9 33 15 34
rect 22 34 23 37
rect 27 37 31 38
rect 36 39 38 42
rect 46 39 48 42
rect 53 39 55 42
rect 36 38 48 39
rect 27 34 28 37
rect 22 33 28 34
rect 36 34 37 38
rect 41 37 48 38
rect 52 38 58 39
rect 41 34 44 37
rect 36 33 44 34
rect 13 30 15 33
rect 23 30 25 33
rect 42 30 44 33
rect 52 34 53 38
rect 57 34 58 38
rect 52 33 58 34
rect 52 30 54 33
rect 13 6 15 10
rect 23 6 25 10
rect 42 6 44 10
rect 52 6 54 10
<< ndiffusion >>
rect 5 15 13 30
rect 5 11 7 15
rect 11 11 13 15
rect 5 10 13 11
rect 15 22 23 30
rect 15 18 17 22
rect 21 18 23 22
rect 15 10 23 18
rect 25 15 42 30
rect 25 11 32 15
rect 36 11 42 15
rect 25 10 42 11
rect 44 29 52 30
rect 44 25 46 29
rect 50 25 52 29
rect 44 22 52 25
rect 44 18 46 22
rect 50 18 52 22
rect 44 10 52 18
rect 54 22 62 30
rect 54 18 57 22
rect 61 18 62 22
rect 54 15 62 18
rect 54 11 57 15
rect 61 11 62 15
rect 54 10 62 11
<< pdiffusion >>
rect 7 55 12 70
rect 5 54 12 55
rect 5 50 6 54
rect 10 50 12 54
rect 5 47 12 50
rect 5 43 6 47
rect 10 43 12 47
rect 5 42 12 43
rect 14 42 19 70
rect 21 69 29 70
rect 21 65 23 69
rect 27 65 29 69
rect 21 62 29 65
rect 21 58 23 62
rect 27 58 29 62
rect 21 42 29 58
rect 31 42 36 70
rect 38 62 46 70
rect 38 58 40 62
rect 44 58 46 62
rect 38 55 46 58
rect 38 51 40 55
rect 44 51 46 55
rect 38 42 46 51
rect 48 42 53 70
rect 55 69 62 70
rect 55 65 57 69
rect 61 65 62 69
rect 55 62 62 65
rect 55 58 57 62
rect 61 58 62 62
rect 55 42 62 58
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect -2 69 66 78
rect -2 68 23 69
rect 22 65 23 68
rect 27 68 57 69
rect 27 65 28 68
rect 22 62 28 65
rect 56 65 57 68
rect 61 68 66 69
rect 61 65 62 68
rect 22 58 23 62
rect 27 58 28 62
rect 40 62 46 63
rect 44 58 46 62
rect 56 62 62 65
rect 56 58 57 62
rect 61 58 62 62
rect 40 55 46 58
rect 5 50 6 54
rect 10 51 40 54
rect 44 51 46 55
rect 10 50 46 51
rect 5 47 11 50
rect 2 22 6 47
rect 10 43 11 47
rect 22 42 55 46
rect 10 38 18 39
rect 14 34 18 38
rect 22 38 28 42
rect 49 38 55 42
rect 22 34 23 38
rect 27 34 28 38
rect 33 34 37 38
rect 41 34 42 38
rect 49 34 53 38
rect 57 34 58 38
rect 10 33 18 34
rect 14 30 18 33
rect 33 30 39 34
rect 14 26 39 30
rect 46 29 51 30
rect 50 25 51 29
rect 46 22 51 25
rect 2 18 17 22
rect 21 18 46 22
rect 50 18 51 22
rect 57 22 61 23
rect 57 15 61 18
rect 6 12 7 15
rect -2 11 7 12
rect 11 12 12 15
rect 31 12 32 15
rect 11 11 32 12
rect 36 12 37 15
rect 36 11 57 12
rect 61 11 66 12
rect -2 2 66 11
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
<< ntransistor >>
rect 13 10 15 30
rect 23 10 25 30
rect 42 10 44 30
rect 52 10 54 30
<< ptransistor >>
rect 12 42 14 70
rect 19 42 21 70
rect 29 42 31 70
rect 36 42 38 70
rect 46 42 48 70
rect 53 42 55 70
<< polycontact >>
rect 10 34 14 38
rect 23 34 27 38
rect 37 34 41 38
rect 53 34 57 38
<< ndcontact >>
rect 7 11 11 15
rect 17 18 21 22
rect 32 11 36 15
rect 46 25 50 29
rect 46 18 50 22
rect 57 18 61 22
rect 57 11 61 15
<< pdcontact >>
rect 6 50 10 54
rect 6 43 10 47
rect 23 65 27 69
rect 23 58 27 62
rect 40 58 44 62
rect 40 51 44 55
rect 57 65 61 69
rect 57 58 61 62
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
<< psubstratepdiff >>
rect 0 2 64 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 64 2
rect 0 -3 64 -2
<< nsubstratendiff >>
rect 0 82 64 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 64 82
rect 0 77 64 78
<< labels >>
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 20 12 20 6 z
rlabel metal1 20 28 20 28 6 b
rlabel ndcontact 20 20 20 20 6 z
rlabel polycontact 12 36 12 36 6 b
rlabel metal1 20 52 20 52 6 z
rlabel metal1 12 52 12 52 6 z
rlabel metal1 32 6 32 6 6 vss
rlabel metal1 28 28 28 28 6 b
rlabel metal1 28 20 28 20 6 z
rlabel metal1 36 20 36 20 6 z
rlabel metal1 36 32 36 32 6 b
rlabel metal1 28 44 28 44 6 a
rlabel metal1 36 44 36 44 6 a
rlabel metal1 36 52 36 52 6 z
rlabel metal1 28 52 28 52 6 z
rlabel metal1 32 74 32 74 6 vdd
rlabel metal1 44 20 44 20 6 z
rlabel metal1 44 44 44 44 6 a
rlabel metal1 44 60 44 60 6 z
rlabel metal1 52 40 52 40 6 a
<< end >>
