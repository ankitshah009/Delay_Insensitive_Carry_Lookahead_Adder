magic
tech scmos
timestamp 1179387568
<< checkpaint >>
rect -22 -22 94 94
<< ab >>
rect 0 0 72 72
<< pwell >>
rect -4 -4 76 32
<< nwell >>
rect -4 32 76 76
<< polysilicon >>
rect 32 62 34 67
rect 42 62 44 67
rect 49 62 51 67
rect 13 58 15 62
rect 21 58 23 62
rect 13 36 15 42
rect 21 39 23 42
rect 9 35 15 36
rect 9 31 10 35
rect 14 31 15 35
rect 9 30 15 31
rect 19 38 25 39
rect 61 57 63 61
rect 61 38 63 41
rect 19 34 20 38
rect 24 34 25 38
rect 19 33 25 34
rect 32 33 34 38
rect 42 35 44 38
rect 9 26 11 30
rect 19 26 21 33
rect 29 31 34 33
rect 39 34 45 35
rect 29 26 31 31
rect 39 30 40 34
rect 44 30 45 34
rect 39 29 45 30
rect 43 24 45 29
rect 49 30 51 38
rect 61 37 70 38
rect 61 36 65 37
rect 64 33 65 36
rect 69 33 70 37
rect 64 32 70 33
rect 49 28 57 30
rect 55 27 57 28
rect 55 26 63 27
rect 43 21 47 24
rect 19 14 21 19
rect 9 7 11 12
rect 29 4 31 19
rect 45 18 47 21
rect 55 22 58 26
rect 62 22 63 26
rect 55 21 63 22
rect 55 18 57 21
rect 45 8 47 12
rect 55 8 57 12
rect 68 4 70 32
rect 29 2 70 4
<< ndiffusion >>
rect 4 18 9 26
rect 2 17 9 18
rect 2 13 3 17
rect 7 13 9 17
rect 2 12 9 13
rect 11 24 19 26
rect 11 20 13 24
rect 17 20 19 24
rect 11 19 19 20
rect 21 25 29 26
rect 21 21 23 25
rect 27 21 29 25
rect 21 19 29 21
rect 31 19 41 26
rect 11 12 16 19
rect 33 18 41 19
rect 33 12 45 18
rect 47 17 55 18
rect 47 13 49 17
rect 53 13 55 17
rect 47 12 55 13
rect 57 17 64 18
rect 57 13 59 17
rect 63 13 64 17
rect 57 12 64 13
rect 33 11 43 12
rect 33 7 38 11
rect 42 7 43 11
rect 33 6 43 7
<< pdiffusion >>
rect 4 68 11 69
rect 4 64 6 68
rect 10 64 11 68
rect 53 68 59 69
rect 4 58 11 64
rect 53 64 54 68
rect 58 64 59 68
rect 53 62 59 64
rect 25 58 32 62
rect 4 42 13 58
rect 15 42 21 58
rect 23 57 32 58
rect 23 53 25 57
rect 29 53 32 57
rect 23 42 32 53
rect 27 38 32 42
rect 34 43 42 62
rect 34 39 36 43
rect 40 39 42 43
rect 34 38 42 39
rect 44 38 49 62
rect 51 57 59 62
rect 51 41 61 57
rect 63 56 70 57
rect 63 52 65 56
rect 69 52 70 56
rect 63 51 70 52
rect 63 41 68 51
rect 51 38 59 41
<< metal1 >>
rect -2 68 74 72
rect -2 64 6 68
rect 10 64 54 68
rect 58 64 64 68
rect 68 64 74 68
rect 2 57 31 58
rect 2 54 25 57
rect 2 24 6 54
rect 24 53 25 54
rect 29 54 31 57
rect 36 56 69 59
rect 36 55 65 56
rect 29 53 30 54
rect 36 50 40 55
rect 65 51 69 52
rect 10 46 40 50
rect 10 35 14 46
rect 31 39 36 43
rect 40 39 41 43
rect 31 38 35 39
rect 19 34 20 38
rect 24 34 35 38
rect 50 35 54 51
rect 58 43 62 51
rect 58 39 70 43
rect 65 37 70 39
rect 10 27 27 31
rect 23 25 27 27
rect 2 20 13 24
rect 17 20 18 24
rect 23 20 27 21
rect 31 20 35 34
rect 40 34 54 35
rect 44 30 54 34
rect 40 29 54 30
rect 58 27 62 35
rect 69 33 70 37
rect 65 32 70 33
rect 66 31 70 32
rect 58 26 70 27
rect 62 22 70 26
rect 58 21 70 22
rect 31 17 54 20
rect 2 13 3 17
rect 7 16 49 17
rect 7 13 35 16
rect 48 13 49 16
rect 53 13 54 17
rect 58 13 59 17
rect 63 13 64 17
rect 38 11 42 12
rect -2 4 21 8
rect 25 7 38 8
rect 58 8 64 13
rect 42 7 74 8
rect 25 4 74 7
rect -2 0 74 4
<< ntransistor >>
rect 9 12 11 26
rect 19 19 21 26
rect 29 19 31 26
rect 45 12 47 18
rect 55 12 57 18
<< ptransistor >>
rect 13 42 15 58
rect 21 42 23 58
rect 32 38 34 62
rect 42 38 44 62
rect 49 38 51 62
rect 61 41 63 57
<< polycontact >>
rect 10 31 14 35
rect 20 34 24 38
rect 40 30 44 34
rect 65 33 69 37
rect 58 22 62 26
<< ndcontact >>
rect 3 13 7 17
rect 13 20 17 24
rect 23 21 27 25
rect 49 13 53 17
rect 59 13 63 17
rect 38 7 42 11
<< pdcontact >>
rect 6 64 10 68
rect 54 64 58 68
rect 25 53 29 57
rect 36 39 40 43
rect 65 52 69 56
<< psubstratepcontact >>
rect 21 4 25 8
<< nsubstratencontact >>
rect 64 64 68 68
<< psubstratepdiff >>
rect 20 8 26 9
rect 20 4 21 8
rect 25 4 26 8
rect 20 3 26 4
<< nsubstratendiff >>
rect 63 68 69 69
rect 63 64 64 68
rect 68 64 69 68
rect 63 63 69 64
<< labels >>
rlabel ptransistor 22 47 22 47 6 an
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 38 12 38 6 bn
rlabel metal1 12 56 12 56 6 z
rlabel metal1 18 15 18 15 6 an
rlabel metal1 25 25 25 25 6 bn
rlabel metal1 27 36 27 36 6 an
rlabel pdcontact 28 56 28 56 6 z
rlabel metal1 20 56 20 56 6 z
rlabel metal1 36 4 36 4 6 vss
rlabel metal1 42 18 42 18 6 an
rlabel metal1 44 32 44 32 6 a2
rlabel metal1 52 40 52 40 6 a2
rlabel metal1 36 41 36 41 6 an
rlabel metal1 36 68 36 68 6 vdd
rlabel metal1 60 28 60 28 6 a1
rlabel metal1 68 24 68 24 6 a1
rlabel metal1 68 40 68 40 6 b
rlabel metal1 60 48 60 48 6 b
rlabel metal1 52 57 52 57 6 bn
<< end >>
