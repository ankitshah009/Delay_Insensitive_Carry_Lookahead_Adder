.subckt iv1v0x2 a vdd vss z
*   SPICE3 file   created from iv1v0x2.ext -      technology: scmos
m00 vdd    vdd    w1     vdd p w=28u  l=2.3636u ad=176p     pd=50u      as=196p     ps=70u
m01 z      a      vdd    vdd p w=28u  l=2.3636u ad=196p     pd=70u      as=176p     ps=50u
m02 vss    vdd    w2     vss n w=20u  l=2.3636u ad=136p     pd=42u      as=140p     ps=54u
m03 z      a      vss    vss n w=20u  l=2.3636u ad=140p     pd=54u      as=136p     ps=42u
C0  a      vdd    0.075f
C1  vss    z      0.104f
C2  vss    a      0.011f
C3  z      a      0.279f
C4  vss    vdd    0.007f
C5  z      vdd    0.126f
C7  z      vss    0.006f
C8  a      vss    0.045f
.ends
