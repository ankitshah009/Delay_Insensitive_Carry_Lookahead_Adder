magic
tech scmos
timestamp 1179385822
<< checkpaint >>
rect -22 -25 46 105
<< ab >>
rect 0 0 24 80
<< pwell >>
rect -4 -7 28 36
<< nwell >>
rect -4 36 28 87
<< polysilicon >>
rect 9 70 11 74
rect 9 39 11 42
rect 9 38 16 39
rect 9 34 11 38
rect 15 34 16 38
rect 9 33 16 34
rect 9 30 11 33
rect 9 11 11 16
<< ndiffusion >>
rect 2 29 9 30
rect 2 25 3 29
rect 7 25 9 29
rect 2 22 9 25
rect 2 18 3 22
rect 7 18 9 22
rect 2 16 9 18
rect 11 28 19 30
rect 11 24 13 28
rect 17 24 19 28
rect 11 21 19 24
rect 11 17 13 21
rect 17 17 19 21
rect 11 16 19 17
<< pdiffusion >>
rect 4 56 9 70
rect 2 55 9 56
rect 2 51 3 55
rect 7 51 9 55
rect 2 48 9 51
rect 2 44 3 48
rect 7 44 9 48
rect 2 42 9 44
rect 11 69 19 70
rect 11 65 13 69
rect 17 65 19 69
rect 11 62 19 65
rect 11 58 13 62
rect 17 58 19 62
rect 11 42 19 58
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect -2 69 26 78
rect -2 68 13 69
rect 12 65 13 68
rect 17 68 26 69
rect 17 65 18 68
rect 12 62 18 65
rect 12 58 13 62
rect 17 58 18 62
rect 2 51 3 55
rect 7 51 14 55
rect 2 49 14 51
rect 2 48 7 49
rect 2 44 3 48
rect 2 43 7 44
rect 2 30 6 43
rect 18 39 22 55
rect 10 38 22 39
rect 10 34 11 38
rect 15 34 22 38
rect 10 33 22 34
rect 2 29 7 30
rect 2 25 3 29
rect 2 22 7 25
rect 2 18 3 22
rect 2 17 7 18
rect 13 28 17 29
rect 13 21 17 24
rect 13 12 17 17
rect -2 2 26 12
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
<< ntransistor >>
rect 9 16 11 30
<< ptransistor >>
rect 9 42 11 70
<< polycontact >>
rect 11 34 15 38
<< ndcontact >>
rect 3 25 7 29
rect 3 18 7 22
rect 13 24 17 28
rect 13 17 17 21
<< pdcontact >>
rect 3 51 7 55
rect 3 44 7 48
rect 13 65 17 69
rect 13 58 17 62
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
<< psubstratepdiff >>
rect 0 2 24 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 24 2
rect 0 -3 24 -2
<< nsubstratendiff >>
rect 0 82 24 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 24 82
rect 0 77 24 78
<< labels >>
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 6 12 6 6 vss
rlabel polycontact 12 36 12 36 6 a
rlabel metal1 12 52 12 52 6 z
rlabel metal1 12 74 12 74 6 vdd
rlabel metal1 20 44 20 44 6 a
<< end >>
