.subckt xor2v2x05 a b vdd vss z
*   SPICE3 file   created from xor2v2x05.ext -      technology: scmos
m00 z      bn     an     vdd p w=16u  l=2.3636u ad=64p      pd=24u      as=92p      ps=46u
m01 bn     an     z      vdd p w=16u  l=2.3636u ad=64p      pd=24u      as=64p      ps=24u
m02 vdd    b      bn     vdd p w=16u  l=2.3636u ad=110p     pd=36u      as=64p      ps=24u
m03 an     a      vdd    vdd p w=16u  l=2.3636u ad=92p      pd=46u      as=110p     ps=36u
m04 w1     bn     z      vss n w=11u  l=2.3636u ad=27.5p    pd=16u      as=53.3704p ps=27.7037u
m05 vss    an     w1     vss n w=11u  l=2.3636u ad=99.4783p pd=44u      as=27.5p    ps=16u
m06 bn     b      vss    vss n w=6u   l=2.3636u ad=24.8571p pd=13.7143u as=54.2609p ps=24u
m07 z      a      bn     vss n w=8u   l=2.3636u ad=38.8148p pd=20.1481u as=33.1429p ps=18.2857u
m08 an     b      z      vss n w=8u   l=2.3636u ad=33.1429p pd=18.2857u as=38.8148p ps=20.1481u
m09 vss    a      an     vss n w=6u   l=2.3636u ad=54.2609p pd=24u      as=24.8571p ps=13.7143u
C0  vss    vdd    0.003f
C1  a      z      0.003f
C2  z      vdd    0.042f
C3  vss    bn     0.093f
C4  a      an     0.083f
C5  z      bn     0.497f
C6  a      b      0.186f
C7  vdd    an     0.274f
C8  vdd    b      0.080f
C9  an     bn     0.524f
C10 bn     b      0.041f
C11 vss    z      0.274f
C12 a      vdd    0.017f
C13 vss    an     0.089f
C14 w1     bn     0.005f
C15 vss    b      0.029f
C16 a      bn     0.015f
C17 z      an     0.327f
C18 vdd    bn     0.047f
C19 z      b      0.009f
C20 an     b      0.123f
C21 vss    a      0.029f
C22 w1     z      0.010f
C24 a      vss    0.040f
C25 z      vss    0.021f
C27 an     vss    0.039f
C28 bn     vss    0.029f
C29 b      vss    0.061f
.ends
