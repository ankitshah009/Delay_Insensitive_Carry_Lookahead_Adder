magic
tech scmos
timestamp 1179386014
<< checkpaint >>
rect -22 -25 54 105
<< ab >>
rect 0 0 32 80
<< pwell >>
rect -4 -7 36 36
<< nwell >>
rect -4 36 36 87
<< polysilicon >>
rect 9 70 11 74
rect 19 70 21 74
rect 9 39 11 42
rect 19 39 21 42
rect 9 38 22 39
rect 9 34 17 38
rect 21 34 22 38
rect 9 33 22 34
rect 10 30 12 33
rect 20 30 22 33
rect 10 15 12 19
rect 20 15 22 19
<< ndiffusion >>
rect 2 22 10 30
rect 2 18 3 22
rect 7 19 10 22
rect 12 29 20 30
rect 12 25 14 29
rect 18 25 20 29
rect 12 19 20 25
rect 22 25 29 30
rect 22 21 24 25
rect 28 21 29 25
rect 22 19 29 21
rect 7 18 8 19
rect 2 17 8 18
<< pdiffusion >>
rect 2 69 9 70
rect 2 65 3 69
rect 7 65 9 69
rect 2 62 9 65
rect 2 58 3 62
rect 7 58 9 62
rect 2 42 9 58
rect 11 62 19 70
rect 11 58 13 62
rect 17 58 19 62
rect 11 55 19 58
rect 11 51 13 55
rect 17 51 19 55
rect 11 42 19 51
rect 21 69 28 70
rect 21 65 23 69
rect 27 65 28 69
rect 21 62 28 65
rect 21 58 23 62
rect 27 58 28 62
rect 21 42 28 58
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect -2 69 34 78
rect -2 68 3 69
rect 2 65 3 68
rect 7 68 23 69
rect 7 65 8 68
rect 2 62 8 65
rect 22 65 23 68
rect 27 68 34 69
rect 27 65 28 68
rect 2 58 3 62
rect 7 58 8 62
rect 13 62 17 63
rect 22 62 28 65
rect 22 58 23 62
rect 27 58 28 62
rect 13 55 17 58
rect 2 51 13 54
rect 17 51 23 54
rect 2 50 23 51
rect 2 29 6 50
rect 17 39 23 46
rect 17 38 30 39
rect 21 34 30 38
rect 17 33 30 34
rect 2 25 14 29
rect 18 25 19 29
rect 24 25 28 26
rect 2 18 3 22
rect 7 18 8 22
rect 2 12 8 18
rect 24 12 28 21
rect -2 2 34 12
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
<< ntransistor >>
rect 10 19 12 30
rect 20 19 22 30
<< ptransistor >>
rect 9 42 11 70
rect 19 42 21 70
<< polycontact >>
rect 17 34 21 38
<< ndcontact >>
rect 3 18 7 22
rect 14 25 18 29
rect 24 21 28 25
<< pdcontact >>
rect 3 65 7 69
rect 3 58 7 62
rect 13 58 17 62
rect 13 51 17 55
rect 23 65 27 69
rect 23 58 27 62
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
<< psubstratepdiff >>
rect 0 2 32 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 32 2
rect 0 -3 32 -2
<< nsubstratendiff >>
rect 0 82 32 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 32 82
rect 0 77 32 78
<< labels >>
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 52 12 52 6 z
rlabel metal1 16 6 16 6 6 vss
rlabel metal1 20 40 20 40 6 a
rlabel metal1 20 52 20 52 6 z
rlabel metal1 16 74 16 74 6 vdd
rlabel metal1 28 36 28 36 6 a
<< end >>
