magic
tech scmos
timestamp 1180600650
<< checkpaint >>
rect -22 -22 182 122
<< ab >>
rect 0 0 160 100
<< pwell >>
rect -4 -4 164 48
<< nwell >>
rect -4 48 164 104
<< polysilicon >>
rect 13 94 15 98
rect 25 83 27 87
rect 37 84 39 88
rect 73 78 75 82
rect 85 78 87 82
rect 61 72 63 76
rect 13 41 15 55
rect 25 53 27 65
rect 37 63 39 66
rect 37 62 43 63
rect 37 58 38 62
rect 42 58 43 62
rect 37 57 43 58
rect 97 77 99 81
rect 109 77 111 81
rect 145 94 147 98
rect 121 78 123 82
rect 19 52 27 53
rect 19 48 20 52
rect 24 48 27 52
rect 61 53 63 56
rect 73 53 75 56
rect 61 52 75 53
rect 61 51 68 52
rect 19 47 27 48
rect 67 48 68 51
rect 72 51 75 52
rect 85 53 87 56
rect 85 52 93 53
rect 85 51 88 52
rect 72 48 73 51
rect 67 47 73 48
rect 87 48 88 51
rect 92 48 93 52
rect 87 47 93 48
rect 27 42 33 43
rect 27 41 28 42
rect 13 39 28 41
rect 13 25 15 39
rect 27 38 28 39
rect 32 38 33 42
rect 27 37 33 38
rect 37 42 43 43
rect 37 38 38 42
rect 42 38 43 42
rect 37 37 43 38
rect 53 42 59 43
rect 53 38 54 42
rect 58 41 59 42
rect 97 41 99 55
rect 109 43 111 55
rect 121 53 123 56
rect 117 52 123 53
rect 117 48 118 52
rect 122 48 123 52
rect 117 47 123 48
rect 145 43 147 55
rect 58 39 99 41
rect 58 38 59 39
rect 53 37 59 38
rect 19 32 27 33
rect 19 28 20 32
rect 24 28 27 32
rect 37 29 39 37
rect 87 34 93 35
rect 67 32 73 33
rect 67 29 68 32
rect 19 27 27 28
rect 25 24 27 27
rect 61 28 68 29
rect 72 29 73 32
rect 87 31 88 34
rect 85 30 88 31
rect 92 30 93 34
rect 85 29 93 30
rect 72 28 75 29
rect 61 27 75 28
rect 61 24 63 27
rect 73 24 75 27
rect 85 26 87 29
rect 97 27 99 39
rect 107 42 113 43
rect 107 38 108 42
rect 112 41 113 42
rect 127 42 133 43
rect 127 41 128 42
rect 112 39 128 41
rect 112 38 113 39
rect 107 37 113 38
rect 127 38 128 39
rect 132 38 133 42
rect 127 37 133 38
rect 137 42 147 43
rect 137 38 138 42
rect 142 38 147 42
rect 137 37 147 38
rect 117 32 123 33
rect 117 29 118 32
rect 109 28 118 29
rect 122 28 123 32
rect 109 27 123 28
rect 25 11 27 15
rect 37 11 39 15
rect 61 12 63 16
rect 109 24 111 27
rect 121 24 123 27
rect 145 25 147 37
rect 13 2 15 6
rect 73 11 75 15
rect 85 11 87 15
rect 97 11 99 15
rect 109 11 111 15
rect 121 12 123 16
rect 145 2 147 6
<< ndiffusion >>
rect 5 22 13 25
rect 5 18 6 22
rect 10 18 13 22
rect 5 6 13 18
rect 15 24 20 25
rect 29 24 37 29
rect 15 15 25 24
rect 27 15 37 24
rect 39 22 47 29
rect 92 26 97 27
rect 77 24 85 26
rect 39 18 42 22
rect 46 18 47 22
rect 39 15 47 18
rect 53 22 61 24
rect 53 18 54 22
rect 58 18 61 22
rect 53 17 61 18
rect 56 16 61 17
rect 63 16 73 24
rect 15 12 23 15
rect 15 8 18 12
rect 22 8 23 12
rect 65 15 73 16
rect 75 15 85 24
rect 87 24 97 26
rect 87 20 90 24
rect 94 20 97 24
rect 87 15 97 20
rect 99 24 107 27
rect 125 32 133 33
rect 125 28 128 32
rect 132 28 133 32
rect 125 27 133 28
rect 125 24 131 27
rect 99 15 109 24
rect 111 16 121 24
rect 123 16 131 24
rect 140 21 145 25
rect 111 15 119 16
rect 65 12 71 15
rect 15 6 23 8
rect 65 8 66 12
rect 70 8 71 12
rect 113 12 119 15
rect 137 12 145 21
rect 65 7 71 8
rect 113 8 114 12
rect 118 8 119 12
rect 113 7 119 8
rect 137 8 138 12
rect 142 8 145 12
rect 137 6 145 8
rect 147 22 155 25
rect 147 18 150 22
rect 154 18 155 22
rect 147 6 155 18
<< pdiffusion >>
rect 5 82 13 94
rect 5 78 6 82
rect 10 78 13 82
rect 5 72 13 78
rect 5 68 6 72
rect 10 68 13 72
rect 5 62 13 68
rect 5 58 6 62
rect 10 58 13 62
rect 5 55 13 58
rect 15 92 23 94
rect 15 88 18 92
rect 22 88 23 92
rect 41 92 47 93
rect 41 88 42 92
rect 46 88 47 92
rect 15 83 23 88
rect 41 84 47 88
rect 65 92 71 93
rect 65 88 66 92
rect 70 88 71 92
rect 113 92 119 93
rect 29 83 37 84
rect 15 65 25 83
rect 27 72 37 83
rect 27 68 30 72
rect 34 68 37 72
rect 27 66 37 68
rect 39 66 47 84
rect 65 78 71 88
rect 113 88 114 92
rect 118 88 119 92
rect 65 72 73 78
rect 27 65 32 66
rect 15 55 23 65
rect 53 62 61 72
rect 53 58 54 62
rect 58 58 61 62
rect 53 56 61 58
rect 63 56 73 72
rect 75 72 85 78
rect 75 68 78 72
rect 82 68 85 72
rect 75 56 85 68
rect 87 77 95 78
rect 113 78 119 88
rect 137 92 145 94
rect 137 88 138 92
rect 142 88 145 92
rect 137 82 145 88
rect 137 78 138 82
rect 142 78 145 82
rect 113 77 121 78
rect 87 62 97 77
rect 87 58 90 62
rect 94 58 97 62
rect 87 56 97 58
rect 92 55 97 56
rect 99 72 109 77
rect 99 68 102 72
rect 106 68 109 72
rect 99 62 109 68
rect 99 58 102 62
rect 106 58 109 62
rect 99 55 109 58
rect 111 56 121 77
rect 123 61 131 78
rect 137 72 145 78
rect 137 68 138 72
rect 142 68 145 72
rect 137 67 145 68
rect 123 60 133 61
rect 123 56 128 60
rect 132 56 133 60
rect 111 55 116 56
rect 127 55 133 56
rect 140 55 145 67
rect 147 82 155 94
rect 147 78 150 82
rect 154 78 155 82
rect 147 72 155 78
rect 147 68 150 72
rect 154 68 155 72
rect 147 62 155 68
rect 147 58 150 62
rect 154 58 155 62
rect 147 55 155 58
<< metal1 >>
rect -2 96 162 100
rect -2 92 54 96
rect 58 92 78 96
rect 82 92 90 96
rect 94 92 102 96
rect 106 92 126 96
rect 130 92 162 96
rect -2 88 18 92
rect 22 88 42 92
rect 46 88 66 92
rect 70 88 114 92
rect 118 88 138 92
rect 142 88 162 92
rect 8 82 12 83
rect 5 78 6 82
rect 10 78 12 82
rect 8 72 12 78
rect 5 68 6 72
rect 10 68 12 72
rect 8 62 12 68
rect 5 58 6 62
rect 10 58 12 62
rect 8 22 12 58
rect 5 18 6 22
rect 10 18 12 22
rect 8 17 12 18
rect 18 82 22 83
rect 138 82 142 88
rect 18 78 122 82
rect 18 52 22 78
rect 68 72 72 73
rect 102 72 106 73
rect 29 68 30 72
rect 34 68 35 72
rect 40 68 72 72
rect 77 68 78 72
rect 82 68 102 72
rect 18 48 20 52
rect 24 48 25 52
rect 18 32 22 48
rect 29 42 33 68
rect 40 63 44 68
rect 27 38 28 42
rect 32 38 33 42
rect 18 28 20 32
rect 24 28 25 32
rect 18 17 22 28
rect 29 22 33 38
rect 38 62 44 63
rect 42 58 44 62
rect 54 62 58 63
rect 38 42 42 58
rect 38 37 42 38
rect 54 42 58 58
rect 54 22 58 38
rect 29 18 42 22
rect 46 18 47 22
rect 54 17 58 18
rect 68 52 72 68
rect 102 62 106 68
rect 68 32 72 48
rect 68 17 72 28
rect 78 58 90 62
rect 94 58 95 62
rect 78 22 82 58
rect 102 57 106 58
rect 118 52 122 78
rect 138 72 142 78
rect 138 67 142 68
rect 148 82 152 83
rect 148 78 150 82
rect 154 78 155 82
rect 148 72 152 78
rect 148 68 150 72
rect 154 68 155 72
rect 148 62 152 68
rect 87 48 88 52
rect 92 48 118 52
rect 98 38 108 42
rect 112 38 113 42
rect 98 34 102 38
rect 87 30 88 34
rect 92 30 102 34
rect 118 32 122 48
rect 118 27 122 28
rect 128 60 132 61
rect 128 42 132 56
rect 148 58 150 62
rect 154 58 155 62
rect 128 32 132 38
rect 128 27 132 28
rect 138 42 142 43
rect 89 22 90 24
rect 78 20 90 22
rect 94 22 95 24
rect 138 22 142 38
rect 94 20 142 22
rect 78 18 142 20
rect 148 22 152 58
rect 148 18 150 22
rect 154 18 155 22
rect 148 17 152 18
rect -2 8 18 12
rect 22 8 66 12
rect 70 8 114 12
rect 118 8 138 12
rect 142 8 162 12
rect -2 4 30 8
rect 34 4 42 8
rect 46 4 54 8
rect 58 4 78 8
rect 82 4 90 8
rect 94 4 102 8
rect 106 4 162 8
rect -2 0 162 4
<< ntransistor >>
rect 13 6 15 25
rect 25 15 27 24
rect 37 15 39 29
rect 61 16 63 24
rect 73 15 75 24
rect 85 15 87 26
rect 97 15 99 27
rect 109 15 111 24
rect 121 16 123 24
rect 145 6 147 25
<< ptransistor >>
rect 13 55 15 94
rect 25 65 27 83
rect 37 66 39 84
rect 61 56 63 72
rect 73 56 75 78
rect 85 56 87 78
rect 97 55 99 77
rect 109 55 111 77
rect 121 56 123 78
rect 145 55 147 94
<< polycontact >>
rect 38 58 42 62
rect 20 48 24 52
rect 68 48 72 52
rect 88 48 92 52
rect 28 38 32 42
rect 38 38 42 42
rect 54 38 58 42
rect 118 48 122 52
rect 20 28 24 32
rect 68 28 72 32
rect 88 30 92 34
rect 108 38 112 42
rect 128 38 132 42
rect 138 38 142 42
rect 118 28 122 32
<< ndcontact >>
rect 6 18 10 22
rect 42 18 46 22
rect 54 18 58 22
rect 18 8 22 12
rect 90 20 94 24
rect 128 28 132 32
rect 66 8 70 12
rect 114 8 118 12
rect 138 8 142 12
rect 150 18 154 22
<< pdcontact >>
rect 6 78 10 82
rect 6 68 10 72
rect 6 58 10 62
rect 18 88 22 92
rect 42 88 46 92
rect 66 88 70 92
rect 30 68 34 72
rect 114 88 118 92
rect 54 58 58 62
rect 78 68 82 72
rect 138 88 142 92
rect 138 78 142 82
rect 90 58 94 62
rect 102 68 106 72
rect 102 58 106 62
rect 138 68 142 72
rect 128 56 132 60
rect 150 78 154 82
rect 150 68 154 72
rect 150 58 154 62
<< psubstratepcontact >>
rect 30 4 34 8
rect 42 4 46 8
rect 54 4 58 8
rect 78 4 82 8
rect 90 4 94 8
rect 102 4 106 8
<< nsubstratencontact >>
rect 54 92 58 96
rect 78 92 82 96
rect 90 92 94 96
rect 102 92 106 96
rect 126 92 130 96
<< psubstratepdiff >>
rect 29 8 59 9
rect 29 4 30 8
rect 34 4 42 8
rect 46 4 54 8
rect 58 4 59 8
rect 77 8 107 9
rect 29 3 59 4
rect 77 4 78 8
rect 82 4 90 8
rect 94 4 102 8
rect 106 4 107 8
rect 77 3 107 4
<< nsubstratendiff >>
rect 53 96 59 97
rect 53 92 54 96
rect 58 92 59 96
rect 77 96 107 97
rect 53 86 59 92
rect 77 92 78 96
rect 82 92 90 96
rect 94 92 102 96
rect 106 92 107 96
rect 125 96 131 97
rect 77 91 107 92
rect 125 92 126 96
rect 130 92 131 96
rect 125 86 131 92
<< labels >>
rlabel metal1 20 50 20 50 6 a
rlabel metal1 10 50 10 50 6 cout
rlabel polycontact 40 40 40 40 6 b
rlabel metal1 40 50 40 50 6 b
rlabel polycontact 40 60 40 60 6 b
rlabel metal1 50 70 50 70 6 b
rlabel metal1 60 70 60 70 6 b
rlabel psubstratepcontact 80 6 80 6 6 vss
rlabel metal1 70 45 70 45 6 b
rlabel nsubstratencontact 80 94 80 94 6 vdd
rlabel metal1 150 50 150 50 6 sout
<< end >>
