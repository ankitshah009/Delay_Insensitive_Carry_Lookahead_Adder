magic
tech scmos
timestamp 1179387335
<< checkpaint >>
rect -22 -22 46 94
<< ab >>
rect 0 0 24 72
<< pwell >>
rect -4 -4 28 32
<< nwell >>
rect -4 32 28 76
<< polysilicon >>
rect 12 57 14 61
rect 12 34 14 38
rect 4 33 14 34
rect 4 29 5 33
rect 9 29 14 33
rect 4 28 14 29
rect 12 25 14 28
rect 12 11 14 15
<< ndiffusion >>
rect 3 24 12 25
rect 3 20 5 24
rect 9 20 12 24
rect 3 16 12 20
rect 3 12 5 16
rect 9 15 12 16
rect 14 24 22 25
rect 14 20 17 24
rect 21 20 22 24
rect 14 15 22 20
rect 9 12 10 15
rect 3 8 10 12
rect 3 4 5 8
rect 9 4 10 8
rect 3 3 10 4
<< pdiffusion >>
rect 3 66 10 68
rect 3 62 5 66
rect 9 62 10 66
rect 3 59 10 62
rect 3 55 5 59
rect 9 57 10 59
rect 9 55 12 57
rect 3 52 12 55
rect 3 48 5 52
rect 9 48 12 52
rect 3 38 12 48
rect 14 50 22 57
rect 14 46 17 50
rect 21 46 22 50
rect 14 43 22 46
rect 14 39 17 43
rect 21 39 22 43
rect 14 38 22 39
<< metal1 >>
rect -2 68 26 72
rect -2 66 16 68
rect -2 64 5 66
rect 9 64 16 66
rect 20 64 26 68
rect 5 59 9 62
rect 5 52 9 55
rect 5 47 9 48
rect 17 50 22 59
rect 21 46 22 50
rect 17 43 22 46
rect 2 39 17 43
rect 21 39 22 43
rect 2 37 22 39
rect 4 29 5 33
rect 9 29 10 33
rect 4 24 10 29
rect 4 20 5 24
rect 9 20 10 24
rect 4 16 10 20
rect 4 12 5 16
rect 9 12 10 16
rect 17 24 22 37
rect 21 20 22 24
rect 17 13 22 20
rect 4 8 10 12
rect -2 4 5 8
rect 9 4 16 8
rect 20 4 26 8
rect -2 0 26 4
<< ntransistor >>
rect 12 15 14 25
<< ptransistor >>
rect 12 38 14 57
<< polycontact >>
rect 5 29 9 33
<< ndcontact >>
rect 5 20 9 24
rect 5 12 9 16
rect 17 20 21 24
rect 5 4 9 8
<< pdcontact >>
rect 5 62 9 66
rect 5 55 9 59
rect 5 48 9 52
rect 17 46 21 50
rect 17 39 21 43
<< psubstratepcontact >>
rect 16 4 20 8
<< nsubstratencontact >>
rect 16 64 20 68
<< psubstratepdiff >>
rect 15 8 21 9
rect 15 4 16 8
rect 20 4 21 8
rect 15 3 21 4
<< nsubstratendiff >>
rect 15 68 21 69
rect 15 64 16 68
rect 20 64 21 68
rect 15 63 21 64
<< labels >>
rlabel metal1 4 40 4 40 6 z
rlabel metal1 12 4 12 4 6 vss
rlabel metal1 12 40 12 40 6 z
rlabel metal1 12 68 12 68 6 vdd
rlabel metal1 20 36 20 36 6 z
<< end >>
