magic
tech scmos
timestamp 1179385887
<< checkpaint >>
rect -22 -25 54 105
<< ab >>
rect 0 0 32 80
<< pwell >>
rect -4 -7 36 36
<< nwell >>
rect -4 36 36 87
<< polysilicon >>
rect 9 70 11 74
rect 19 70 21 74
rect 9 39 11 42
rect 19 39 21 42
rect 9 38 21 39
rect 9 34 16 38
rect 20 34 21 38
rect 9 33 21 34
rect 9 30 11 33
rect 19 30 21 33
rect 9 6 11 11
rect 19 6 21 11
<< ndiffusion >>
rect 2 23 9 30
rect 2 19 3 23
rect 7 19 9 23
rect 2 16 9 19
rect 2 12 3 16
rect 7 12 9 16
rect 2 11 9 12
rect 11 29 19 30
rect 11 25 13 29
rect 17 25 19 29
rect 11 22 19 25
rect 11 18 13 22
rect 17 18 19 22
rect 11 11 19 18
rect 21 23 29 30
rect 21 19 23 23
rect 27 19 29 23
rect 21 16 29 19
rect 21 12 23 16
rect 27 12 29 16
rect 21 11 29 12
<< pdiffusion >>
rect 2 69 9 70
rect 2 65 3 69
rect 7 65 9 69
rect 2 62 9 65
rect 2 58 3 62
rect 7 58 9 62
rect 2 42 9 58
rect 11 62 19 70
rect 11 58 13 62
rect 17 58 19 62
rect 11 55 19 58
rect 11 51 13 55
rect 17 51 19 55
rect 11 42 19 51
rect 21 69 29 70
rect 21 65 23 69
rect 27 65 29 69
rect 21 62 29 65
rect 21 58 23 62
rect 27 58 29 62
rect 21 42 29 58
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect -2 69 34 78
rect -2 68 3 69
rect 2 65 3 68
rect 7 68 23 69
rect 7 65 8 68
rect 2 62 8 65
rect 22 65 23 68
rect 27 68 34 69
rect 27 65 28 68
rect 2 58 3 62
rect 7 58 8 62
rect 13 62 17 63
rect 22 62 28 65
rect 22 58 23 62
rect 27 58 28 62
rect 13 55 17 58
rect 2 51 13 54
rect 2 50 17 51
rect 2 30 6 50
rect 26 38 30 47
rect 15 34 16 38
rect 20 34 30 38
rect 2 29 23 30
rect 2 26 13 29
rect 17 26 23 29
rect 2 19 3 23
rect 7 19 8 23
rect 2 16 8 19
rect 13 22 17 25
rect 13 17 17 18
rect 22 19 23 23
rect 27 19 28 23
rect 2 12 3 16
rect 7 12 8 16
rect 22 16 28 19
rect 22 12 23 16
rect 27 12 28 16
rect -2 2 34 12
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
<< ntransistor >>
rect 9 11 11 30
rect 19 11 21 30
<< ptransistor >>
rect 9 42 11 70
rect 19 42 21 70
<< polycontact >>
rect 16 34 20 38
<< ndcontact >>
rect 3 19 7 23
rect 3 12 7 16
rect 13 25 17 29
rect 13 18 17 22
rect 23 19 27 23
rect 23 12 27 16
<< pdcontact >>
rect 3 65 7 69
rect 3 58 7 62
rect 13 58 17 62
rect 13 51 17 55
rect 23 65 27 69
rect 23 58 27 62
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
<< psubstratepdiff >>
rect 0 2 32 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 32 2
rect 0 -3 32 -2
<< nsubstratendiff >>
rect 0 82 32 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 32 82
rect 0 77 32 78
<< labels >>
rlabel metal1 4 40 4 40 6 z
rlabel metal1 12 28 12 28 6 z
rlabel metal1 12 52 12 52 6 z
rlabel metal1 16 6 16 6 6 vss
rlabel metal1 20 36 20 36 6 a
rlabel metal1 20 28 20 28 6 z
rlabel metal1 16 74 16 74 6 vdd
rlabel metal1 28 44 28 44 6 a
<< end >>
