magic
tech scmos
timestamp 1179387461
<< checkpaint >>
rect -22 -22 102 94
<< ab >>
rect 0 0 80 72
<< pwell >>
rect -4 -4 84 32
<< nwell >>
rect -4 32 84 76
<< polysilicon >>
rect 16 59 18 64
rect 26 59 28 64
rect 36 59 38 64
rect 48 59 50 64
rect 58 59 60 64
rect 16 43 18 46
rect 2 42 18 43
rect 2 38 3 42
rect 7 41 18 42
rect 7 38 11 41
rect 2 37 11 38
rect 9 26 11 37
rect 26 35 28 38
rect 16 34 22 35
rect 16 30 17 34
rect 21 30 22 34
rect 16 29 22 30
rect 26 34 32 35
rect 26 30 27 34
rect 31 30 32 34
rect 26 29 32 30
rect 19 26 21 29
rect 26 26 28 29
rect 36 26 38 38
rect 48 35 50 38
rect 58 35 60 38
rect 46 34 54 35
rect 46 30 49 34
rect 53 30 54 34
rect 46 29 54 30
rect 58 34 65 35
rect 58 30 60 34
rect 64 30 65 34
rect 58 29 65 30
rect 46 26 48 29
rect 72 27 78 28
rect 72 24 73 27
rect 69 23 73 24
rect 77 23 78 27
rect 69 22 78 23
rect 69 19 71 22
rect 9 8 11 13
rect 19 8 21 13
rect 26 8 28 13
rect 36 4 38 13
rect 46 8 48 13
rect 69 4 71 8
rect 36 2 71 4
<< ndiffusion >>
rect 2 25 9 26
rect 2 21 3 25
rect 7 21 9 25
rect 2 18 9 21
rect 2 14 3 18
rect 7 14 9 18
rect 2 13 9 14
rect 11 18 19 26
rect 11 14 13 18
rect 17 14 19 18
rect 11 13 19 14
rect 21 13 26 26
rect 28 25 36 26
rect 28 21 30 25
rect 34 21 36 25
rect 28 13 36 21
rect 38 25 46 26
rect 38 21 40 25
rect 44 21 46 25
rect 38 13 46 21
rect 48 19 53 26
rect 48 18 55 19
rect 48 14 50 18
rect 54 14 55 18
rect 48 13 55 14
rect 62 18 69 19
rect 62 14 63 18
rect 67 14 69 18
rect 62 13 69 14
rect 64 8 69 13
rect 71 13 78 19
rect 71 9 73 13
rect 77 9 78 13
rect 71 8 78 9
<< pdiffusion >>
rect 7 68 14 69
rect 7 64 9 68
rect 13 64 14 68
rect 40 68 46 69
rect 40 64 41 68
rect 45 64 46 68
rect 7 59 14 64
rect 40 59 46 64
rect 7 46 16 59
rect 18 58 26 59
rect 18 54 20 58
rect 24 54 26 58
rect 18 51 26 54
rect 18 47 20 51
rect 24 47 26 51
rect 18 46 26 47
rect 21 38 26 46
rect 28 50 36 59
rect 28 46 30 50
rect 34 46 36 50
rect 28 43 36 46
rect 28 39 30 43
rect 34 39 36 43
rect 28 38 36 39
rect 38 38 48 59
rect 50 43 58 59
rect 50 39 52 43
rect 56 39 58 43
rect 50 38 58 39
rect 60 58 67 59
rect 60 54 62 58
rect 66 54 67 58
rect 60 53 67 54
rect 60 38 65 53
<< metal1 >>
rect -2 68 82 72
rect -2 64 9 68
rect 13 64 41 68
rect 45 64 72 68
rect 76 64 82 68
rect 2 54 15 59
rect 19 54 20 58
rect 24 54 62 58
rect 66 54 71 58
rect 2 43 6 54
rect 19 51 24 54
rect 19 50 20 51
rect 10 47 20 50
rect 10 46 24 47
rect 30 50 63 51
rect 34 47 63 50
rect 2 42 7 43
rect 2 38 3 42
rect 2 37 7 38
rect 2 29 6 37
rect 10 26 14 46
rect 30 43 34 46
rect 17 39 30 42
rect 52 43 56 44
rect 17 38 34 39
rect 41 39 52 42
rect 41 38 56 39
rect 17 34 21 38
rect 41 34 45 38
rect 26 30 27 34
rect 31 30 45 34
rect 17 29 21 30
rect 3 25 7 26
rect 10 25 35 26
rect 10 22 30 25
rect 29 21 30 22
rect 34 21 35 25
rect 39 25 45 30
rect 39 21 40 25
rect 44 21 45 25
rect 49 34 54 35
rect 53 30 54 34
rect 59 34 63 47
rect 66 37 78 43
rect 59 30 60 34
rect 64 30 70 34
rect 49 26 54 30
rect 49 22 63 26
rect 3 18 7 21
rect 66 18 70 30
rect 74 28 78 37
rect 73 27 78 28
rect 77 23 78 27
rect 73 21 78 23
rect 12 14 13 18
rect 17 14 50 18
rect 54 14 55 18
rect 62 14 63 18
rect 67 14 70 18
rect 3 8 7 14
rect 73 13 77 14
rect 73 8 77 9
rect -2 0 82 8
<< ntransistor >>
rect 9 13 11 26
rect 19 13 21 26
rect 26 13 28 26
rect 36 13 38 26
rect 46 13 48 26
rect 69 8 71 19
<< ptransistor >>
rect 16 46 18 59
rect 26 38 28 59
rect 36 38 38 59
rect 48 38 50 59
rect 58 38 60 59
<< polycontact >>
rect 3 38 7 42
rect 17 30 21 34
rect 27 30 31 34
rect 49 30 53 34
rect 60 30 64 34
rect 73 23 77 27
<< ndcontact >>
rect 3 21 7 25
rect 3 14 7 18
rect 13 14 17 18
rect 30 21 34 25
rect 40 21 44 25
rect 50 14 54 18
rect 63 14 67 18
rect 73 9 77 13
<< pdcontact >>
rect 9 64 13 68
rect 41 64 45 68
rect 20 54 24 58
rect 20 47 24 51
rect 30 46 34 50
rect 30 39 34 43
rect 52 39 56 43
rect 62 54 66 58
<< nsubstratencontact >>
rect 72 64 76 68
<< nsubstratendiff >>
rect 71 68 77 69
rect 71 64 72 68
rect 76 64 77 68
rect 71 40 77 64
<< labels >>
rlabel polycontact 19 32 19 32 6 a2n
rlabel polycontact 29 32 29 32 6 a1n
rlabel polycontact 61 32 61 32 6 a2n
rlabel metal1 4 44 4 44 6 b
rlabel metal1 20 24 20 24 6 z
rlabel metal1 28 24 28 24 6 z
rlabel metal1 19 35 19 35 6 a2n
rlabel metal1 12 36 12 36 6 z
rlabel metal1 20 48 20 48 6 z
rlabel metal1 28 56 28 56 6 z
rlabel metal1 12 56 12 56 6 b
rlabel metal1 40 4 40 4 6 vss
rlabel metal1 43 31 43 31 6 a1n
rlabel metal1 35 32 35 32 6 a1n
rlabel metal1 32 44 32 44 6 a2n
rlabel metal1 44 56 44 56 6 z
rlabel metal1 36 56 36 56 6 z
rlabel metal1 40 68 40 68 6 vdd
rlabel metal1 60 24 60 24 6 a1
rlabel metal1 52 28 52 28 6 a1
rlabel pdcontact 54 41 54 41 6 a1n
rlabel metal1 60 56 60 56 6 z
rlabel metal1 52 56 52 56 6 z
rlabel ndcontact 66 16 66 16 6 a2n
rlabel metal1 76 32 76 32 6 a2
rlabel metal1 64 32 64 32 6 a2n
rlabel metal1 68 40 68 40 6 a2
rlabel metal1 68 56 68 56 6 z
<< end >>
