.subckt aoi211v5x05 a1 a2 b c vdd vss z
*   SPICE3 file   created from aoi211v5x05.ext -      technology: scmos
m00 w1     c      z      vdd p w=27u  l=2.3636u ad=67.5p    pd=32u      as=163p     ps=68u
m01 n1     b      w1     vdd p w=27u  l=2.3636u ad=121p     pd=46u      as=67.5p    ps=32u
m02 vdd    a1     n1     vdd p w=27u  l=2.3636u ad=108p     pd=35u      as=121p     ps=46u
m03 n1     a2     vdd    vdd p w=27u  l=2.3636u ad=121p     pd=46u      as=108p     ps=35u
m04 z      c      vss    vss n w=6u   l=2.3636u ad=30p      pd=17.1429u as=72p      ps=30.2857u
m05 vss    b      z      vss n w=6u   l=2.3636u ad=72p      pd=30.2857u as=30p      ps=17.1429u
m06 w2     a1     vss    vss n w=9u   l=2.3636u ad=22.5p    pd=14u      as=108p     ps=45.4286u
m07 z      a2     w2     vss n w=9u   l=2.3636u ad=45p      pd=25.7143u as=22.5p    ps=14u
C0  n1     a2     0.145f
C1  vdd    a1     0.021f
C2  vss    b      0.015f
C3  vdd    c      0.017f
C4  z      a2     0.044f
C5  n1     b      0.106f
C6  z      b      0.083f
C7  a2     a1     0.175f
C8  w1     c      0.002f
C9  a1     b      0.101f
C10 a2     c      0.031f
C11 vdd    w1     0.005f
C12 vss    z      0.271f
C13 b      c      0.200f
C14 vdd    a2     0.050f
C15 vss    a1     0.038f
C16 n1     z      0.032f
C17 vss    c      0.030f
C18 n1     a1     0.029f
C19 vdd    b      0.032f
C20 n1     c      0.001f
C21 z      a1     0.139f
C22 w1     b      0.009f
C23 a2     b      0.097f
C24 z      c      0.278f
C25 vdd    n1     0.190f
C26 w2     z      0.010f
C27 a1     c      0.054f
C28 vss    a2     0.014f
C29 w2     a1     0.003f
C30 vdd    z      0.075f
C33 z      vss    0.018f
C34 a2     vss    0.020f
C35 a1     vss    0.025f
C36 b      vss    0.019f
C37 c      vss    0.023f
.ends
