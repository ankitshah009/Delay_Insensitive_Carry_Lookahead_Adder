magic
tech scmos
timestamp 1170759800
<< checkpaint >>
rect -22 -26 54 114
<< ab >>
rect 0 0 32 88
<< pwell >>
rect -4 -8 36 40
<< nwell >>
rect -4 40 36 96
<< polysilicon >>
rect 2 77 11 83
rect 9 74 11 77
rect 21 77 30 83
rect 21 74 23 77
rect 9 43 11 46
rect 21 43 23 46
rect 2 42 14 43
rect 2 38 6 42
rect 10 38 14 42
rect 2 37 14 38
rect 18 42 30 43
rect 18 38 22 42
rect 26 38 30 42
rect 18 37 30 38
rect 9 34 11 37
rect 21 34 23 37
rect 9 11 11 14
rect 2 5 11 11
rect 21 11 23 14
rect 21 5 30 11
<< ndiffusion >>
rect 2 21 9 34
rect 2 17 3 21
rect 7 17 9 21
rect 2 14 9 17
rect 11 14 21 34
rect 23 22 30 34
rect 23 18 25 22
rect 29 18 30 22
rect 23 14 30 18
rect 13 2 19 14
<< pdiffusion >>
rect 13 74 19 86
rect 2 71 9 74
rect 2 67 3 71
rect 7 67 9 71
rect 2 46 9 67
rect 11 51 21 74
rect 11 47 14 51
rect 18 47 21 51
rect 11 46 21 47
rect 23 71 30 74
rect 23 67 25 71
rect 29 67 30 71
rect 23 46 30 67
<< metal1 >>
rect -2 86 2 90
rect 10 86 22 90
rect 30 86 34 90
rect 6 82 10 86
rect 6 71 10 78
rect 2 67 3 71
rect 7 67 10 71
rect 22 82 26 86
rect 22 71 26 78
rect 22 67 25 71
rect 29 67 30 71
rect 14 51 18 55
rect 6 42 10 47
rect 6 33 10 38
rect 14 22 18 47
rect 22 42 26 47
rect 22 33 26 38
rect 2 17 3 21
rect 7 17 10 21
rect 14 18 25 22
rect 29 18 30 22
rect 6 10 10 17
rect 6 2 10 6
rect -2 -2 2 2
rect 10 -2 22 2
rect 30 -2 34 2
<< metal2 >>
rect -2 86 6 90
rect 10 86 22 90
rect 26 86 34 90
rect -2 82 34 86
rect -2 78 6 82
rect 10 78 22 82
rect 26 78 34 82
rect -2 76 34 78
rect -2 10 34 12
rect -2 6 6 10
rect 10 6 34 10
rect -2 2 34 6
rect -2 -2 6 2
rect 10 -2 22 2
rect 26 -2 34 2
<< ntransistor >>
rect 9 14 11 34
rect 21 14 23 34
<< ptransistor >>
rect 9 46 11 74
rect 21 46 23 74
<< polycontact >>
rect 6 38 10 42
rect 22 38 26 42
<< ndcontact >>
rect 3 17 7 21
rect 25 18 29 22
<< pdcontact >>
rect 3 67 7 71
rect 14 47 18 51
rect 25 67 29 71
<< m2contact >>
rect 6 86 10 90
rect 22 86 26 90
rect 6 78 10 82
rect 22 78 26 82
rect 6 6 10 10
rect 6 -2 10 2
rect 22 -2 26 2
<< psubstratepcontact >>
rect 2 -2 6 2
rect 26 -2 30 2
<< nsubstratencontact >>
rect 2 86 6 90
rect 26 86 30 90
<< psubstratepdiff >>
rect 0 2 7 3
rect 25 2 32 3
rect 0 -2 2 2
rect 6 -2 7 2
rect 0 -3 7 -2
rect 25 -2 26 2
rect 30 -2 32 2
rect 25 -3 32 -2
<< nsubstratendiff >>
rect 0 90 7 91
rect 0 86 2 90
rect 6 86 7 90
rect 25 90 32 91
rect 25 86 26 90
rect 30 86 32 90
rect 0 85 7 86
rect 25 85 32 86
<< labels >>
rlabel polycontact 8 40 8 40 6 a
rlabel metal1 16 40 16 40 6 z
rlabel metal1 24 20 24 20 6 z
rlabel polycontact 24 40 24 40 6 b
rlabel metal2 16 6 16 6 6 vss
rlabel metal2 16 82 16 82 6 vdd
<< end >>
