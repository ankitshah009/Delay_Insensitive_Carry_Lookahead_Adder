magic
tech scmos
timestamp 1179386415
<< checkpaint >>
rect -22 -22 94 94
<< ab >>
rect 0 0 72 72
<< pwell >>
rect -4 -4 76 32
<< nwell >>
rect -4 32 76 76
<< polysilicon >>
rect 9 62 11 67
rect 19 62 21 67
rect 29 62 31 67
rect 39 62 41 67
rect 50 52 52 57
rect 60 52 62 57
rect 9 35 11 38
rect 19 35 21 38
rect 29 35 31 38
rect 39 35 41 38
rect 50 35 52 38
rect 60 35 62 38
rect 9 34 15 35
rect 9 30 10 34
rect 14 30 15 34
rect 9 29 15 30
rect 19 34 31 35
rect 19 30 26 34
rect 30 30 31 34
rect 19 29 31 30
rect 12 26 14 29
rect 19 26 21 29
rect 29 26 31 29
rect 36 34 52 35
rect 36 30 42 34
rect 46 33 52 34
rect 56 34 62 35
rect 46 30 47 33
rect 36 29 47 30
rect 56 30 57 34
rect 61 30 62 34
rect 56 29 62 30
rect 36 26 38 29
rect 12 8 14 13
rect 19 8 21 13
rect 29 8 31 13
rect 36 8 38 13
<< ndiffusion >>
rect 3 13 12 26
rect 14 13 19 26
rect 21 18 29 26
rect 21 14 23 18
rect 27 14 29 18
rect 21 13 29 14
rect 31 13 36 26
rect 38 13 47 26
rect 3 8 10 13
rect 40 8 47 13
rect 3 4 5 8
rect 9 4 10 8
rect 3 3 10 4
rect 40 4 41 8
rect 45 4 47 8
rect 40 3 47 4
<< pdiffusion >>
rect 2 61 9 62
rect 2 57 3 61
rect 7 57 9 61
rect 2 38 9 57
rect 11 58 19 62
rect 11 54 13 58
rect 17 54 19 58
rect 11 50 19 54
rect 11 46 13 50
rect 17 46 19 50
rect 11 38 19 46
rect 21 61 29 62
rect 21 57 23 61
rect 27 57 29 61
rect 21 38 29 57
rect 31 58 39 62
rect 31 54 33 58
rect 37 54 39 58
rect 31 50 39 54
rect 31 46 33 50
rect 37 46 39 50
rect 31 38 39 46
rect 41 61 48 62
rect 41 57 43 61
rect 47 57 48 61
rect 41 52 48 57
rect 41 38 50 52
rect 52 50 60 52
rect 52 46 54 50
rect 58 46 60 50
rect 52 38 60 46
rect 62 51 70 52
rect 62 47 64 51
rect 68 47 70 51
rect 62 43 70 47
rect 62 39 64 43
rect 68 39 70 43
rect 62 38 70 39
<< metal1 >>
rect -2 68 74 72
rect -2 64 53 68
rect 57 64 64 68
rect 68 64 74 68
rect 3 61 7 64
rect 23 61 27 64
rect 3 56 7 57
rect 13 58 17 59
rect 43 61 47 64
rect 23 56 27 57
rect 33 58 38 59
rect 13 50 17 54
rect 37 54 38 58
rect 43 56 47 57
rect 33 50 38 54
rect 64 51 68 64
rect 2 46 13 50
rect 17 46 33 50
rect 37 46 54 50
rect 58 46 59 50
rect 2 18 6 46
rect 64 43 68 47
rect 25 38 57 42
rect 64 38 68 39
rect 10 34 21 35
rect 14 30 21 34
rect 25 34 31 38
rect 25 30 26 34
rect 30 30 31 34
rect 41 30 42 34
rect 46 30 47 34
rect 53 30 57 38
rect 61 30 63 34
rect 10 29 21 30
rect 17 26 21 29
rect 41 26 47 30
rect 17 22 47 26
rect 2 14 23 18
rect 27 14 31 18
rect -2 4 5 8
rect 9 4 41 8
rect 45 4 53 8
rect 57 4 64 8
rect 68 4 74 8
rect -2 0 74 4
<< ntransistor >>
rect 12 13 14 26
rect 19 13 21 26
rect 29 13 31 26
rect 36 13 38 26
<< ptransistor >>
rect 9 38 11 62
rect 19 38 21 62
rect 29 38 31 62
rect 39 38 41 62
rect 50 38 52 52
rect 60 38 62 52
<< polycontact >>
rect 10 30 14 34
rect 26 30 30 34
rect 42 30 46 34
rect 57 30 61 34
<< ndcontact >>
rect 23 14 27 18
rect 5 4 9 8
rect 41 4 45 8
<< pdcontact >>
rect 3 57 7 61
rect 13 54 17 58
rect 13 46 17 50
rect 23 57 27 61
rect 33 54 37 58
rect 33 46 37 50
rect 43 57 47 61
rect 54 46 58 50
rect 64 47 68 51
rect 64 39 68 43
<< psubstratepcontact >>
rect 53 4 57 8
rect 64 4 68 8
<< nsubstratencontact >>
rect 53 64 57 68
rect 64 64 68 68
<< psubstratepdiff >>
rect 52 8 69 9
rect 52 4 53 8
rect 57 4 64 8
rect 68 4 69 8
rect 52 3 69 4
<< nsubstratendiff >>
rect 52 68 69 69
rect 52 64 53 68
rect 57 64 64 68
rect 68 64 69 68
rect 52 63 69 64
<< labels >>
rlabel metal1 4 32 4 32 6 z
rlabel metal1 20 16 20 16 6 z
rlabel metal1 12 16 12 16 6 z
rlabel metal1 20 24 20 24 6 a
rlabel polycontact 12 32 12 32 6 a
rlabel metal1 12 48 12 48 6 z
rlabel metal1 20 48 20 48 6 z
rlabel metal1 36 4 36 4 6 vss
rlabel metal1 28 16 28 16 6 z
rlabel metal1 28 24 28 24 6 a
rlabel metal1 36 24 36 24 6 a
rlabel metal1 28 36 28 36 6 b
rlabel metal1 36 40 36 40 6 b
rlabel metal1 28 48 28 48 6 z
rlabel metal1 36 52 36 52 6 z
rlabel metal1 36 68 36 68 6 vdd
rlabel metal1 44 28 44 28 6 a
rlabel metal1 44 40 44 40 6 b
rlabel metal1 52 40 52 40 6 b
rlabel metal1 44 48 44 48 6 z
rlabel metal1 52 48 52 48 6 z
rlabel polycontact 60 32 60 32 6 b
<< end >>
