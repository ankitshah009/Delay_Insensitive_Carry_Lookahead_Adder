magic
tech scmos
timestamp 1180600758
<< checkpaint >>
rect -22 -22 82 122
<< ab >>
rect 0 0 60 100
<< pwell >>
rect -4 -4 64 48
<< nwell >>
rect -4 48 64 104
<< polysilicon >>
rect 11 94 13 98
rect 23 94 25 98
rect 47 75 49 79
rect 11 43 13 55
rect 23 53 25 56
rect 23 52 43 53
rect 23 51 38 52
rect 37 48 38 51
rect 42 48 43 52
rect 37 47 43 48
rect 7 42 13 43
rect 7 38 8 42
rect 12 38 13 42
rect 7 37 13 38
rect 17 42 23 43
rect 17 38 18 42
rect 22 41 23 42
rect 47 41 49 55
rect 22 39 49 41
rect 22 38 25 39
rect 17 37 25 38
rect 11 25 13 37
rect 23 25 25 37
rect 47 25 49 39
rect 47 11 49 15
rect 11 2 13 6
rect 23 2 25 6
<< ndiffusion >>
rect 3 12 11 25
rect 3 8 4 12
rect 8 8 11 12
rect 3 6 11 8
rect 13 6 23 25
rect 25 22 33 25
rect 25 18 28 22
rect 32 18 33 22
rect 25 6 33 18
rect 39 22 47 25
rect 39 18 40 22
rect 44 18 47 22
rect 39 15 47 18
rect 49 22 57 25
rect 49 18 52 22
rect 56 18 57 22
rect 49 15 57 18
<< pdiffusion >>
rect 3 92 11 94
rect 3 88 4 92
rect 8 88 11 92
rect 3 55 11 88
rect 13 56 23 94
rect 25 82 33 94
rect 25 78 28 82
rect 32 78 33 82
rect 25 72 33 78
rect 25 68 28 72
rect 32 68 33 72
rect 25 62 33 68
rect 25 58 28 62
rect 32 58 33 62
rect 25 56 33 58
rect 39 72 47 75
rect 39 68 40 72
rect 44 68 47 72
rect 39 62 47 68
rect 39 58 40 62
rect 44 58 47 62
rect 13 55 18 56
rect 39 55 47 58
rect 49 72 57 75
rect 49 68 52 72
rect 56 68 57 72
rect 49 62 57 68
rect 49 58 52 62
rect 56 58 57 62
rect 49 55 57 58
<< metal1 >>
rect -2 96 62 100
rect -2 92 40 96
rect 44 92 52 96
rect 56 92 62 96
rect -2 88 4 92
rect 8 88 62 92
rect 8 42 12 83
rect 8 17 12 38
rect 18 42 22 83
rect 18 17 22 38
rect 28 82 32 83
rect 28 72 32 78
rect 28 62 32 68
rect 28 22 32 58
rect 40 72 44 73
rect 40 62 44 68
rect 40 52 44 58
rect 52 72 56 88
rect 52 62 56 68
rect 52 57 56 58
rect 37 48 38 52
rect 42 48 44 52
rect 28 17 32 18
rect 40 22 44 48
rect 40 17 44 18
rect 52 22 56 23
rect 52 12 56 18
rect -2 8 4 12
rect 8 8 62 12
rect -2 4 40 8
rect 44 4 52 8
rect 56 4 62 8
rect -2 0 62 4
<< ntransistor >>
rect 11 6 13 25
rect 23 6 25 25
rect 47 15 49 25
<< ptransistor >>
rect 11 55 13 94
rect 23 56 25 94
rect 47 55 49 75
<< polycontact >>
rect 38 48 42 52
rect 8 38 12 42
rect 18 38 22 42
<< ndcontact >>
rect 4 8 8 12
rect 28 18 32 22
rect 40 18 44 22
rect 52 18 56 22
<< pdcontact >>
rect 4 88 8 92
rect 28 78 32 82
rect 28 68 32 72
rect 28 58 32 62
rect 40 68 44 72
rect 40 58 44 62
rect 52 68 56 72
rect 52 58 56 62
<< psubstratepcontact >>
rect 40 4 44 8
rect 52 4 56 8
<< nsubstratencontact >>
rect 40 92 44 96
rect 52 92 56 96
<< psubstratepdiff >>
rect 39 8 57 9
rect 39 4 40 8
rect 44 4 52 8
rect 56 4 57 8
rect 39 3 57 4
<< nsubstratendiff >>
rect 39 96 57 97
rect 39 92 40 96
rect 44 92 52 96
rect 56 92 57 96
rect 39 91 57 92
<< labels >>
rlabel metal1 10 50 10 50 6 i
rlabel metal1 20 50 20 50 6 cmd
rlabel metal1 30 6 30 6 6 vss
rlabel metal1 30 50 30 50 6 nq
rlabel metal1 30 94 30 94 6 vdd
<< end >>
