.subckt nr4_x1 a b c d vdd vss z
*   SPICE3 file   created from nr4_x1.ext -      technology: scmos
m00 w1     d      vdd    vdd p w=39u  l=2.3636u ad=117p     pd=45u      as=312p     ps=94u
m01 w2     b      w1     vdd p w=39u  l=2.3636u ad=117p     pd=45u      as=117p     ps=45u
m02 w3     c      w2     vdd p w=39u  l=2.3636u ad=117p     pd=45u      as=117p     ps=45u
m03 z      a      w3     vdd p w=39u  l=2.3636u ad=195p     pd=49u      as=117p     ps=45u
m04 w4     a      z      vdd p w=39u  l=2.3636u ad=117p     pd=45u      as=195p     ps=49u
m05 w5     c      w4     vdd p w=39u  l=2.3636u ad=117p     pd=45u      as=117p     ps=45u
m06 w6     b      w5     vdd p w=39u  l=2.3636u ad=117p     pd=45u      as=117p     ps=45u
m07 vdd    d      w6     vdd p w=39u  l=2.3636u ad=312p     pd=94u      as=117p     ps=45u
m08 z      d      vss    vss n w=11u  l=2.3636u ad=55p      pd=21u      as=86p      ps=33.5u
m09 vss    b      z      vss n w=11u  l=2.3636u ad=86p      pd=33.5u    as=55p      ps=21u
m10 z      c      vss    vss n w=11u  l=2.3636u ad=55p      pd=21u      as=86p      ps=33.5u
m11 vss    a      z      vss n w=11u  l=2.3636u ad=86p      pd=33.5u    as=55p      ps=21u
C0  w6     vdd    0.011f
C1  z      w3     0.013f
C2  vss    a      0.026f
C3  vdd    d      0.445f
C4  a      b      0.156f
C5  z      w1     0.027f
C6  w4     vdd    0.011f
C7  vss    b      0.145f
C8  c      d      0.179f
C9  z      a      0.263f
C10 w6     d      0.027f
C11 w4     c      0.011f
C12 w3     vdd    0.011f
C13 vss    z      0.243f
C14 z      b      0.167f
C15 w4     d      0.012f
C16 w2     a      0.018f
C17 w1     vdd    0.011f
C18 vdd    a      0.032f
C19 w3     d      0.012f
C20 vdd    b      0.010f
C21 w1     d      0.012f
C22 a      c      0.339f
C23 vss    c      0.037f
C24 z      w2     0.013f
C25 w5     vdd    0.011f
C26 a      d      0.133f
C27 c      b      0.379f
C28 z      vdd    0.094f
C29 vss    d      0.025f
C30 b      d      0.161f
C31 z      c      0.112f
C32 w2     vdd    0.011f
C33 w5     d      0.028f
C34 z      d      0.431f
C35 w2     d      0.012f
C36 vdd    c      0.014f
C38 z      vss    0.015f
C40 a      vss    0.043f
C41 c      vss    0.050f
C42 b      vss    0.065f
C43 d      vss    0.050f
.ends
