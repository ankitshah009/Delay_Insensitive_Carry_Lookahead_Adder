magic
tech scmos
timestamp 1179386724
<< checkpaint >>
rect -22 -22 54 94
<< ab >>
rect 0 0 32 72
<< pwell >>
rect -4 -4 36 32
<< nwell >>
rect -4 32 36 76
<< polysilicon >>
rect 12 66 14 70
rect 19 66 21 70
rect 12 43 14 46
rect 9 42 15 43
rect 9 38 10 42
rect 14 38 15 42
rect 9 37 15 38
rect 10 25 12 37
rect 19 34 21 46
rect 19 33 25 34
rect 19 29 20 33
rect 24 29 25 33
rect 19 28 25 29
rect 20 25 22 28
rect 10 14 12 19
rect 20 14 22 19
<< ndiffusion >>
rect 2 24 10 25
rect 2 20 3 24
rect 7 20 10 24
rect 2 19 10 20
rect 12 24 20 25
rect 12 20 14 24
rect 18 20 20 24
rect 12 19 20 20
rect 22 24 30 25
rect 22 20 25 24
rect 29 20 30 24
rect 22 19 30 20
<< pdiffusion >>
rect 7 60 12 66
rect 5 59 12 60
rect 5 55 6 59
rect 10 55 12 59
rect 5 54 12 55
rect 7 46 12 54
rect 14 46 19 66
rect 21 65 30 66
rect 21 61 25 65
rect 29 61 30 65
rect 21 58 30 61
rect 21 54 25 58
rect 29 54 30 58
rect 21 46 30 54
<< metal1 >>
rect -2 65 34 72
rect -2 64 25 65
rect 29 64 34 65
rect 2 33 6 59
rect 10 55 11 59
rect 25 58 29 61
rect 25 53 29 54
rect 18 46 22 51
rect 10 42 22 46
rect 10 37 14 38
rect 26 35 30 43
rect 18 33 30 35
rect 2 29 14 33
rect 18 29 20 33
rect 24 29 30 33
rect 3 24 7 25
rect 10 20 14 29
rect 25 24 29 25
rect 18 20 19 24
rect 3 8 7 20
rect 25 8 29 20
rect -2 4 4 8
rect 8 4 24 8
rect 28 4 34 8
rect -2 0 34 4
<< ntransistor >>
rect 10 19 12 25
rect 20 19 22 25
<< ptransistor >>
rect 12 46 14 66
rect 19 46 21 66
<< polycontact >>
rect 10 38 14 42
rect 20 29 24 33
<< ndcontact >>
rect 3 20 7 24
rect 14 20 18 24
rect 25 20 29 24
<< pdcontact >>
rect 6 55 10 59
rect 25 61 29 65
rect 25 54 29 58
<< psubstratepcontact >>
rect 4 4 8 8
rect 24 4 28 8
<< psubstratepdiff >>
rect 3 8 29 9
rect 3 4 4 8
rect 8 4 24 8
rect 28 4 29 8
rect 3 3 29 4
<< labels >>
rlabel metal1 4 44 4 44 6 z
rlabel metal1 12 24 12 24 6 z
rlabel polycontact 12 40 12 40 6 b
rlabel metal1 16 4 16 4 6 vss
rlabel metal1 20 32 20 32 6 a
rlabel metal1 20 48 20 48 6 b
rlabel metal1 16 68 16 68 6 vdd
rlabel metal1 28 36 28 36 6 a
<< end >>
