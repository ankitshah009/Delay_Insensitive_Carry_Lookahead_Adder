.subckt oai21v0x2 a1 a2 b vdd vss z
*   SPICE3 file   created from oai21v0x2.ext -      technology: scmos
m00 vdd    b      z      vdd p w=28u  l=2.3636u ad=177.333p pd=50u      as=134.333p ps=48u
m01 w1     a1     vdd    vdd p w=28u  l=2.3636u ad=70p      pd=33u      as=177.333p ps=50u
m02 z      a2     w1     vdd p w=28u  l=2.3636u ad=134.333p pd=48u      as=70p      ps=33u
m03 w2     a2     z      vdd p w=28u  l=2.3636u ad=70p      pd=33u      as=134.333p ps=48u
m04 vdd    a1     w2     vdd p w=28u  l=2.3636u ad=177.333p pd=50u      as=70p      ps=33u
m05 z      b      n1     vss n w=18u  l=2.3636u ad=90p      pd=32.4u    as=90p      ps=41.1429u
m06 n1     b      z      vss n w=12u  l=2.3636u ad=60p      pd=27.4286u as=60p      ps=21.6u
m07 vss    a2     n1     vss n w=20u  l=2.3636u ad=140p     pd=34u      as=100p     ps=45.7143u
m08 n1     a1     vss    vss n w=20u  l=2.3636u ad=100p     pd=45.7143u as=140p     ps=34u
C0  a1     b      0.145f
C1  a2     vdd    0.029f
C2  vss    z      0.047f
C3  b      vdd    0.058f
C4  n1     a2     0.032f
C5  vss    a1     0.102f
C6  n1     b      0.035f
C7  w2     vdd    0.005f
C8  z      a1     0.068f
C9  vss    n1     0.339f
C10 a2     b      0.066f
C11 z      vdd    0.264f
C12 a1     vdd    0.061f
C13 vss    a2     0.020f
C14 n1     z      0.217f
C15 w2     a2     0.020f
C16 n1     a1     0.272f
C17 w1     z      0.010f
C18 vss    b      0.024f
C19 n1     vdd    0.008f
C20 z      a2     0.113f
C21 z      b      0.256f
C22 a2     a1     0.285f
C23 w1     vdd    0.005f
C25 z      vss    0.010f
C26 a2     vss    0.027f
C27 a1     vss    0.036f
C28 b      vss    0.023f
.ends
