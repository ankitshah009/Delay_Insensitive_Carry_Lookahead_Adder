magic
tech scmos
timestamp 1179385016
<< checkpaint >>
rect -22 -25 62 105
<< ab >>
rect 0 0 40 80
<< pwell >>
rect -4 -7 44 36
<< nwell >>
rect -4 36 44 87
<< polysilicon >>
rect 9 70 11 74
rect 19 67 21 72
rect 29 67 31 72
rect 9 39 11 42
rect 19 39 21 50
rect 29 47 31 50
rect 29 46 35 47
rect 29 42 30 46
rect 34 42 35 46
rect 29 41 35 42
rect 9 38 15 39
rect 9 34 10 38
rect 14 34 15 38
rect 9 33 15 34
rect 19 38 25 39
rect 19 34 20 38
rect 24 34 25 38
rect 19 33 25 34
rect 9 30 11 33
rect 22 30 24 33
rect 29 30 31 41
rect 9 11 11 16
rect 22 11 24 16
rect 29 11 31 16
<< ndiffusion >>
rect 2 29 9 30
rect 2 25 3 29
rect 7 25 9 29
rect 2 21 9 25
rect 2 17 3 21
rect 7 17 9 21
rect 2 16 9 17
rect 11 16 22 30
rect 24 16 29 30
rect 31 22 36 30
rect 31 21 38 22
rect 31 17 33 21
rect 37 17 38 21
rect 31 16 38 17
rect 13 12 20 16
rect 13 8 14 12
rect 18 8 20 12
rect 13 7 20 8
<< pdiffusion >>
rect 4 63 9 70
rect 2 62 9 63
rect 2 58 3 62
rect 7 58 9 62
rect 2 55 9 58
rect 2 51 3 55
rect 7 51 9 55
rect 2 50 9 51
rect 4 42 9 50
rect 11 67 17 70
rect 11 66 19 67
rect 11 62 13 66
rect 17 62 19 66
rect 11 50 19 62
rect 21 62 29 67
rect 21 58 23 62
rect 27 58 29 62
rect 21 55 29 58
rect 21 51 23 55
rect 27 51 29 55
rect 21 50 29 51
rect 31 66 38 67
rect 31 62 33 66
rect 37 62 38 66
rect 31 50 38 62
rect 11 42 17 50
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect -2 68 42 78
rect 13 66 17 68
rect 2 62 7 63
rect 2 58 3 62
rect 33 66 37 68
rect 13 61 17 62
rect 23 62 27 63
rect 2 55 7 58
rect 2 51 3 55
rect 33 61 37 62
rect 23 55 27 58
rect 2 50 7 51
rect 10 51 23 54
rect 10 50 27 51
rect 2 30 6 50
rect 10 38 14 50
rect 25 42 30 46
rect 34 42 38 55
rect 17 34 20 38
rect 24 34 31 38
rect 10 30 14 34
rect 2 29 7 30
rect 2 25 3 29
rect 10 26 22 30
rect 2 23 7 25
rect 2 21 14 23
rect 2 17 3 21
rect 7 17 14 21
rect 18 21 22 26
rect 26 25 31 34
rect 18 17 33 21
rect 37 17 38 21
rect -2 8 14 12
rect 18 8 42 12
rect -2 2 42 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
<< ntransistor >>
rect 9 16 11 30
rect 22 16 24 30
rect 29 16 31 30
<< ptransistor >>
rect 9 42 11 70
rect 19 50 21 67
rect 29 50 31 67
<< polycontact >>
rect 30 42 34 46
rect 10 34 14 38
rect 20 34 24 38
<< ndcontact >>
rect 3 25 7 29
rect 3 17 7 21
rect 33 17 37 21
rect 14 8 18 12
<< pdcontact >>
rect 3 58 7 62
rect 3 51 7 55
rect 13 62 17 66
rect 23 58 27 62
rect 23 51 27 55
rect 33 62 37 66
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
<< psubstratepdiff >>
rect 0 2 40 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 40 2
rect 0 -3 40 -2
<< nsubstratendiff >>
rect 0 82 40 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 40 82
rect 0 77 40 78
<< labels >>
rlabel polycontact 12 36 12 36 6 zn
rlabel metal1 4 40 4 40 6 z
rlabel metal1 12 20 12 20 6 z
rlabel metal1 12 40 12 40 6 zn
rlabel metal1 20 6 20 6 6 vss
rlabel metal1 20 36 20 36 6 a
rlabel metal1 28 32 28 32 6 a
rlabel metal1 28 44 28 44 6 b
rlabel metal1 25 56 25 56 6 zn
rlabel metal1 20 74 20 74 6 vdd
rlabel metal1 28 19 28 19 6 zn
rlabel metal1 36 52 36 52 6 b
<< end >>
