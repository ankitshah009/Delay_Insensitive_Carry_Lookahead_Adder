magic
tech scmos
timestamp 1179385595
<< checkpaint >>
rect -22 -22 78 94
<< ab >>
rect 0 0 56 72
<< pwell >>
rect -4 -4 60 32
<< nwell >>
rect -4 32 60 76
<< polysilicon >>
rect 9 66 11 70
rect 19 66 21 70
rect 29 66 31 70
rect 39 66 41 70
rect 9 35 11 38
rect 19 35 21 38
rect 29 35 31 38
rect 39 35 41 38
rect 9 34 24 35
rect 9 30 12 34
rect 16 30 19 34
rect 23 30 24 34
rect 9 29 24 30
rect 29 34 41 35
rect 29 30 36 34
rect 40 30 41 34
rect 29 29 41 30
rect 9 26 11 29
rect 19 26 21 29
rect 29 26 31 29
rect 39 26 41 29
rect 9 7 11 12
rect 19 7 21 12
rect 39 11 41 16
rect 29 3 31 8
<< ndiffusion >>
rect 2 17 9 26
rect 2 13 3 17
rect 7 13 9 17
rect 2 12 9 13
rect 11 25 19 26
rect 11 21 13 25
rect 17 21 19 25
rect 11 18 19 21
rect 11 14 13 18
rect 17 14 19 18
rect 11 12 19 14
rect 21 17 29 26
rect 21 13 23 17
rect 27 13 29 17
rect 21 12 29 13
rect 23 8 29 12
rect 31 25 39 26
rect 31 21 33 25
rect 37 21 39 25
rect 31 16 39 21
rect 41 21 48 26
rect 41 17 43 21
rect 47 17 48 21
rect 41 16 48 17
rect 31 8 36 16
<< pdiffusion >>
rect 2 65 9 66
rect 2 61 3 65
rect 7 61 9 65
rect 2 58 9 61
rect 2 54 3 58
rect 7 54 9 58
rect 2 38 9 54
rect 11 58 19 66
rect 11 54 13 58
rect 17 54 19 58
rect 11 51 19 54
rect 11 47 13 51
rect 17 47 19 51
rect 11 38 19 47
rect 21 65 29 66
rect 21 61 23 65
rect 27 61 29 65
rect 21 58 29 61
rect 21 54 23 58
rect 27 54 29 58
rect 21 38 29 54
rect 31 50 39 66
rect 31 46 33 50
rect 37 46 39 50
rect 31 43 39 46
rect 31 39 33 43
rect 37 39 39 43
rect 31 38 39 39
rect 41 65 48 66
rect 41 61 43 65
rect 47 61 48 65
rect 41 58 48 61
rect 41 54 43 58
rect 47 54 48 58
rect 41 38 48 54
<< metal1 >>
rect -2 65 58 72
rect -2 64 3 65
rect 2 61 3 64
rect 7 64 23 65
rect 7 61 8 64
rect 2 58 8 61
rect 27 64 43 65
rect 2 54 3 58
rect 7 54 8 58
rect 13 58 17 59
rect 13 51 17 54
rect 23 58 27 61
rect 42 61 43 64
rect 47 64 58 65
rect 47 61 48 64
rect 42 58 48 61
rect 42 54 43 58
rect 47 54 48 58
rect 23 53 27 54
rect 2 47 13 51
rect 33 50 37 51
rect 17 47 23 50
rect 2 46 23 47
rect 2 26 6 46
rect 33 43 37 46
rect 23 39 33 42
rect 23 38 37 39
rect 11 30 12 34
rect 16 30 19 34
rect 2 25 17 26
rect 2 21 13 25
rect 23 25 27 38
rect 42 34 46 51
rect 33 30 36 34
rect 40 30 46 34
rect 23 21 33 25
rect 37 21 38 25
rect 43 21 47 22
rect 13 18 17 21
rect 2 13 3 17
rect 7 13 8 17
rect 13 13 17 14
rect 22 13 23 17
rect 27 13 28 17
rect 2 8 8 13
rect 22 8 28 13
rect 43 8 47 17
rect -2 4 41 8
rect 45 4 48 8
rect 52 4 58 8
rect -2 0 58 4
<< ntransistor >>
rect 9 12 11 26
rect 19 12 21 26
rect 29 8 31 26
rect 39 16 41 26
<< ptransistor >>
rect 9 38 11 66
rect 19 38 21 66
rect 29 38 31 66
rect 39 38 41 66
<< polycontact >>
rect 12 30 16 34
rect 19 30 23 34
rect 36 30 40 34
<< ndcontact >>
rect 3 13 7 17
rect 13 21 17 25
rect 13 14 17 18
rect 23 13 27 17
rect 33 21 37 25
rect 43 17 47 21
<< pdcontact >>
rect 3 61 7 65
rect 3 54 7 58
rect 13 54 17 58
rect 13 47 17 51
rect 23 61 27 65
rect 23 54 27 58
rect 33 46 37 50
rect 33 39 37 43
rect 43 61 47 65
rect 43 54 47 58
<< psubstratepcontact >>
rect 41 4 45 8
rect 48 4 52 8
<< psubstratepdiff >>
rect 40 8 53 9
rect 40 4 41 8
rect 45 4 48 8
rect 52 4 53 8
rect 40 3 53 4
<< labels >>
rlabel polysilicon 16 32 16 32 6 an
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 24 12 24 6 z
rlabel metal1 19 32 19 32 6 an
rlabel metal1 12 48 12 48 6 z
rlabel metal1 20 48 20 48 6 z
rlabel metal1 28 4 28 4 6 vss
rlabel metal1 30 23 30 23 6 an
rlabel metal1 36 32 36 32 6 a
rlabel metal1 35 44 35 44 6 an
rlabel metal1 28 68 28 68 6 vdd
rlabel metal1 44 44 44 44 6 a
<< end >>
