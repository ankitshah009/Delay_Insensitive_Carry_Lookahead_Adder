magic
tech scmos
timestamp 1179387273
<< checkpaint >>
rect -22 -25 86 105
<< ab >>
rect 0 0 64 80
<< pwell >>
rect -4 -7 68 36
<< nwell >>
rect -4 36 68 87
<< polysilicon >>
rect 28 70 30 74
rect 35 70 37 74
rect 42 70 44 74
rect 49 70 51 74
rect 9 61 11 65
rect 9 40 11 49
rect 28 40 30 43
rect 9 39 15 40
rect 9 35 10 39
rect 14 35 15 39
rect 9 34 15 35
rect 19 39 30 40
rect 19 35 20 39
rect 24 38 30 39
rect 24 35 25 38
rect 19 34 25 35
rect 35 34 37 43
rect 9 25 11 34
rect 19 25 21 34
rect 29 33 37 34
rect 29 29 32 33
rect 36 29 37 33
rect 29 28 37 29
rect 42 31 44 43
rect 49 40 51 43
rect 49 39 58 40
rect 49 38 53 39
rect 52 35 53 38
rect 57 35 58 39
rect 52 34 58 35
rect 42 30 48 31
rect 29 25 31 28
rect 42 26 43 30
rect 47 26 48 30
rect 42 25 48 26
rect 42 22 44 25
rect 52 22 54 34
rect 9 15 11 19
rect 19 15 21 19
rect 29 14 31 19
rect 42 11 44 16
rect 52 11 54 16
<< ndiffusion >>
rect 2 24 9 25
rect 2 20 3 24
rect 7 20 9 24
rect 2 19 9 20
rect 11 19 19 25
rect 21 24 29 25
rect 21 20 23 24
rect 27 20 29 24
rect 21 19 29 20
rect 31 22 40 25
rect 31 19 42 22
rect 13 13 17 19
rect 33 16 42 19
rect 44 21 52 22
rect 44 17 46 21
rect 50 17 52 21
rect 44 16 52 17
rect 54 16 62 22
rect 13 12 19 13
rect 13 8 14 12
rect 18 8 19 12
rect 13 7 19 8
rect 33 12 40 16
rect 33 8 34 12
rect 38 8 40 12
rect 56 12 62 16
rect 33 7 40 8
rect 56 8 57 12
rect 61 8 62 12
rect 56 7 62 8
<< pdiffusion >>
rect 13 64 19 65
rect 13 61 14 64
rect 4 55 9 61
rect 2 54 9 55
rect 2 50 3 54
rect 7 50 9 54
rect 2 49 9 50
rect 11 60 14 61
rect 18 60 19 64
rect 11 59 19 60
rect 11 49 17 59
rect 23 55 28 70
rect 21 54 28 55
rect 21 50 22 54
rect 26 50 28 54
rect 21 49 28 50
rect 23 43 28 49
rect 30 43 35 70
rect 37 43 42 70
rect 44 43 49 70
rect 51 69 59 70
rect 51 65 53 69
rect 57 65 59 69
rect 51 62 59 65
rect 51 58 53 62
rect 57 58 59 62
rect 51 43 59 58
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect -2 69 66 78
rect -2 68 53 69
rect 14 64 18 68
rect 52 65 53 68
rect 57 68 66 69
rect 57 65 58 68
rect 14 59 18 60
rect 2 54 7 55
rect 2 50 3 54
rect 2 49 7 50
rect 11 50 22 54
rect 26 50 27 54
rect 2 25 6 49
rect 11 40 15 50
rect 34 46 38 63
rect 52 62 58 65
rect 52 58 53 62
rect 57 58 58 62
rect 10 39 15 40
rect 14 35 15 39
rect 10 34 15 35
rect 20 42 38 46
rect 42 46 46 55
rect 42 42 57 46
rect 20 39 24 42
rect 53 39 57 42
rect 20 34 24 35
rect 32 34 47 38
rect 53 34 57 35
rect 11 30 15 34
rect 32 33 38 34
rect 11 26 27 30
rect 2 24 7 25
rect 2 20 3 24
rect 23 24 27 26
rect 36 29 38 33
rect 32 25 38 29
rect 42 26 43 30
rect 47 26 62 30
rect 7 20 16 22
rect 2 17 16 20
rect 27 20 46 21
rect 23 17 46 20
rect 50 17 51 21
rect 58 17 62 26
rect -2 8 14 12
rect 18 8 34 12
rect 38 8 57 12
rect 61 8 66 12
rect -2 2 66 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
<< ntransistor >>
rect 9 19 11 25
rect 19 19 21 25
rect 29 19 31 25
rect 42 16 44 22
rect 52 16 54 22
<< ptransistor >>
rect 9 49 11 61
rect 28 43 30 70
rect 35 43 37 70
rect 42 43 44 70
rect 49 43 51 70
<< polycontact >>
rect 10 35 14 39
rect 20 35 24 39
rect 32 29 36 33
rect 53 35 57 39
rect 43 26 47 30
<< ndcontact >>
rect 3 20 7 24
rect 23 20 27 24
rect 46 17 50 21
rect 14 8 18 12
rect 34 8 38 12
rect 57 8 61 12
<< pdcontact >>
rect 3 50 7 54
rect 14 60 18 64
rect 22 50 26 54
rect 53 65 57 69
rect 53 58 57 62
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
<< psubstratepdiff >>
rect 0 2 64 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 64 2
rect 0 -3 64 -2
<< nsubstratendiff >>
rect 0 82 64 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 64 82
rect 0 77 64 78
<< labels >>
rlabel polycontact 12 37 12 37 6 zn
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 20 12 20 6 z
rlabel metal1 13 40 13 40 6 zn
rlabel metal1 32 6 32 6 6 vss
rlabel ndcontact 25 23 25 23 6 zn
rlabel metal1 36 32 36 32 6 c
rlabel metal1 28 44 28 44 6 d
rlabel metal1 19 52 19 52 6 zn
rlabel metal1 36 56 36 56 6 d
rlabel metal1 32 74 32 74 6 vdd
rlabel metal1 37 19 37 19 6 zn
rlabel metal1 44 36 44 36 6 c
rlabel metal1 44 52 44 52 6 a
rlabel metal1 52 28 52 28 6 b
rlabel metal1 60 20 60 20 6 b
rlabel metal1 52 44 52 44 6 a
<< end >>
