magic
tech scmos
timestamp 1179386339
<< checkpaint >>
rect -22 -25 118 105
<< ab >>
rect 0 0 96 80
<< pwell >>
rect -4 -7 100 36
<< nwell >>
rect -4 36 100 87
<< polysilicon >>
rect 9 68 11 73
rect 19 68 21 73
rect 29 68 31 73
rect 39 68 41 73
rect 49 68 51 73
rect 59 68 61 73
rect 69 60 71 65
rect 79 60 81 65
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 39 39 41 42
rect 9 38 15 39
rect 9 34 10 38
rect 14 34 15 38
rect 9 33 15 34
rect 19 38 31 39
rect 19 34 26 38
rect 30 34 31 38
rect 19 33 31 34
rect 35 38 41 39
rect 35 34 36 38
rect 40 35 41 38
rect 49 35 51 42
rect 59 39 61 42
rect 69 39 71 42
rect 79 39 81 42
rect 59 38 71 39
rect 40 34 54 35
rect 35 33 54 34
rect 12 30 14 33
rect 19 30 21 33
rect 29 30 31 33
rect 36 30 38 33
rect 52 30 54 33
rect 59 34 60 38
rect 64 34 71 38
rect 59 33 71 34
rect 75 38 81 39
rect 75 34 76 38
rect 80 34 81 38
rect 75 33 81 34
rect 59 30 61 33
rect 69 30 71 33
rect 76 30 78 33
rect 12 6 14 10
rect 19 6 21 10
rect 29 6 31 10
rect 36 6 38 10
rect 52 6 54 10
rect 59 6 61 10
rect 69 6 71 10
rect 76 6 78 10
<< ndiffusion >>
rect 3 15 12 30
rect 3 11 5 15
rect 9 11 12 15
rect 3 10 12 11
rect 14 10 19 30
rect 21 22 29 30
rect 21 18 23 22
rect 27 18 29 22
rect 21 10 29 18
rect 31 10 36 30
rect 38 15 52 30
rect 38 11 43 15
rect 47 11 52 15
rect 38 10 52 11
rect 54 10 59 30
rect 61 22 69 30
rect 61 18 63 22
rect 67 18 69 22
rect 61 10 69 18
rect 71 10 76 30
rect 78 22 86 30
rect 78 18 80 22
rect 84 18 86 22
rect 78 15 86 18
rect 78 11 80 15
rect 84 11 86 15
rect 78 10 86 11
<< pdiffusion >>
rect 2 67 9 68
rect 2 63 3 67
rect 7 63 9 67
rect 2 42 9 63
rect 11 61 19 68
rect 11 57 13 61
rect 17 57 19 61
rect 11 54 19 57
rect 11 50 13 54
rect 17 50 19 54
rect 11 42 19 50
rect 21 67 29 68
rect 21 63 23 67
rect 27 63 29 67
rect 21 42 29 63
rect 31 62 39 68
rect 31 58 33 62
rect 37 58 39 62
rect 31 54 39 58
rect 31 50 33 54
rect 37 50 39 54
rect 31 42 39 50
rect 41 67 49 68
rect 41 63 43 67
rect 47 63 49 67
rect 41 42 49 63
rect 51 54 59 68
rect 51 50 53 54
rect 57 50 59 54
rect 51 47 59 50
rect 51 43 53 47
rect 57 43 59 47
rect 51 42 59 43
rect 61 60 67 68
rect 61 59 69 60
rect 61 55 63 59
rect 67 55 69 59
rect 61 42 69 55
rect 71 54 79 60
rect 71 50 73 54
rect 77 50 79 54
rect 71 47 79 50
rect 71 43 73 47
rect 77 43 79 47
rect 71 42 79 43
rect 81 59 88 60
rect 81 55 83 59
rect 87 55 88 59
rect 81 42 88 55
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect -2 68 98 78
rect 3 67 7 68
rect 3 62 7 63
rect 23 67 27 68
rect 43 67 47 68
rect 23 62 27 63
rect 33 62 38 63
rect 43 62 47 63
rect 13 61 17 62
rect 13 55 17 57
rect 2 54 17 55
rect 37 58 38 62
rect 33 54 38 58
rect 63 59 67 68
rect 83 59 87 68
rect 63 54 67 55
rect 73 54 79 55
rect 83 54 87 55
rect 2 50 13 54
rect 17 50 33 54
rect 37 50 53 54
rect 57 50 58 54
rect 2 22 6 50
rect 53 47 58 50
rect 25 42 49 46
rect 57 46 58 47
rect 77 50 79 54
rect 73 47 79 50
rect 57 43 73 46
rect 77 43 79 47
rect 53 42 79 43
rect 10 38 14 39
rect 25 38 31 42
rect 45 38 49 42
rect 25 34 26 38
rect 30 34 31 38
rect 35 34 36 38
rect 40 34 41 38
rect 45 34 60 38
rect 64 34 65 38
rect 75 34 76 38
rect 80 34 81 38
rect 10 30 14 34
rect 35 30 41 34
rect 75 30 81 34
rect 10 26 87 30
rect 2 18 23 22
rect 27 18 63 22
rect 67 18 71 22
rect 79 18 80 22
rect 84 18 85 22
rect 79 15 85 18
rect 4 12 5 15
rect -2 11 5 12
rect 9 12 10 15
rect 42 12 43 15
rect 9 11 43 12
rect 47 12 48 15
rect 79 12 80 15
rect 47 11 80 12
rect 84 12 85 15
rect 84 11 98 12
rect -2 2 98 11
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
<< ntransistor >>
rect 12 10 14 30
rect 19 10 21 30
rect 29 10 31 30
rect 36 10 38 30
rect 52 10 54 30
rect 59 10 61 30
rect 69 10 71 30
rect 76 10 78 30
<< ptransistor >>
rect 9 42 11 68
rect 19 42 21 68
rect 29 42 31 68
rect 39 42 41 68
rect 49 42 51 68
rect 59 42 61 68
rect 69 42 71 60
rect 79 42 81 60
<< polycontact >>
rect 10 34 14 38
rect 26 34 30 38
rect 36 34 40 38
rect 60 34 64 38
rect 76 34 80 38
<< ndcontact >>
rect 5 11 9 15
rect 23 18 27 22
rect 43 11 47 15
rect 63 18 67 22
rect 80 18 84 22
rect 80 11 84 15
<< pdcontact >>
rect 3 63 7 67
rect 13 57 17 61
rect 13 50 17 54
rect 23 63 27 67
rect 33 58 37 62
rect 33 50 37 54
rect 43 63 47 67
rect 53 50 57 54
rect 53 43 57 47
rect 63 55 67 59
rect 73 50 77 54
rect 73 43 77 47
rect 83 55 87 59
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
rect 90 -2 94 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
rect 90 78 94 82
<< psubstratepdiff >>
rect 0 2 96 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 96 2
rect 0 -3 96 -2
<< nsubstratendiff >>
rect 0 82 96 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 96 82
rect 0 77 96 78
<< labels >>
rlabel metal1 12 20 12 20 6 z
rlabel metal1 4 40 4 40 6 z
rlabel polycontact 12 36 12 36 6 a
rlabel metal1 12 52 12 52 6 z
rlabel metal1 20 20 20 20 6 z
rlabel metal1 20 28 20 28 6 a
rlabel metal1 28 20 28 20 6 z
rlabel metal1 28 28 28 28 6 a
rlabel polycontact 28 36 28 36 6 b
rlabel metal1 28 40 28 40 6 b
rlabel metal1 28 52 28 52 6 z
rlabel metal1 20 52 20 52 6 z
rlabel metal1 48 6 48 6 6 vss
rlabel metal1 36 20 36 20 6 z
rlabel metal1 36 28 36 28 6 a
rlabel metal1 44 20 44 20 6 z
rlabel metal1 44 28 44 28 6 a
rlabel metal1 52 20 52 20 6 z
rlabel metal1 52 28 52 28 6 a
rlabel metal1 36 44 36 44 6 b
rlabel metal1 44 44 44 44 6 b
rlabel metal1 52 36 52 36 6 b
rlabel metal1 44 52 44 52 6 z
rlabel metal1 52 52 52 52 6 z
rlabel metal1 36 56 36 56 6 z
rlabel metal1 48 74 48 74 6 vdd
rlabel metal1 60 20 60 20 6 z
rlabel metal1 60 28 60 28 6 a
rlabel metal1 68 20 68 20 6 z
rlabel metal1 68 28 68 28 6 a
rlabel metal1 76 28 76 28 6 a
rlabel metal1 60 36 60 36 6 b
rlabel metal1 60 44 60 44 6 z
rlabel metal1 68 44 68 44 6 z
rlabel metal1 76 48 76 48 6 z
rlabel metal1 84 28 84 28 6 a
<< end >>
