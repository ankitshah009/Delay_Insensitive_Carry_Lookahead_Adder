.subckt nd4v0x3 a b c d vdd vss z
*   SPICE3 file   created from nd4v0x3.ext -      technology: scmos
m00 z      a      vdd    vdd p w=18u  l=2.3636u ad=72p      pd=27u      as=100.688p ps=35.4375u
m01 vdd    b      z      vdd p w=18u  l=2.3636u ad=100.688p pd=35.4375u as=72p      ps=27u
m02 z      c      vdd    vdd p w=16u  l=2.3636u ad=64p      pd=24u      as=89.5p    ps=31.5u
m03 vdd    d      z      vdd p w=16u  l=2.3636u ad=89.5p    pd=31.5u    as=64p      ps=24u
m04 z      d      vdd    vdd p w=16u  l=2.3636u ad=64p      pd=24u      as=89.5p    ps=31.5u
m05 vdd    c      z      vdd p w=16u  l=2.3636u ad=89.5p    pd=31.5u    as=64p      ps=24u
m06 z      b      vdd    vdd p w=14u  l=2.3636u ad=56p      pd=21u      as=78.3125p ps=27.5625u
m07 vdd    a      z      vdd p w=14u  l=2.3636u ad=78.3125p pd=27.5625u as=56p      ps=21u
m08 w1     a      vss    vss n w=19u  l=2.3636u ad=47.5p    pd=24u      as=168.5p   ps=57u
m09 w2     b      w1     vss n w=19u  l=2.3636u ad=47.5p    pd=24u      as=47.5p    ps=24u
m10 w3     c      w2     vss n w=19u  l=2.3636u ad=47.5p    pd=24u      as=47.5p    ps=24u
m11 z      d      w3     vss n w=19u  l=2.3636u ad=76p      pd=27u      as=47.5p    ps=24u
m12 w4     d      z      vss n w=19u  l=2.3636u ad=47.5p    pd=24u      as=76p      ps=27u
m13 w5     c      w4     vss n w=19u  l=2.3636u ad=47.5p    pd=24u      as=47.5p    ps=24u
m14 w6     b      w5     vss n w=19u  l=2.3636u ad=47.5p    pd=24u      as=47.5p    ps=24u
m15 vss    a      w6     vss n w=19u  l=2.3636u ad=168.5p   pd=57u      as=47.5p    ps=24u
C0  vss    a      0.197f
C1  vdd    c      0.057f
C2  z      b      0.548f
C3  w3     vss    0.004f
C4  w5     vss    0.004f
C5  d      b      0.149f
C6  vdd    a      0.069f
C7  w1     vss    0.004f
C8  w2     z      0.010f
C9  c      a      0.215f
C10 vss    z      0.303f
C11 vss    d      0.027f
C12 w3     a      0.007f
C13 z      vdd    0.693f
C14 w5     a      0.009f
C15 w1     a      0.006f
C16 vdd    d      0.022f
C17 z      c      0.129f
C18 vss    b      0.062f
C19 w4     vss    0.004f
C20 w6     vss    0.004f
C21 vdd    b      0.200f
C22 d      c      0.337f
C23 z      a      0.352f
C24 w2     vss    0.004f
C25 w3     z      0.010f
C26 c      b      0.519f
C27 d      a      0.196f
C28 w1     z      0.010f
C29 b      a      0.464f
C30 w4     a      0.008f
C31 vss    vdd    0.007f
C32 w6     a      0.010f
C33 z      d      0.077f
C34 w2     a      0.007f
C35 vss    c      0.042f
C37 z      vss    0.020f
C39 d      vss    0.036f
C40 c      vss    0.053f
C41 b      vss    0.070f
C42 a      vss    0.057f
.ends
