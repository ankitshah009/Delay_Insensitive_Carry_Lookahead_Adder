magic
tech scmos
timestamp 1180600661
<< checkpaint >>
rect -22 -22 62 122
<< ab >>
rect 0 0 40 100
<< pwell >>
rect -4 -4 44 48
<< nwell >>
rect -4 48 44 104
<< polysilicon >>
rect 13 94 15 98
rect 25 94 27 98
rect 13 33 15 55
rect 25 33 27 67
rect 7 32 27 33
rect 7 28 8 32
rect 12 28 27 32
rect 7 27 27 28
rect 13 24 15 27
rect 25 24 27 27
rect 13 2 15 6
rect 25 2 27 6
<< ndiffusion >>
rect 5 12 13 24
rect 5 8 6 12
rect 10 8 13 12
rect 5 6 13 8
rect 15 22 25 24
rect 15 18 18 22
rect 22 18 25 22
rect 15 6 25 18
rect 27 22 35 24
rect 27 18 30 22
rect 34 18 35 22
rect 27 12 35 18
rect 27 8 30 12
rect 34 8 35 12
rect 27 6 35 8
<< pdiffusion >>
rect 5 92 13 94
rect 5 88 6 92
rect 10 88 13 92
rect 5 55 13 88
rect 15 82 25 94
rect 15 78 18 82
rect 22 78 25 82
rect 15 72 25 78
rect 15 68 18 72
rect 22 68 25 72
rect 15 67 25 68
rect 27 92 35 94
rect 27 88 30 92
rect 34 88 35 92
rect 27 82 35 88
rect 27 78 30 82
rect 34 78 35 82
rect 27 72 35 78
rect 27 68 30 72
rect 34 68 35 72
rect 27 67 35 68
rect 15 62 23 67
rect 15 58 18 62
rect 22 58 23 62
rect 15 55 23 58
<< metal1 >>
rect -2 92 42 100
rect -2 88 6 92
rect 10 88 30 92
rect 34 88 42 92
rect 8 32 12 83
rect 8 17 12 28
rect 18 82 22 83
rect 18 72 22 78
rect 18 62 22 68
rect 30 82 34 88
rect 30 72 34 78
rect 30 67 34 68
rect 18 22 22 58
rect 18 17 22 18
rect 30 22 34 23
rect 30 12 34 18
rect -2 8 6 12
rect 10 8 30 12
rect 34 8 42 12
rect -2 0 42 8
<< ntransistor >>
rect 13 6 15 24
rect 25 6 27 24
<< ptransistor >>
rect 13 55 15 94
rect 25 67 27 94
<< polycontact >>
rect 8 28 12 32
<< ndcontact >>
rect 6 8 10 12
rect 18 18 22 22
rect 30 18 34 22
rect 30 8 34 12
<< pdcontact >>
rect 6 88 10 92
rect 18 78 22 82
rect 18 68 22 72
rect 30 88 34 92
rect 30 78 34 82
rect 30 68 34 72
rect 18 58 22 62
<< labels >>
rlabel metal1 10 50 10 50 6 i
rlabel metal1 20 6 20 6 6 vss
rlabel metal1 20 50 20 50 6 nq
rlabel metal1 20 94 20 94 6 vdd
<< end >>
