.subckt cgi2bv0x3 a b c vdd vss z
*   SPICE3 file   created from cgi2bv0x3.ext -      technology: scmos
m00 vdd    b      bn     vdd p w=8u   l=2.3636u ad=37.2658p pd=11.2405u as=34.5p    ps=12.75u
m01 bn     b      vdd    vdd p w=28u  l=2.3636u ad=120.75p  pd=44.625u  as=130.43p  ps=39.3418u
m02 vdd    b      bn     vdd p w=28u  l=2.3636u ad=130.43p  pd=39.3418u as=120.75p  ps=44.625u
m03 n1     bn     vdd    vdd p w=28u  l=2.3636u ad=118p     pd=39.7778u as=130.43p  ps=39.3418u
m04 vdd    bn     n1     vdd p w=28u  l=2.3636u ad=130.43p  pd=39.3418u as=118p     ps=39.7778u
m05 n1     bn     vdd    vdd p w=28u  l=2.3636u ad=118p     pd=39.7778u as=130.43p  ps=39.3418u
m06 z      c      n1     vdd p w=28u  l=2.3636u ad=112p     pd=36u      as=118p     ps=39.7778u
m07 n1     c      z      vdd p w=28u  l=2.3636u ad=118p     pd=39.7778u as=112p     ps=36u
m08 z      c      n1     vdd p w=28u  l=2.3636u ad=112p     pd=36u      as=118p     ps=39.7778u
m09 w1     bn     z      vdd p w=28u  l=2.3636u ad=70p      pd=33u      as=112p     ps=36u
m10 vdd    a      w1     vdd p w=28u  l=2.3636u ad=130.43p  pd=39.3418u as=70p      ps=33u
m11 w2     a      vdd    vdd p w=28u  l=2.3636u ad=70p      pd=33u      as=130.43p  ps=39.3418u
m12 z      bn     w2     vdd p w=28u  l=2.3636u ad=112p     pd=36u      as=70p      ps=33u
m13 w3     bn     z      vdd p w=28u  l=2.3636u ad=70p      pd=33u      as=112p     ps=36u
m14 vdd    a      w3     vdd p w=28u  l=2.3636u ad=130.43p  pd=39.3418u as=70p      ps=33u
m15 n1     a      vdd    vdd p w=28u  l=2.3636u ad=118p     pd=39.7778u as=130.43p  ps=39.3418u
m16 vdd    a      n1     vdd p w=28u  l=2.3636u ad=130.43p  pd=39.3418u as=118p     ps=39.7778u
m17 n1     a      vdd    vdd p w=28u  l=2.3636u ad=118p     pd=39.7778u as=130.43p  ps=39.3418u
m18 bn     b      vss    vss n w=16u  l=2.3636u ad=64p      pd=24u      as=95.6923p ps=33.2308u
m19 vss    b      bn     vss n w=16u  l=2.3636u ad=95.6923p pd=33.2308u as=64p      ps=24u
m20 n3     bn     vss    vss n w=14u  l=2.3636u ad=56p      pd=21.2258u as=83.7308p ps=29.0769u
m21 vss    bn     n3     vss n w=14u  l=2.3636u ad=83.7308p pd=29.0769u as=56p      ps=21.2258u
m22 n3     bn     vss    vss n w=14u  l=2.3636u ad=56p      pd=21.2258u as=83.7308p ps=29.0769u
m23 z      c      n3     vss n w=14u  l=2.3636u ad=56p      pd=22u      as=56p      ps=21.2258u
m24 n3     c      z      vss n w=14u  l=2.3636u ad=56p      pd=21.2258u as=56p      ps=22u
m25 z      c      n3     vss n w=14u  l=2.3636u ad=56p      pd=22u      as=56p      ps=21.2258u
m26 w4     bn     z      vss n w=14u  l=2.3636u ad=35p      pd=19u      as=56p      ps=22u
m27 vss    a      w4     vss n w=14u  l=2.3636u ad=83.7308p pd=29.0769u as=35p      ps=19u
m28 w5     a      vss    vss n w=14u  l=2.3636u ad=35p      pd=19u      as=83.7308p ps=29.0769u
m29 z      bn     w5     vss n w=14u  l=2.3636u ad=56p      pd=22u      as=35p      ps=19u
m30 w6     bn     z      vss n w=14u  l=2.3636u ad=35p      pd=19u      as=56p      ps=22u
m31 vss    a      w6     vss n w=14u  l=2.3636u ad=83.7308p pd=29.0769u as=35p      ps=19u
m32 n3     a      vss    vss n w=20u  l=2.3636u ad=80p      pd=30.3226u as=119.615p ps=41.5385u
m33 vss    a      n3     vss n w=20u  l=2.3636u ad=119.615p pd=41.5385u as=80p      ps=30.3226u
C0  z      bn     0.233f
C1  n1     c      0.073f
C2  w2     vdd    0.005f
C3  n3     z      0.755f
C4  z      vdd    0.291f
C5  a      bn     0.567f
C6  vss    n1     0.050f
C7  n3     a      0.088f
C8  w5     bn     0.008f
C9  w3     z      0.010f
C10 a      vdd    0.094f
C11 c      b      0.008f
C12 w5     n3     0.010f
C13 vss    c      0.024f
C14 n3     bn     0.343f
C15 w3     a      0.007f
C16 w1     z      0.010f
C17 w2     n1     0.010f
C18 bn     vdd    0.250f
C19 n3     vdd    0.033f
C20 vss    b      0.102f
C21 z      n1     0.851f
C22 w6     z      0.010f
C23 z      c      0.186f
C24 n1     a      0.128f
C25 w3     vdd    0.005f
C26 n1     bn     0.109f
C27 w1     vdd    0.005f
C28 a      c      0.064f
C29 n3     n1     0.124f
C30 vss    z      0.217f
C31 n1     vdd    1.036f
C32 c      bn     0.266f
C33 w6     n3     0.010f
C34 vss    a      0.057f
C35 n3     c      0.071f
C36 w4     bn     0.008f
C37 w2     z      0.010f
C38 w3     n1     0.010f
C39 c      vdd    0.025f
C40 bn     b      0.337f
C41 w4     n3     0.010f
C42 n3     b      0.004f
C43 vss    bn     0.354f
C44 w2     a      0.007f
C45 w1     n1     0.010f
C46 b      vdd    0.041f
C47 n3     vss    0.867f
C48 vss    vdd    0.026f
C49 z      a      0.546f
C51 z      vss    0.006f
C52 a      vss    0.085f
C53 c      vss    0.044f
C54 bn     vss    0.121f
C55 b      vss    0.047f
.ends
