magic
tech scmos
timestamp 1183911755
<< checkpaint >>
rect -22 -22 166 94
<< ab >>
rect 0 0 144 72
<< pwell >>
rect -4 -4 148 32
<< nwell >>
rect -4 32 148 76
<< polysilicon >>
rect 9 66 11 70
rect 55 68 111 70
rect 55 60 57 68
rect 65 60 67 64
rect 75 60 77 64
rect 82 60 84 68
rect 92 60 94 64
rect 99 60 101 64
rect 19 52 21 57
rect 38 54 40 59
rect 45 54 47 59
rect 9 34 11 38
rect 19 35 21 38
rect 19 34 34 35
rect 9 33 15 34
rect 19 33 29 34
rect 9 29 10 33
rect 14 29 15 33
rect 9 28 15 29
rect 27 30 29 33
rect 33 30 34 34
rect 27 29 34 30
rect 9 24 11 28
rect 27 26 29 29
rect 38 19 40 48
rect 45 44 47 48
rect 45 43 51 44
rect 45 39 46 43
rect 50 39 51 43
rect 45 38 51 39
rect 55 34 57 48
rect 45 32 57 34
rect 45 19 47 32
rect 65 29 67 48
rect 75 44 77 54
rect 71 43 77 44
rect 71 39 72 43
rect 76 39 77 43
rect 71 38 77 39
rect 65 28 71 29
rect 51 27 57 28
rect 51 23 52 27
rect 56 23 57 27
rect 51 22 57 23
rect 55 19 57 22
rect 65 24 66 28
rect 70 24 71 28
rect 65 23 71 24
rect 65 19 67 23
rect 75 19 77 38
rect 82 34 84 54
rect 109 58 111 68
rect 129 59 131 64
rect 92 44 94 47
rect 88 43 94 44
rect 88 39 89 43
rect 93 39 94 43
rect 88 38 94 39
rect 99 35 101 47
rect 109 44 111 47
rect 129 45 131 49
rect 122 44 131 45
rect 109 42 117 44
rect 115 35 117 42
rect 122 40 123 44
rect 127 40 131 44
rect 122 39 131 40
rect 99 34 105 35
rect 82 32 94 34
rect 82 27 88 28
rect 82 23 83 27
rect 87 23 88 27
rect 82 22 88 23
rect 82 19 84 22
rect 92 19 94 32
rect 99 30 100 34
rect 104 30 105 34
rect 99 29 105 30
rect 115 34 121 35
rect 115 30 116 34
rect 120 30 121 34
rect 115 29 121 30
rect 99 19 101 29
rect 119 26 121 29
rect 129 26 131 39
rect 27 14 29 19
rect 119 15 121 20
rect 129 14 131 19
rect 9 7 11 10
rect 38 7 40 13
rect 45 8 47 13
rect 9 5 40 7
rect 55 4 57 13
rect 65 8 67 13
rect 75 8 77 13
rect 82 4 84 13
rect 92 8 94 13
rect 99 8 101 13
rect 55 2 84 4
<< ndiffusion >>
rect 20 25 27 26
rect 2 23 9 24
rect 2 19 3 23
rect 7 19 9 23
rect 2 18 9 19
rect 4 10 9 18
rect 11 16 16 24
rect 20 21 21 25
rect 25 21 27 25
rect 20 20 27 21
rect 22 19 27 20
rect 29 19 36 26
rect 112 25 119 26
rect 112 21 113 25
rect 117 21 119 25
rect 112 20 119 21
rect 121 25 129 26
rect 121 21 123 25
rect 127 21 129 25
rect 121 20 129 21
rect 11 15 18 16
rect 11 11 13 15
rect 17 11 18 15
rect 31 18 38 19
rect 31 14 32 18
rect 36 14 38 18
rect 31 13 38 14
rect 40 13 45 19
rect 47 18 55 19
rect 47 14 49 18
rect 53 14 55 18
rect 47 13 55 14
rect 57 18 65 19
rect 57 14 59 18
rect 63 14 65 18
rect 57 13 65 14
rect 67 18 75 19
rect 67 14 69 18
rect 73 14 75 18
rect 67 13 75 14
rect 77 13 82 19
rect 84 18 92 19
rect 84 14 86 18
rect 90 14 92 18
rect 84 13 92 14
rect 94 13 99 19
rect 101 18 108 19
rect 101 14 103 18
rect 107 14 108 18
rect 123 19 129 20
rect 131 25 138 26
rect 131 21 133 25
rect 137 21 138 25
rect 131 19 138 21
rect 101 13 108 14
rect 11 10 18 11
<< pdiffusion >>
rect 4 52 9 66
rect 2 50 9 52
rect 2 46 3 50
rect 7 46 9 50
rect 2 43 9 46
rect 2 39 3 43
rect 7 39 9 43
rect 2 38 9 39
rect 11 65 18 66
rect 11 61 13 65
rect 17 61 18 65
rect 11 60 18 61
rect 11 52 17 60
rect 50 54 55 60
rect 30 53 38 54
rect 11 51 19 52
rect 11 47 13 51
rect 17 47 19 51
rect 11 38 19 47
rect 21 44 26 52
rect 30 49 31 53
rect 35 49 38 53
rect 30 48 38 49
rect 40 48 45 54
rect 47 53 55 54
rect 47 49 49 53
rect 53 49 55 53
rect 47 48 55 49
rect 57 53 65 60
rect 57 49 59 53
rect 63 49 65 53
rect 57 48 65 49
rect 67 59 75 60
rect 67 55 69 59
rect 73 55 75 59
rect 67 54 75 55
rect 77 54 82 60
rect 84 59 92 60
rect 84 55 86 59
rect 90 55 92 59
rect 84 54 92 55
rect 67 48 73 54
rect 21 43 28 44
rect 21 39 23 43
rect 27 39 28 43
rect 21 38 28 39
rect 87 47 92 54
rect 94 47 99 60
rect 101 58 106 60
rect 122 58 129 59
rect 101 57 109 58
rect 101 53 103 57
rect 107 53 109 57
rect 101 47 109 53
rect 111 53 116 58
rect 122 54 123 58
rect 127 54 129 58
rect 111 52 118 53
rect 111 48 113 52
rect 117 48 118 52
rect 122 49 129 54
rect 131 55 136 59
rect 131 54 138 55
rect 131 50 133 54
rect 137 50 138 54
rect 131 49 138 50
rect 111 47 118 48
<< metal1 >>
rect -2 68 146 72
rect -2 65 27 68
rect -2 64 13 65
rect 17 64 27 65
rect 31 64 37 68
rect 41 64 118 68
rect 122 64 146 68
rect 13 51 17 61
rect 2 50 7 51
rect 2 46 3 50
rect 31 53 35 64
rect 69 59 73 64
rect 69 54 73 55
rect 81 55 86 59
rect 90 55 91 59
rect 102 57 108 64
rect 59 53 63 54
rect 31 48 35 49
rect 38 49 49 53
rect 53 49 54 53
rect 13 46 17 47
rect 2 43 7 46
rect 2 39 3 43
rect 7 39 15 42
rect 2 38 15 39
rect 21 39 23 43
rect 27 39 28 43
rect 2 24 6 38
rect 21 33 25 39
rect 38 34 42 49
rect 59 43 63 49
rect 45 39 46 43
rect 9 29 10 33
rect 14 29 25 33
rect 28 30 29 34
rect 33 30 44 34
rect 21 25 25 29
rect 2 23 7 24
rect 2 19 3 23
rect 21 20 25 21
rect 2 18 7 19
rect 32 18 36 19
rect 13 15 17 16
rect 13 8 17 11
rect 40 18 44 30
rect 50 28 54 43
rect 59 39 72 43
rect 76 39 77 43
rect 50 27 56 28
rect 50 23 52 27
rect 50 22 56 23
rect 59 18 63 39
rect 81 36 85 55
rect 102 53 103 57
rect 107 53 108 57
rect 122 58 128 64
rect 122 54 123 58
rect 127 54 128 58
rect 133 54 137 55
rect 113 52 117 53
rect 76 32 85 36
rect 89 48 113 50
rect 89 46 117 48
rect 89 43 93 46
rect 121 44 127 50
rect 121 42 123 44
rect 76 29 80 32
rect 66 28 80 29
rect 89 28 93 39
rect 97 34 103 42
rect 113 40 123 42
rect 113 38 127 40
rect 133 34 137 50
rect 97 30 100 34
rect 104 30 111 34
rect 115 30 116 34
rect 120 30 137 34
rect 70 24 80 28
rect 66 23 80 24
rect 40 14 49 18
rect 53 14 54 18
rect 32 8 36 14
rect 59 13 63 14
rect 69 18 73 19
rect 76 18 80 23
rect 83 27 93 28
rect 87 26 93 27
rect 87 25 118 26
rect 87 23 113 25
rect 83 22 113 23
rect 112 21 113 22
rect 117 21 118 25
rect 123 25 127 26
rect 76 14 86 18
rect 90 14 91 18
rect 102 14 103 18
rect 107 14 108 18
rect 69 8 73 14
rect 102 8 108 14
rect 123 8 127 21
rect 133 25 137 30
rect 133 20 137 21
rect -2 4 119 8
rect 123 4 130 8
rect 134 4 146 8
rect -2 0 146 4
<< ntransistor >>
rect 9 10 11 24
rect 27 19 29 26
rect 119 20 121 26
rect 38 13 40 19
rect 45 13 47 19
rect 55 13 57 19
rect 65 13 67 19
rect 75 13 77 19
rect 82 13 84 19
rect 92 13 94 19
rect 99 13 101 19
rect 129 19 131 26
<< ptransistor >>
rect 9 38 11 66
rect 19 38 21 52
rect 38 48 40 54
rect 45 48 47 54
rect 55 48 57 60
rect 65 48 67 60
rect 75 54 77 60
rect 82 54 84 60
rect 92 47 94 60
rect 99 47 101 60
rect 109 47 111 58
rect 129 49 131 59
<< polycontact >>
rect 10 29 14 33
rect 29 30 33 34
rect 46 39 50 43
rect 72 39 76 43
rect 52 23 56 27
rect 66 24 70 28
rect 89 39 93 43
rect 123 40 127 44
rect 83 23 87 27
rect 100 30 104 34
rect 116 30 120 34
<< ndcontact >>
rect 3 19 7 23
rect 21 21 25 25
rect 113 21 117 25
rect 123 21 127 25
rect 13 11 17 15
rect 32 14 36 18
rect 49 14 53 18
rect 59 14 63 18
rect 69 14 73 18
rect 86 14 90 18
rect 103 14 107 18
rect 133 21 137 25
<< pdcontact >>
rect 3 46 7 50
rect 3 39 7 43
rect 13 61 17 65
rect 13 47 17 51
rect 31 49 35 53
rect 49 49 53 53
rect 59 49 63 53
rect 69 55 73 59
rect 86 55 90 59
rect 23 39 27 43
rect 103 53 107 57
rect 123 54 127 58
rect 113 48 117 52
rect 133 50 137 54
<< psubstratepcontact >>
rect 119 4 123 8
rect 130 4 134 8
<< nsubstratencontact >>
rect 27 64 31 68
rect 37 64 41 68
rect 118 64 122 68
<< psubstratepdiff >>
rect 112 8 141 9
rect 112 4 119 8
rect 123 4 130 8
rect 134 4 141 8
rect 112 3 141 4
<< nsubstratendiff >>
rect 22 68 46 69
rect 22 64 27 68
rect 31 64 37 68
rect 41 64 46 68
rect 22 63 46 64
rect 117 68 123 69
rect 117 64 118 68
rect 122 64 123 68
rect 117 63 123 64
<< labels >>
rlabel polycontact 12 31 12 31 6 zn
rlabel polycontact 30 32 30 32 6 n4
rlabel polycontact 54 25 54 25 6 ci
rlabel polycontact 48 41 48 41 6 ci
rlabel polycontact 68 26 68 26 6 n1
rlabel polycontact 85 25 85 25 6 ci
rlabel polycontact 91 41 91 41 6 ci
rlabel polycontact 74 41 74 41 6 n2
rlabel polycontact 118 32 118 32 6 cn
rlabel metal1 17 31 17 31 6 zn
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 40 12 40 6 z
rlabel metal1 23 31 23 31 6 zn
rlabel metal1 47 16 47 16 6 n4
rlabel polycontact 53 25 53 25 6 ci
rlabel metal1 36 32 36 32 6 n4
rlabel polycontact 49 41 49 41 6 ci
rlabel metal1 46 51 46 51 6 n4
rlabel metal1 72 4 72 4 6 vss
rlabel metal1 73 26 73 26 6 n1
rlabel metal1 68 41 68 41 6 n2
rlabel metal1 61 33 61 33 6 n2
rlabel metal1 72 68 72 68 6 vdd
rlabel metal1 83 16 83 16 6 n1
rlabel metal1 108 32 108 32 6 d
rlabel metal1 100 36 100 36 6 d
rlabel metal1 91 36 91 36 6 ci
rlabel metal1 86 57 86 57 6 n1
rlabel metal1 100 24 100 24 6 ci
rlabel metal1 126 32 126 32 6 cn
rlabel metal1 116 40 116 40 6 cp
rlabel metal1 124 44 124 44 6 cp
rlabel metal1 135 37 135 37 6 cn
rlabel pdcontact 115 49 115 49 6 ci
<< end >>
