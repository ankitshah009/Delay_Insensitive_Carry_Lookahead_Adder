magic
tech scmos
timestamp 1179387261
<< checkpaint >>
rect -22 -22 78 94
<< ab >>
rect 0 0 56 72
<< pwell >>
rect -4 -4 60 32
<< nwell >>
rect -4 32 60 76
<< polysilicon >>
rect 9 60 11 65
rect 22 55 24 60
rect 29 55 31 60
rect 36 55 38 60
rect 9 31 11 48
rect 22 42 24 45
rect 17 41 24 42
rect 17 37 18 41
rect 22 37 24 41
rect 17 36 24 37
rect 9 30 15 31
rect 9 26 10 30
rect 14 26 15 30
rect 9 25 15 26
rect 9 21 11 25
rect 19 21 21 36
rect 29 35 31 45
rect 36 42 38 45
rect 36 40 43 42
rect 29 34 35 35
rect 29 30 30 34
rect 34 30 35 34
rect 29 29 35 30
rect 29 21 31 29
rect 41 27 43 40
rect 41 26 47 27
rect 41 22 42 26
rect 46 22 47 26
rect 41 21 47 22
rect 41 18 43 21
rect 9 10 11 15
rect 19 11 21 15
rect 29 11 31 15
rect 41 7 43 12
<< ndiffusion >>
rect 2 20 9 21
rect 2 16 3 20
rect 7 16 9 20
rect 2 15 9 16
rect 11 20 19 21
rect 11 16 13 20
rect 17 16 19 20
rect 11 15 19 16
rect 21 20 29 21
rect 21 16 23 20
rect 27 16 29 20
rect 21 15 29 16
rect 31 18 39 21
rect 31 15 41 18
rect 33 12 41 15
rect 43 17 50 18
rect 43 13 45 17
rect 49 13 50 17
rect 43 12 50 13
rect 33 8 39 12
rect 33 4 34 8
rect 38 4 39 8
rect 33 3 39 4
<< pdiffusion >>
rect 13 68 20 69
rect 13 64 14 68
rect 18 64 20 68
rect 13 60 20 64
rect 2 59 9 60
rect 2 55 3 59
rect 7 55 9 59
rect 2 54 9 55
rect 4 48 9 54
rect 11 55 20 60
rect 11 48 22 55
rect 13 45 22 48
rect 24 45 29 55
rect 31 45 36 55
rect 38 51 43 55
rect 38 50 45 51
rect 38 46 40 50
rect 44 46 45 50
rect 38 45 45 46
<< metal1 >>
rect -2 68 58 72
rect -2 64 14 68
rect 18 64 25 68
rect 29 64 44 68
rect 48 64 58 68
rect 2 55 3 59
rect 7 55 15 59
rect 2 54 15 55
rect 2 21 6 54
rect 10 46 40 50
rect 44 46 45 50
rect 10 30 14 46
rect 17 41 31 42
rect 17 37 18 41
rect 22 38 31 41
rect 22 37 23 38
rect 17 30 23 37
rect 41 34 47 42
rect 29 30 30 34
rect 34 30 47 34
rect 14 26 27 27
rect 10 23 27 26
rect 2 20 7 21
rect 23 20 27 23
rect 33 22 42 26
rect 46 22 47 26
rect 2 16 3 20
rect 2 15 7 16
rect 12 16 13 20
rect 17 16 18 20
rect 2 13 6 15
rect 12 8 18 16
rect 27 16 45 17
rect 23 13 45 16
rect 49 13 50 17
rect -2 4 14 8
rect 18 4 24 8
rect 28 4 34 8
rect 38 4 58 8
rect -2 0 58 4
<< ntransistor >>
rect 9 15 11 21
rect 19 15 21 21
rect 29 15 31 21
rect 41 12 43 18
<< ptransistor >>
rect 9 48 11 60
rect 22 45 24 55
rect 29 45 31 55
rect 36 45 38 55
<< polycontact >>
rect 18 37 22 41
rect 10 26 14 30
rect 30 30 34 34
rect 42 22 46 26
<< ndcontact >>
rect 3 16 7 20
rect 13 16 17 20
rect 23 16 27 20
rect 45 13 49 17
rect 34 4 38 8
<< pdcontact >>
rect 14 64 18 68
rect 3 55 7 59
rect 40 46 44 50
<< psubstratepcontact >>
rect 14 4 18 8
rect 24 4 28 8
<< nsubstratencontact >>
rect 25 64 29 68
rect 44 64 48 68
<< psubstratepdiff >>
rect 13 8 29 9
rect 13 4 14 8
rect 18 4 24 8
rect 28 4 29 8
rect 13 3 29 4
<< nsubstratendiff >>
rect 24 68 49 69
rect 24 64 25 68
rect 29 64 44 68
rect 48 64 49 68
rect 24 63 49 64
<< labels >>
rlabel polycontact 12 28 12 28 6 zn
rlabel metal1 4 36 4 36 6 z
rlabel metal1 25 20 25 20 6 zn
rlabel metal1 20 36 20 36 6 a
rlabel metal1 12 36 12 36 6 zn
rlabel metal1 12 56 12 56 6 z
rlabel metal1 28 4 28 4 6 vss
rlabel metal1 36 24 36 24 6 c
rlabel metal1 36 32 36 32 6 b
rlabel metal1 28 40 28 40 6 a
rlabel metal1 28 68 28 68 6 vdd
rlabel metal1 36 15 36 15 6 zn
rlabel polycontact 44 24 44 24 6 c
rlabel metal1 44 36 44 36 6 b
rlabel metal1 27 48 27 48 6 zn
<< end >>
