magic
tech scmos
timestamp 1179387075
<< checkpaint >>
rect -22 -25 78 105
<< ab >>
rect 0 0 56 80
<< pwell >>
rect -4 -7 60 36
<< nwell >>
rect -4 36 60 87
<< polysilicon >>
rect 13 68 15 73
rect 21 68 23 73
rect 31 68 33 73
rect 39 68 41 73
rect 13 47 15 52
rect 21 47 23 52
rect 9 46 15 47
rect 9 42 10 46
rect 14 42 15 46
rect 9 41 15 42
rect 20 46 26 47
rect 20 42 21 46
rect 25 42 26 46
rect 20 41 26 42
rect 9 23 11 41
rect 20 30 22 41
rect 31 39 33 52
rect 39 49 41 52
rect 39 48 46 49
rect 39 44 41 48
rect 45 44 46 48
rect 39 43 46 44
rect 30 38 36 39
rect 30 34 31 38
rect 35 34 36 38
rect 30 33 36 34
rect 30 30 32 33
rect 20 18 22 23
rect 30 18 32 23
rect 41 22 43 43
rect 9 11 11 16
rect 41 10 43 15
<< ndiffusion >>
rect 13 29 20 30
rect 13 25 14 29
rect 18 25 20 29
rect 13 23 20 25
rect 22 28 30 30
rect 22 24 24 28
rect 28 24 30 28
rect 22 23 30 24
rect 32 23 39 30
rect 2 21 9 23
rect 2 17 3 21
rect 7 17 9 21
rect 2 16 9 17
rect 11 16 17 23
rect 34 22 39 23
rect 34 15 41 22
rect 43 21 50 22
rect 43 17 45 21
rect 49 17 50 21
rect 43 15 50 17
rect 34 13 39 15
rect 33 12 39 13
rect 33 8 34 12
rect 38 8 39 12
rect 33 7 39 8
<< pdiffusion >>
rect 4 72 11 73
rect 4 68 6 72
rect 10 68 11 72
rect 4 52 13 68
rect 15 52 21 68
rect 23 63 31 68
rect 23 59 25 63
rect 29 59 31 63
rect 23 52 31 59
rect 33 52 39 68
rect 41 67 48 68
rect 41 63 43 67
rect 47 63 48 67
rect 41 52 48 63
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect -2 72 58 78
rect -2 68 6 72
rect 10 68 58 72
rect 43 67 47 68
rect 2 59 25 63
rect 29 59 30 63
rect 2 57 14 59
rect 2 30 6 57
rect 10 46 14 47
rect 18 46 22 55
rect 34 54 38 63
rect 43 62 47 63
rect 34 50 47 54
rect 41 48 47 50
rect 18 42 21 46
rect 25 42 31 46
rect 45 44 47 48
rect 41 42 47 44
rect 10 38 14 42
rect 10 34 23 38
rect 30 34 31 38
rect 35 34 39 38
rect 33 31 39 34
rect 2 29 19 30
rect 2 25 14 29
rect 18 25 19 29
rect 24 28 28 29
rect 33 25 46 31
rect 24 21 28 24
rect 2 17 3 21
rect 7 17 45 21
rect 49 17 50 21
rect -2 8 34 12
rect 38 8 58 12
rect -2 2 58 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
<< ntransistor >>
rect 20 23 22 30
rect 30 23 32 30
rect 9 16 11 23
rect 41 15 43 22
<< ptransistor >>
rect 13 52 15 68
rect 21 52 23 68
rect 31 52 33 68
rect 39 52 41 68
<< polycontact >>
rect 10 42 14 46
rect 21 42 25 46
rect 41 44 45 48
rect 31 34 35 38
<< ndcontact >>
rect 14 25 18 29
rect 24 24 28 28
rect 3 17 7 21
rect 45 17 49 21
rect 34 8 38 12
<< pdcontact >>
rect 6 68 10 72
rect 25 59 29 63
rect 43 63 47 67
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
<< psubstratepdiff >>
rect 0 2 56 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 56 2
rect 0 -3 56 -2
<< nsubstratendiff >>
rect 0 82 56 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 56 82
rect 0 77 56 78
<< labels >>
rlabel metal1 4 44 4 44 6 z
rlabel metal1 12 28 12 28 6 z
rlabel polycontact 12 44 12 44 6 b1
rlabel metal1 12 60 12 60 6 z
rlabel metal1 28 6 28 6 6 vss
rlabel metal1 26 23 26 23 6 n3
rlabel metal1 20 36 20 36 6 b1
rlabel metal1 28 44 28 44 6 b2
rlabel metal1 20 52 20 52 6 b2
rlabel metal1 28 74 28 74 6 vdd
rlabel metal1 44 28 44 28 6 a2
rlabel metal1 36 32 36 32 6 a2
rlabel metal1 44 48 44 48 6 a1
rlabel metal1 36 60 36 60 6 a1
rlabel metal1 26 19 26 19 6 n3
<< end >>
