magic
tech scmos
timestamp 1179385459
<< checkpaint >>
rect -22 -25 126 105
<< ab >>
rect 0 0 104 80
<< pwell >>
rect -4 -7 108 36
<< nwell >>
rect -4 36 108 87
<< polysilicon >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 39 70 41 74
rect 49 70 51 74
rect 59 65 61 70
rect 69 61 71 65
rect 79 61 81 65
rect 89 61 91 65
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 39 39 41 42
rect 9 38 41 39
rect 9 37 36 38
rect 29 34 36 37
rect 40 34 41 38
rect 29 33 41 34
rect 29 30 31 33
rect 39 30 41 33
rect 49 39 51 42
rect 59 39 61 42
rect 49 38 61 39
rect 49 34 53 38
rect 57 34 61 38
rect 49 33 61 34
rect 49 30 51 33
rect 59 30 61 33
rect 69 39 71 42
rect 79 39 81 42
rect 89 39 91 42
rect 69 38 91 39
rect 69 34 82 38
rect 86 34 91 38
rect 69 33 91 34
rect 69 30 71 33
rect 79 30 81 33
rect 29 6 31 10
rect 39 6 41 10
rect 49 6 51 10
rect 59 6 61 10
rect 69 9 71 14
rect 79 9 81 14
<< ndiffusion >>
rect 21 22 29 30
rect 21 18 23 22
rect 27 18 29 22
rect 21 15 29 18
rect 21 11 23 15
rect 27 11 29 15
rect 21 10 29 11
rect 31 29 39 30
rect 31 25 33 29
rect 37 25 39 29
rect 31 22 39 25
rect 31 18 33 22
rect 37 18 39 22
rect 31 10 39 18
rect 41 22 49 30
rect 41 18 43 22
rect 47 18 49 22
rect 41 15 49 18
rect 41 11 43 15
rect 47 11 49 15
rect 41 10 49 11
rect 51 29 59 30
rect 51 25 53 29
rect 57 25 59 29
rect 51 22 59 25
rect 51 18 53 22
rect 57 18 59 22
rect 51 10 59 18
rect 61 28 69 30
rect 61 24 63 28
rect 67 24 69 28
rect 61 20 69 24
rect 61 16 63 20
rect 67 16 69 20
rect 61 14 69 16
rect 71 29 79 30
rect 71 25 73 29
rect 77 25 79 29
rect 71 21 79 25
rect 71 17 73 21
rect 77 17 79 21
rect 71 14 79 17
rect 81 27 88 30
rect 81 23 83 27
rect 87 23 88 27
rect 81 19 88 23
rect 81 15 83 19
rect 87 15 88 19
rect 81 14 88 15
rect 61 10 67 14
<< pdiffusion >>
rect 2 69 9 70
rect 2 65 3 69
rect 7 65 9 69
rect 2 62 9 65
rect 2 58 3 62
rect 7 58 9 62
rect 2 55 9 58
rect 2 51 3 55
rect 7 51 9 55
rect 2 42 9 51
rect 11 54 19 70
rect 11 50 13 54
rect 17 50 19 54
rect 11 47 19 50
rect 11 43 13 47
rect 17 43 19 47
rect 11 42 19 43
rect 21 69 29 70
rect 21 65 23 69
rect 27 65 29 69
rect 21 61 29 65
rect 21 57 23 61
rect 27 57 29 61
rect 21 42 29 57
rect 31 54 39 70
rect 31 50 33 54
rect 37 50 39 54
rect 31 47 39 50
rect 31 43 33 47
rect 37 43 39 47
rect 31 42 39 43
rect 41 69 49 70
rect 41 65 43 69
rect 47 65 49 69
rect 41 61 49 65
rect 41 57 43 61
rect 47 57 49 61
rect 41 42 49 57
rect 51 65 56 70
rect 51 54 59 65
rect 51 50 53 54
rect 57 50 59 54
rect 51 47 59 50
rect 51 43 53 47
rect 57 43 59 47
rect 51 42 59 43
rect 61 61 67 65
rect 61 60 69 61
rect 61 56 63 60
rect 67 56 69 60
rect 61 53 69 56
rect 61 49 63 53
rect 67 49 69 53
rect 61 42 69 49
rect 71 54 79 61
rect 71 50 73 54
rect 77 50 79 54
rect 71 47 79 50
rect 71 43 73 47
rect 77 43 79 47
rect 71 42 79 43
rect 81 60 89 61
rect 81 56 83 60
rect 87 56 89 60
rect 81 53 89 56
rect 81 49 83 53
rect 87 49 89 53
rect 81 42 89 49
rect 91 55 96 61
rect 91 54 98 55
rect 91 50 93 54
rect 97 50 98 54
rect 91 47 98 50
rect 91 43 93 47
rect 97 43 98 47
rect 91 42 98 43
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect -2 69 106 78
rect -2 68 3 69
rect 7 68 23 69
rect 3 62 7 65
rect 3 55 7 58
rect 27 68 43 69
rect 23 61 27 65
rect 23 56 27 57
rect 47 68 106 69
rect 43 61 47 65
rect 43 56 47 57
rect 62 60 68 68
rect 62 56 63 60
rect 67 56 68 60
rect 3 50 7 51
rect 13 54 17 55
rect 13 47 17 50
rect 9 43 13 46
rect 33 54 38 55
rect 37 50 38 54
rect 33 47 38 50
rect 17 43 33 46
rect 37 46 38 47
rect 53 54 57 55
rect 53 47 57 50
rect 62 53 68 56
rect 82 60 88 68
rect 82 56 83 60
rect 87 56 88 60
rect 62 49 63 53
rect 67 49 68 53
rect 73 54 77 55
rect 37 43 53 46
rect 9 42 57 43
rect 73 47 77 50
rect 82 53 88 56
rect 82 49 83 53
rect 87 49 88 53
rect 93 54 97 55
rect 93 47 97 50
rect 77 43 93 46
rect 73 42 97 43
rect 26 30 30 42
rect 73 38 77 42
rect 35 34 36 38
rect 40 34 53 38
rect 57 34 77 38
rect 81 34 82 38
rect 86 34 95 38
rect 26 29 57 30
rect 73 29 77 34
rect 26 26 33 29
rect 37 26 53 29
rect 37 25 38 26
rect 33 22 38 25
rect 53 22 57 25
rect 22 18 23 22
rect 27 18 28 22
rect 22 15 28 18
rect 37 18 38 22
rect 33 17 38 18
rect 42 18 43 22
rect 47 18 48 22
rect 22 12 23 15
rect -2 11 23 12
rect 27 12 28 15
rect 42 15 48 18
rect 53 17 57 18
rect 63 28 67 29
rect 63 20 67 24
rect 42 12 43 15
rect 27 11 43 12
rect 47 12 48 15
rect 73 21 77 25
rect 73 16 77 17
rect 83 27 87 28
rect 90 25 95 34
rect 83 19 87 23
rect 63 12 67 16
rect 83 12 87 15
rect 47 11 106 12
rect -2 2 106 11
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
<< ntransistor >>
rect 29 10 31 30
rect 39 10 41 30
rect 49 10 51 30
rect 59 10 61 30
rect 69 14 71 30
rect 79 14 81 30
<< ptransistor >>
rect 9 42 11 70
rect 19 42 21 70
rect 29 42 31 70
rect 39 42 41 70
rect 49 42 51 70
rect 59 42 61 65
rect 69 42 71 61
rect 79 42 81 61
rect 89 42 91 61
<< polycontact >>
rect 36 34 40 38
rect 53 34 57 38
rect 82 34 86 38
<< ndcontact >>
rect 23 18 27 22
rect 23 11 27 15
rect 33 25 37 29
rect 33 18 37 22
rect 43 18 47 22
rect 43 11 47 15
rect 53 25 57 29
rect 53 18 57 22
rect 63 24 67 28
rect 63 16 67 20
rect 73 25 77 29
rect 73 17 77 21
rect 83 23 87 27
rect 83 15 87 19
<< pdcontact >>
rect 3 65 7 69
rect 3 58 7 62
rect 3 51 7 55
rect 13 50 17 54
rect 13 43 17 47
rect 23 65 27 69
rect 23 57 27 61
rect 33 50 37 54
rect 33 43 37 47
rect 43 65 47 69
rect 43 57 47 61
rect 53 50 57 54
rect 53 43 57 47
rect 63 56 67 60
rect 63 49 67 53
rect 73 50 77 54
rect 73 43 77 47
rect 83 56 87 60
rect 83 49 87 53
rect 93 50 97 54
rect 93 43 97 47
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
rect 90 -2 94 2
rect 98 -2 102 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
rect 90 78 94 82
rect 98 78 102 82
<< psubstratepdiff >>
rect 0 2 104 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 104 2
rect 0 -3 104 -2
<< nsubstratendiff >>
rect 0 82 104 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 104 82
rect 0 77 104 78
<< labels >>
rlabel polysilicon 35 36 35 36 6 an
rlabel polycontact 55 36 55 36 6 an
rlabel metal1 12 44 12 44 6 z
rlabel metal1 36 24 36 24 6 z
rlabel metal1 20 44 20 44 6 z
rlabel metal1 28 40 28 40 6 z
rlabel metal1 36 48 36 48 6 z
rlabel metal1 52 6 52 6 6 vss
rlabel metal1 44 28 44 28 6 z
rlabel metal1 52 28 52 28 6 z
rlabel metal1 44 44 44 44 6 z
rlabel metal1 52 44 52 44 6 z
rlabel metal1 52 74 52 74 6 vdd
rlabel polycontact 56 36 56 36 6 an
rlabel metal1 75 35 75 35 6 an
rlabel metal1 92 32 92 32 6 a
rlabel polycontact 84 36 84 36 6 a
rlabel metal1 95 48 95 48 6 an
<< end >>
