magic
tech scmos
timestamp 1179386719
<< checkpaint >>
rect -22 -25 70 105
<< ab >>
rect 0 0 48 80
<< pwell >>
rect -4 -7 52 36
<< nwell >>
rect -4 36 52 87
<< polysilicon >>
rect 12 63 14 68
rect 19 63 21 68
rect 33 60 35 65
rect 12 42 14 48
rect 9 41 15 42
rect 9 37 10 41
rect 14 37 15 41
rect 9 36 15 37
rect 11 22 13 36
rect 19 31 21 48
rect 33 42 35 48
rect 25 41 35 42
rect 25 37 26 41
rect 30 37 35 41
rect 25 36 35 37
rect 17 30 23 31
rect 33 30 35 36
rect 17 26 18 30
rect 22 26 23 30
rect 17 25 23 26
rect 21 22 23 25
rect 33 19 35 24
rect 11 9 13 14
rect 21 9 23 14
<< ndiffusion >>
rect 25 24 33 30
rect 35 29 42 30
rect 35 25 37 29
rect 41 25 42 29
rect 35 24 42 25
rect 25 22 31 24
rect 3 14 11 22
rect 13 21 21 22
rect 13 17 15 21
rect 19 17 21 21
rect 13 14 21 17
rect 23 20 31 22
rect 23 16 26 20
rect 30 16 31 20
rect 23 14 31 16
rect 3 12 9 14
rect 3 8 4 12
rect 8 8 9 12
rect 3 7 9 8
<< pdiffusion >>
rect 5 62 12 63
rect 5 58 6 62
rect 10 58 12 62
rect 5 57 12 58
rect 7 48 12 57
rect 14 48 19 63
rect 21 62 31 63
rect 21 58 26 62
rect 30 60 31 62
rect 30 58 33 60
rect 21 55 33 58
rect 21 51 27 55
rect 31 51 33 55
rect 21 48 33 51
rect 35 54 40 60
rect 35 53 42 54
rect 35 49 37 53
rect 41 49 42 53
rect 35 48 42 49
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect -2 68 50 78
rect 2 62 14 63
rect 2 58 6 62
rect 10 58 14 62
rect 2 57 14 58
rect 26 62 32 68
rect 30 58 32 62
rect 2 22 6 57
rect 26 55 32 58
rect 18 47 22 55
rect 26 51 27 55
rect 31 51 32 55
rect 37 53 41 54
rect 10 43 22 47
rect 10 41 14 43
rect 26 41 30 47
rect 10 33 14 37
rect 18 37 26 39
rect 18 33 30 37
rect 37 30 41 49
rect 17 26 18 30
rect 22 29 41 30
rect 22 26 37 29
rect 37 24 41 25
rect 2 21 23 22
rect 2 17 15 21
rect 19 17 23 21
rect 26 20 30 21
rect 26 12 30 16
rect -2 8 4 12
rect 8 8 50 12
rect -2 2 50 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
<< ntransistor >>
rect 33 24 35 30
rect 11 14 13 22
rect 21 14 23 22
<< ptransistor >>
rect 12 48 14 63
rect 19 48 21 63
rect 33 48 35 60
<< polycontact >>
rect 10 37 14 41
rect 26 37 30 41
rect 18 26 22 30
<< ndcontact >>
rect 37 25 41 29
rect 15 17 19 21
rect 26 16 30 20
rect 4 8 8 12
<< pdcontact >>
rect 6 58 10 62
rect 26 58 30 62
rect 27 51 31 55
rect 37 49 41 53
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
<< psubstratepdiff >>
rect 0 2 48 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 48 2
rect 0 -3 48 -2
<< nsubstratendiff >>
rect 0 82 48 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 48 82
rect 0 77 48 78
<< labels >>
rlabel polycontact 20 28 20 28 6 an
rlabel metal1 4 40 4 40 6 z
rlabel metal1 20 20 20 20 6 z
rlabel metal1 12 20 12 20 6 z
rlabel metal1 20 36 20 36 6 a
rlabel polycontact 12 40 12 40 6 b
rlabel metal1 20 52 20 52 6 b
rlabel metal1 12 60 12 60 6 z
rlabel metal1 24 6 24 6 6 vss
rlabel polycontact 28 40 28 40 6 a
rlabel metal1 24 74 24 74 6 vdd
rlabel metal1 29 28 29 28 6 an
rlabel metal1 39 39 39 39 6 an
<< end >>
