magic
tech scmos
timestamp 1185094813
<< checkpaint >>
rect -22 -22 42 122
<< ab >>
rect 0 0 20 100
<< pwell >>
rect -4 -4 24 48
<< nwell >>
rect -4 48 24 104
<< metal1 >>
rect -2 96 22 100
rect -2 92 4 96
rect 8 92 12 96
rect 16 92 22 96
rect -2 88 22 92
rect -2 8 22 12
rect -2 4 4 8
rect 8 4 12 8
rect 16 4 22 8
rect -2 0 22 4
<< psubstratepcontact >>
rect 4 4 8 8
rect 12 4 16 8
<< nsubstratencontact >>
rect 4 92 8 96
rect 12 92 16 96
<< psubstratepdiff >>
rect 3 8 17 39
rect 3 4 4 8
rect 8 4 12 8
rect 16 4 17 8
rect 3 3 17 4
<< nsubstratendiff >>
rect 3 96 17 97
rect 3 92 4 96
rect 8 92 12 96
rect 16 92 17 96
rect 3 55 17 92
<< labels >>
rlabel metal1 10 6 10 6 6 vss
rlabel metal1 10 94 10 94 6 vdd
<< end >>
