magic
tech scmos
timestamp 1179387569
<< checkpaint >>
rect -22 -25 94 105
<< ab >>
rect 0 0 72 80
<< pwell >>
rect -4 -7 76 36
<< nwell >>
rect -4 36 76 87
<< polysilicon >>
rect 32 66 34 71
rect 42 66 44 71
rect 49 66 51 71
rect 13 62 15 66
rect 21 62 23 66
rect 13 40 15 46
rect 21 43 23 46
rect 9 39 15 40
rect 9 35 10 39
rect 14 35 15 39
rect 9 34 15 35
rect 19 42 25 43
rect 61 61 63 65
rect 61 42 63 45
rect 19 38 20 42
rect 24 38 25 42
rect 19 37 25 38
rect 32 37 34 42
rect 42 39 44 42
rect 9 30 11 34
rect 19 30 21 37
rect 29 35 34 37
rect 39 38 45 39
rect 29 30 31 35
rect 39 34 40 38
rect 44 34 45 38
rect 39 33 45 34
rect 43 28 45 33
rect 49 34 51 42
rect 61 41 70 42
rect 61 40 65 41
rect 64 37 65 40
rect 69 37 70 41
rect 64 36 70 37
rect 49 32 57 34
rect 55 31 57 32
rect 55 30 63 31
rect 43 25 47 28
rect 19 18 21 23
rect 9 11 11 16
rect 29 8 31 23
rect 45 22 47 25
rect 55 26 58 30
rect 62 26 63 30
rect 55 25 63 26
rect 55 22 57 25
rect 45 12 47 16
rect 55 12 57 16
rect 68 8 70 36
rect 29 6 70 8
<< ndiffusion >>
rect 4 22 9 30
rect 2 21 9 22
rect 2 17 3 21
rect 7 17 9 21
rect 2 16 9 17
rect 11 28 19 30
rect 11 24 13 28
rect 17 24 19 28
rect 11 23 19 24
rect 21 29 29 30
rect 21 25 23 29
rect 27 25 29 29
rect 21 23 29 25
rect 31 23 41 30
rect 11 16 16 23
rect 33 22 41 23
rect 33 16 45 22
rect 47 21 55 22
rect 47 17 49 21
rect 53 17 55 21
rect 47 16 55 17
rect 57 21 64 22
rect 57 17 59 21
rect 63 17 64 21
rect 57 16 64 17
rect 33 15 43 16
rect 33 11 38 15
rect 42 11 43 15
rect 33 10 43 11
<< pdiffusion >>
rect 4 72 11 73
rect 4 68 6 72
rect 10 68 11 72
rect 53 72 59 73
rect 4 62 11 68
rect 53 68 54 72
rect 58 68 59 72
rect 53 66 59 68
rect 25 62 32 66
rect 4 46 13 62
rect 15 46 21 62
rect 23 61 32 62
rect 23 57 25 61
rect 29 57 32 61
rect 23 46 32 57
rect 27 42 32 46
rect 34 47 42 66
rect 34 43 36 47
rect 40 43 42 47
rect 34 42 42 43
rect 44 42 49 66
rect 51 61 59 66
rect 51 45 61 61
rect 63 60 70 61
rect 63 56 65 60
rect 69 56 70 60
rect 63 55 70 56
rect 63 45 68 55
rect 51 42 59 45
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect -2 72 74 78
rect -2 68 6 72
rect 10 68 54 72
rect 58 68 74 72
rect 2 61 31 62
rect 2 58 25 61
rect 2 28 6 58
rect 24 57 25 58
rect 29 58 31 61
rect 36 60 69 63
rect 36 59 65 60
rect 29 57 30 58
rect 36 54 40 59
rect 65 55 69 56
rect 10 50 40 54
rect 10 39 14 50
rect 31 43 36 47
rect 40 43 41 47
rect 31 42 35 43
rect 19 38 20 42
rect 24 38 35 42
rect 50 39 54 55
rect 58 47 62 55
rect 58 43 70 47
rect 65 41 70 43
rect 10 31 27 35
rect 23 29 27 31
rect 2 24 13 28
rect 17 24 18 28
rect 23 24 27 25
rect 31 24 35 38
rect 40 38 54 39
rect 44 34 54 38
rect 40 33 54 34
rect 58 31 62 39
rect 69 37 70 41
rect 65 36 70 37
rect 66 35 70 36
rect 58 30 70 31
rect 62 26 70 30
rect 58 25 70 26
rect 31 21 54 24
rect 2 17 3 21
rect 7 20 49 21
rect 7 17 35 20
rect 48 17 49 20
rect 53 17 54 21
rect 58 17 59 21
rect 63 17 64 21
rect 38 15 42 16
rect -2 11 38 12
rect 58 12 64 17
rect 42 11 74 12
rect -2 2 74 11
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
<< ntransistor >>
rect 9 16 11 30
rect 19 23 21 30
rect 29 23 31 30
rect 45 16 47 22
rect 55 16 57 22
<< ptransistor >>
rect 13 46 15 62
rect 21 46 23 62
rect 32 42 34 66
rect 42 42 44 66
rect 49 42 51 66
rect 61 45 63 61
<< polycontact >>
rect 10 35 14 39
rect 20 38 24 42
rect 40 34 44 38
rect 65 37 69 41
rect 58 26 62 30
<< ndcontact >>
rect 3 17 7 21
rect 13 24 17 28
rect 23 25 27 29
rect 49 17 53 21
rect 59 17 63 21
rect 38 11 42 15
<< pdcontact >>
rect 6 68 10 72
rect 54 68 58 72
rect 25 57 29 61
rect 36 43 40 47
rect 65 56 69 60
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
<< psubstratepdiff >>
rect 0 2 72 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 72 2
rect 0 -3 72 -2
<< nsubstratendiff >>
rect 0 82 72 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 72 82
rect 0 77 72 78
<< labels >>
rlabel ptransistor 22 51 22 51 6 an
rlabel metal1 4 40 4 40 6 z
rlabel metal1 25 29 25 29 6 bn
rlabel metal1 12 42 12 42 6 bn
rlabel metal1 12 60 12 60 6 z
rlabel metal1 20 60 20 60 6 z
rlabel metal1 36 6 36 6 6 vss
rlabel metal1 18 19 18 19 6 an
rlabel metal1 27 40 27 40 6 an
rlabel metal1 36 45 36 45 6 an
rlabel pdcontact 28 60 28 60 6 z
rlabel metal1 36 74 36 74 6 vdd
rlabel ndcontact 51 20 51 20 6 an
rlabel metal1 44 36 44 36 6 a2
rlabel metal1 52 44 52 44 6 a2
rlabel metal1 68 28 68 28 6 a1
rlabel metal1 60 32 60 32 6 a1
rlabel metal1 68 44 68 44 6 b
rlabel metal1 60 52 60 52 6 b
rlabel pdcontact 67 59 67 59 6 bn
<< end >>
