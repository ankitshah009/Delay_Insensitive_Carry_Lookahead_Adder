magic
tech scmos
timestamp 1179386685
<< checkpaint >>
rect -22 -25 78 105
<< ab >>
rect 0 0 56 80
<< pwell >>
rect -4 -7 60 36
<< nwell >>
rect -4 36 60 87
<< polysilicon >>
rect 10 70 12 74
rect 17 70 19 74
rect 27 70 29 74
rect 34 70 36 74
rect 44 66 46 71
rect 10 39 12 42
rect 17 39 19 42
rect 27 39 29 42
rect 34 39 36 42
rect 4 38 13 39
rect 4 34 5 38
rect 9 34 13 38
rect 4 33 13 34
rect 17 38 29 39
rect 17 34 18 38
rect 22 37 29 38
rect 33 38 39 39
rect 22 34 23 37
rect 17 33 23 34
rect 33 34 34 38
rect 38 34 39 38
rect 33 33 39 34
rect 11 30 13 33
rect 21 30 23 33
rect 44 31 46 42
rect 44 30 50 31
rect 44 27 45 30
rect 33 26 45 27
rect 49 26 50 30
rect 33 25 50 26
rect 33 22 35 25
rect 11 10 13 15
rect 21 10 23 15
rect 33 6 35 10
<< ndiffusion >>
rect 2 15 11 30
rect 13 29 21 30
rect 13 25 15 29
rect 19 25 21 29
rect 13 15 21 25
rect 23 22 31 30
rect 23 15 33 22
rect 2 12 9 15
rect 2 8 4 12
rect 8 8 9 12
rect 25 12 33 15
rect 2 7 9 8
rect 25 8 26 12
rect 30 10 33 12
rect 35 21 42 22
rect 35 17 37 21
rect 41 17 42 21
rect 35 16 42 17
rect 35 10 40 16
rect 30 8 31 10
rect 25 7 31 8
<< pdiffusion >>
rect 2 69 10 70
rect 2 65 4 69
rect 8 65 10 69
rect 2 62 10 65
rect 2 58 4 62
rect 8 58 10 62
rect 2 42 10 58
rect 12 42 17 70
rect 19 61 27 70
rect 19 57 21 61
rect 25 57 27 61
rect 19 54 27 57
rect 19 50 21 54
rect 25 50 27 54
rect 19 42 27 50
rect 29 42 34 70
rect 36 66 42 70
rect 36 65 44 66
rect 36 61 38 65
rect 42 61 44 65
rect 36 57 44 61
rect 36 53 38 57
rect 42 53 44 57
rect 36 42 44 53
rect 46 55 51 66
rect 46 54 53 55
rect 46 50 48 54
rect 52 50 53 54
rect 46 47 53 50
rect 46 43 48 47
rect 52 43 53 47
rect 46 42 53 43
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect -2 69 58 78
rect -2 68 4 69
rect 3 65 4 68
rect 8 68 58 69
rect 8 65 9 68
rect 3 62 9 65
rect 38 65 42 68
rect 3 58 4 62
rect 8 58 9 62
rect 21 61 25 62
rect 21 55 25 57
rect 38 57 42 61
rect 17 54 30 55
rect 17 50 21 54
rect 25 50 30 54
rect 38 52 42 53
rect 48 54 52 55
rect 9 42 22 46
rect 5 38 9 39
rect 5 21 9 34
rect 18 38 22 42
rect 18 33 22 34
rect 26 29 30 50
rect 48 47 52 50
rect 48 39 52 43
rect 14 25 15 29
rect 19 25 30 29
rect 34 38 52 39
rect 38 35 52 38
rect 34 21 38 34
rect 42 30 54 31
rect 42 26 45 30
rect 49 26 54 30
rect 42 25 54 26
rect 5 17 37 21
rect 41 17 42 21
rect 50 17 54 25
rect -2 8 4 12
rect 8 8 26 12
rect 30 8 58 12
rect -2 2 58 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
<< ntransistor >>
rect 11 15 13 30
rect 21 15 23 30
rect 33 10 35 22
<< ptransistor >>
rect 10 42 12 70
rect 17 42 19 70
rect 27 42 29 70
rect 34 42 36 70
rect 44 42 46 66
<< polycontact >>
rect 5 34 9 38
rect 18 34 22 38
rect 34 34 38 38
rect 45 26 49 30
<< ndcontact >>
rect 15 25 19 29
rect 4 8 8 12
rect 26 8 30 12
rect 37 17 41 21
<< pdcontact >>
rect 4 65 8 69
rect 4 58 8 62
rect 21 57 25 61
rect 21 50 25 54
rect 38 61 42 65
rect 38 53 42 57
rect 48 50 52 54
rect 48 43 52 47
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
<< psubstratepdiff >>
rect 0 2 56 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 56 2
rect 0 -3 56 -2
<< nsubstratendiff >>
rect 0 82 56 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 56 82
rect 0 77 56 78
<< labels >>
rlabel polycontact 8 36 8 36 6 an
rlabel polycontact 36 36 36 36 6 an
rlabel metal1 7 28 7 28 6 an
rlabel metal1 12 44 12 44 6 b
rlabel metal1 20 52 20 52 6 z
rlabel metal1 28 6 28 6 6 vss
rlabel metal1 36 28 36 28 6 an
rlabel metal1 23 19 23 19 6 an
rlabel metal1 28 40 28 40 6 z
rlabel metal1 28 74 28 74 6 vdd
rlabel metal1 44 28 44 28 6 a
rlabel metal1 52 24 52 24 6 a
rlabel pdcontact 50 45 50 45 6 an
<< end >>
