magic
tech scmos
timestamp 1179385781
<< checkpaint >>
rect -22 -25 86 105
<< ab >>
rect 0 0 64 80
<< pwell >>
rect -4 -7 68 36
<< nwell >>
rect -4 36 68 87
<< polysilicon >>
rect 9 68 11 74
rect 20 72 26 73
rect 20 68 21 72
rect 25 68 26 72
rect 20 67 26 68
rect 9 47 11 50
rect 9 46 18 47
rect 9 45 13 46
rect 12 42 13 45
rect 17 42 18 46
rect 12 30 18 42
rect 22 40 26 67
rect 36 61 38 66
rect 43 61 45 66
rect 36 50 38 53
rect 43 50 45 53
rect 32 49 38 50
rect 32 45 33 49
rect 37 45 38 49
rect 32 44 38 45
rect 42 49 48 50
rect 42 45 43 49
rect 47 45 48 49
rect 42 44 48 45
rect 22 38 37 40
rect 9 28 18 30
rect 23 33 29 34
rect 23 29 24 33
rect 28 29 29 33
rect 23 28 29 29
rect 33 32 37 38
rect 33 28 49 32
rect 9 25 11 28
rect 16 25 18 28
rect 26 25 28 28
rect 33 25 35 28
rect 40 25 42 28
rect 47 25 49 28
rect 26 14 28 19
rect 33 14 35 19
rect 40 14 42 19
rect 47 15 49 19
rect 9 6 11 10
rect 16 6 18 10
<< ndiffusion >>
rect 2 24 9 25
rect 2 20 3 24
rect 7 20 9 24
rect 2 10 9 20
rect 11 10 16 25
rect 18 24 26 25
rect 18 20 20 24
rect 24 20 26 24
rect 18 19 26 20
rect 28 19 33 25
rect 35 19 40 25
rect 42 19 47 25
rect 49 24 56 25
rect 49 20 51 24
rect 55 20 56 24
rect 49 19 56 20
rect 18 10 24 19
<< pdiffusion >>
rect 2 63 9 68
rect 2 59 3 63
rect 7 59 9 63
rect 2 55 9 59
rect 2 51 3 55
rect 7 51 9 55
rect 2 50 9 51
rect 11 67 18 68
rect 11 63 13 67
rect 17 63 18 67
rect 11 50 18 63
rect 28 72 34 73
rect 28 68 29 72
rect 33 68 34 72
rect 28 61 34 68
rect 28 53 36 61
rect 38 53 43 61
rect 45 58 56 61
rect 45 54 51 58
rect 55 54 56 58
rect 45 53 56 54
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect -2 72 66 78
rect -2 68 21 72
rect 25 68 29 72
rect 33 68 66 72
rect 12 67 18 68
rect 12 63 13 67
rect 17 63 18 67
rect 2 59 3 63
rect 7 59 8 63
rect 12 60 18 63
rect 2 56 8 59
rect 22 58 56 63
rect 22 57 51 58
rect 2 55 18 56
rect 2 51 3 55
rect 7 51 18 55
rect 2 50 18 51
rect 2 38 8 50
rect 22 46 28 57
rect 50 54 51 57
rect 55 54 56 58
rect 12 42 13 46
rect 17 42 28 46
rect 33 49 39 50
rect 37 45 39 49
rect 33 38 39 45
rect 2 32 19 38
rect 23 34 39 38
rect 43 49 47 53
rect 23 33 29 34
rect 2 24 8 32
rect 23 29 24 33
rect 28 29 29 33
rect 23 28 29 29
rect 2 20 3 24
rect 7 20 8 24
rect 2 17 8 20
rect 19 20 20 24
rect 24 20 25 24
rect 19 12 25 20
rect 43 12 47 45
rect 50 24 56 54
rect 50 20 51 24
rect 55 20 56 24
rect 50 17 56 20
rect -2 2 66 12
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
<< ntransistor >>
rect 9 10 11 25
rect 16 10 18 25
rect 26 19 28 25
rect 33 19 35 25
rect 40 19 42 25
rect 47 19 49 25
<< ptransistor >>
rect 9 50 11 68
rect 36 53 38 61
rect 43 53 45 61
<< polycontact >>
rect 21 68 25 72
rect 13 42 17 46
rect 33 45 37 49
rect 43 45 47 49
rect 24 29 28 33
<< ndcontact >>
rect 3 20 7 24
rect 20 20 24 24
rect 51 20 55 24
<< pdcontact >>
rect 3 59 7 63
rect 3 51 7 55
rect 13 63 17 67
rect 29 68 33 72
rect 51 54 55 58
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
<< psubstratepdiff >>
rect 0 2 64 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 64 2
rect 0 -3 64 -2
<< nsubstratendiff >>
rect 0 82 64 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 64 82
rect 0 77 64 78
<< labels >>
rlabel polysilicon 15 37 15 37 6 an
rlabel metal1 12 36 12 36 6 z
rlabel metal1 4 40 4 40 6 z
rlabel metal1 12 52 12 52 6 z
rlabel metal1 28 36 28 36 6 a
rlabel metal1 20 44 20 44 6 an
rlabel metal1 32 6 32 6 6 vss
rlabel metal1 36 40 36 40 6 a
rlabel metal1 32 74 32 74 6 vdd
rlabel metal1 53 40 53 40 6 an
<< end >>
