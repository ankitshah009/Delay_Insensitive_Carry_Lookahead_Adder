.subckt an12_x1 i0 i1 q vdd vss
*   SPICE3 file   created from an12_x1.ext -      technology: scmos
m00 w1     i0     q      vdd p w=40u  l=2.3636u ad=120p     pd=46u      as=400p     ps=104u
m01 vdd    w2     w1     vdd p w=40u  l=2.3636u ad=240p     pd=66.6667u as=120p     ps=46u
m02 w2     i1     vdd    vdd p w=20u  l=2.3636u ad=160p     pd=56u      as=120p     ps=33.3333u
m03 q      i0     vss    vss n w=10u  l=2.3636u ad=50p      pd=20u      as=92p      ps=36u
m04 vss    w2     q      vss n w=10u  l=2.3636u ad=92p      pd=36u      as=50p      ps=20u
m05 w2     i1     vss    vss n w=10u  l=2.3636u ad=80p      pd=36u      as=92p      ps=36u
C0  q      vdd    0.077f
C1  i1     i0     0.430f
C2  q      i0     0.435f
C3  vdd    w2     0.023f
C4  w2     i0     0.168f
C5  i1     q      0.159f
C6  vss    i0     0.017f
C7  w1     vdd    0.014f
C8  i1     w2     0.408f
C9  q      w2     0.061f
C10 w1     i0     0.041f
C11 vdd    i0     0.041f
C12 vss    i1     0.067f
C13 vss    q      0.152f
C14 i1     vdd    0.094f
C15 vss    w2     0.051f
C17 i1     vss    0.042f
C18 q      vss    0.028f
C20 w2     vss    0.040f
C21 i0     vss    0.037f
.ends
