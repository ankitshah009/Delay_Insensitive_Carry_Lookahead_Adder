magic
tech scmos
timestamp 1179387105
<< checkpaint >>
rect -22 -22 78 94
<< ab >>
rect 0 0 56 72
<< pwell >>
rect -4 -4 60 32
<< nwell >>
rect -4 32 60 76
<< polysilicon >>
rect 23 66 25 70
rect 30 66 32 70
rect 37 66 39 70
rect 13 57 15 62
rect 13 35 15 46
rect 23 36 25 39
rect 9 34 15 35
rect 9 30 10 34
rect 14 30 15 34
rect 9 29 15 30
rect 19 35 26 36
rect 19 31 21 35
rect 25 31 26 35
rect 19 30 26 31
rect 9 19 11 29
rect 19 19 21 30
rect 30 28 32 39
rect 37 36 39 39
rect 37 35 47 36
rect 37 34 42 35
rect 41 31 42 34
rect 46 31 47 35
rect 41 30 47 31
rect 30 27 37 28
rect 30 23 32 27
rect 36 23 37 27
rect 30 22 37 23
rect 31 19 33 22
rect 41 19 43 30
rect 9 5 11 10
rect 19 5 21 10
rect 31 5 33 10
rect 41 5 43 10
<< ndiffusion >>
rect 2 18 9 19
rect 2 14 3 18
rect 7 14 9 18
rect 2 13 9 14
rect 4 10 9 13
rect 11 17 19 19
rect 11 13 13 17
rect 17 13 19 17
rect 11 10 19 13
rect 21 10 31 19
rect 33 17 41 19
rect 33 13 35 17
rect 39 13 41 17
rect 33 10 41 13
rect 43 15 50 19
rect 43 11 45 15
rect 49 11 50 15
rect 43 10 50 11
rect 23 8 29 10
rect 23 4 24 8
rect 28 4 29 8
rect 23 3 29 4
<< pdiffusion >>
rect 5 58 11 59
rect 5 54 6 58
rect 10 57 11 58
rect 18 57 23 66
rect 10 54 13 57
rect 5 46 13 54
rect 15 51 23 57
rect 15 47 17 51
rect 21 47 23 51
rect 15 46 23 47
rect 18 39 23 46
rect 25 39 30 66
rect 32 39 37 66
rect 39 65 48 66
rect 39 61 42 65
rect 46 61 48 65
rect 39 58 48 61
rect 39 54 42 58
rect 46 54 48 58
rect 39 39 48 54
<< metal1 >>
rect -2 68 58 72
rect -2 64 4 68
rect 8 65 58 68
rect 8 64 42 65
rect 5 58 11 64
rect 41 61 42 64
rect 46 64 58 65
rect 46 61 47 64
rect 5 54 6 58
rect 10 54 11 58
rect 2 47 17 51
rect 21 47 22 51
rect 2 45 14 47
rect 2 19 6 45
rect 26 43 30 59
rect 41 58 47 61
rect 41 54 42 58
rect 46 54 47 58
rect 34 45 47 51
rect 18 37 30 43
rect 20 35 26 37
rect 42 35 47 45
rect 10 34 14 35
rect 20 31 21 35
rect 25 31 26 35
rect 10 26 14 30
rect 34 28 38 35
rect 46 31 47 35
rect 42 30 47 31
rect 32 27 38 28
rect 10 22 23 26
rect 36 26 38 27
rect 36 23 47 26
rect 32 22 47 23
rect 34 21 47 22
rect 2 18 7 19
rect 2 14 3 18
rect 2 13 7 14
rect 12 13 13 17
rect 17 13 35 17
rect 39 13 40 17
rect 45 15 49 16
rect 45 8 49 11
rect -2 4 24 8
rect 28 4 58 8
rect -2 0 58 4
<< ntransistor >>
rect 9 10 11 19
rect 19 10 21 19
rect 31 10 33 19
rect 41 10 43 19
<< ptransistor >>
rect 13 46 15 57
rect 23 39 25 66
rect 30 39 32 66
rect 37 39 39 66
<< polycontact >>
rect 10 30 14 34
rect 21 31 25 35
rect 42 31 46 35
rect 32 23 36 27
<< ndcontact >>
rect 3 14 7 18
rect 13 13 17 17
rect 35 13 39 17
rect 45 11 49 15
rect 24 4 28 8
<< pdcontact >>
rect 6 54 10 58
rect 17 47 21 51
rect 42 61 46 65
rect 42 54 46 58
<< nsubstratencontact >>
rect 4 64 8 68
<< nsubstratendiff >>
rect 3 68 9 69
rect 3 64 4 68
rect 8 64 9 68
rect 3 63 9 64
<< labels >>
rlabel metal1 4 32 4 32 6 z
rlabel polycontact 12 32 12 32 6 b
rlabel metal1 20 24 20 24 6 b
rlabel metal1 20 40 20 40 6 a3
rlabel metal1 12 48 12 48 6 z
rlabel metal1 28 4 28 4 6 vss
rlabel metal1 26 15 26 15 6 n3
rlabel metal1 36 28 36 28 6 a2
rlabel metal1 28 48 28 48 6 a3
rlabel metal1 36 48 36 48 6 a1
rlabel metal1 28 68 28 68 6 vdd
rlabel metal1 44 24 44 24 6 a2
rlabel metal1 44 44 44 44 6 a1
<< end >>
