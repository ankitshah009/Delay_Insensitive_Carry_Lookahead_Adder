magic
tech scmos
timestamp 1179386636
<< checkpaint >>
rect -22 -25 78 105
<< ab >>
rect 0 0 56 80
<< pwell >>
rect -4 -7 60 36
<< nwell >>
rect -4 36 60 87
<< polysilicon >>
rect 9 63 11 68
rect 19 63 21 68
rect 29 63 31 68
rect 39 63 41 68
rect 9 38 11 53
rect 19 48 21 53
rect 16 47 24 48
rect 16 43 17 47
rect 21 43 24 47
rect 16 42 24 43
rect 9 37 15 38
rect 9 33 10 37
rect 14 34 15 37
rect 14 33 17 34
rect 9 32 17 33
rect 15 29 17 32
rect 22 29 24 42
rect 29 47 31 53
rect 29 46 35 47
rect 29 42 30 46
rect 34 42 35 46
rect 29 41 35 42
rect 29 29 31 41
rect 39 38 41 53
rect 39 37 47 38
rect 39 34 42 37
rect 36 33 42 34
rect 46 33 47 37
rect 36 32 47 33
rect 36 29 38 32
rect 15 12 17 17
rect 22 12 24 17
rect 29 12 31 17
rect 36 12 38 17
<< ndiffusion >>
rect 10 23 15 29
rect 8 22 15 23
rect 8 18 9 22
rect 13 18 15 22
rect 8 17 15 18
rect 17 17 22 29
rect 24 17 29 29
rect 31 17 36 29
rect 38 22 49 29
rect 38 18 43 22
rect 47 18 49 22
rect 38 17 49 18
<< pdiffusion >>
rect 2 62 9 63
rect 2 58 3 62
rect 7 58 9 62
rect 2 53 9 58
rect 11 59 19 63
rect 11 55 13 59
rect 17 55 19 59
rect 11 53 19 55
rect 21 62 29 63
rect 21 58 23 62
rect 27 58 29 62
rect 21 53 29 58
rect 31 59 39 63
rect 31 55 33 59
rect 37 55 39 59
rect 31 53 39 55
rect 41 62 49 63
rect 41 58 44 62
rect 48 58 49 62
rect 41 53 49 58
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect -2 68 58 78
rect 2 62 8 68
rect 2 58 3 62
rect 7 58 8 62
rect 22 62 28 68
rect 13 59 17 60
rect 22 58 23 62
rect 27 58 28 62
rect 33 59 38 63
rect 13 54 17 55
rect 37 55 38 59
rect 43 62 49 68
rect 43 58 44 62
rect 48 58 49 62
rect 33 54 38 55
rect 2 50 38 54
rect 2 22 6 50
rect 42 47 46 55
rect 16 43 17 47
rect 21 43 22 47
rect 10 37 14 39
rect 18 38 22 43
rect 25 42 30 46
rect 34 42 46 47
rect 18 33 30 38
rect 34 33 38 42
rect 42 37 46 39
rect 10 29 14 33
rect 10 25 22 29
rect 2 18 9 22
rect 13 18 14 22
rect 2 17 6 18
rect 18 17 22 25
rect 26 17 30 33
rect 42 29 46 33
rect 34 25 46 29
rect 34 17 38 25
rect 42 18 43 22
rect 47 18 48 22
rect 42 12 48 18
rect -2 2 58 12
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
<< ntransistor >>
rect 15 17 17 29
rect 22 17 24 29
rect 29 17 31 29
rect 36 17 38 29
<< ptransistor >>
rect 9 53 11 63
rect 19 53 21 63
rect 29 53 31 63
rect 39 53 41 63
<< polycontact >>
rect 17 43 21 47
rect 10 33 14 37
rect 30 42 34 46
rect 42 33 46 37
<< ndcontact >>
rect 9 18 13 22
rect 43 18 47 22
<< pdcontact >>
rect 3 58 7 62
rect 13 55 17 59
rect 23 58 27 62
rect 33 55 37 59
rect 44 58 48 62
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
<< psubstratepdiff >>
rect 0 2 56 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 56 2
rect 0 -3 56 -2
<< nsubstratendiff >>
rect 0 82 56 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 56 82
rect 0 77 56 78
<< labels >>
rlabel metal1 4 32 4 32 6 z
rlabel metal1 12 32 12 32 6 d
rlabel metal1 12 52 12 52 6 z
rlabel metal1 28 6 28 6 6 vss
rlabel metal1 20 20 20 20 6 d
rlabel metal1 28 24 28 24 6 c
rlabel metal1 20 36 20 36 6 c
rlabel metal1 28 44 28 44 6 b
rlabel metal1 28 52 28 52 6 z
rlabel metal1 20 52 20 52 6 z
rlabel metal1 28 74 28 74 6 vdd
rlabel metal1 36 20 36 20 6 a
rlabel metal1 44 32 44 32 6 a
rlabel metal1 36 36 36 36 6 b
rlabel metal1 44 52 44 52 6 b
rlabel metal1 36 60 36 60 6 z
<< end >>
