.subckt dfnt1v0x2 cp d vdd vss z
*   SPICE3 file   created from dfnt1v0x2.ext -      technology: scmos
m00 vdd    zn     z      vdd p w=28u  l=2.3636u ad=140.56p  pd=61.04u   as=168p     ps=70u
m01 zn     n4     vdd    vdd p w=14u  l=2.3636u ad=82p      pd=42u      as=70.28p   ps=30.52u
m02 w1     zn     vdd    vdd p w=6u   l=2.3636u ad=15p      pd=11u      as=30.12p   ps=13.08u
m03 n4     ci     w1     vdd p w=6u   l=2.3636u ad=26p      pd=13.3333u as=15p      ps=11u
m04 n2     cn     n4     vdd p w=12u  l=2.3636u ad=48p      pd=20u      as=52p      ps=26.6667u
m05 vdd    n1     n2     vdd p w=12u  l=2.3636u ad=60.24p   pd=26.16u   as=48p      ps=20u
m06 w2     n2     vdd    vdd p w=6u   l=2.3636u ad=15p      pd=11u      as=30.12p   ps=13.08u
m07 n1     cn     w2     vdd p w=6u   l=2.3636u ad=26.2105p pd=13.2632u as=15p      ps=11u
m08 vss    zn     z      vss n w=14u  l=2.3636u ad=76.5172p pd=41.0345u as=82p      ps=42u
m09 vss    n4     zn     vss n w=7u   l=2.3636u ad=38.2586p pd=20.5172u as=47p      ps=28u
m10 w3     ci     n1     vdd p w=13u  l=2.3636u ad=32.5p    pd=18u      as=56.7895p ps=28.7368u
m11 vdd    d      w3     vdd p w=13u  l=2.3636u ad=65.26p   pd=28.34u   as=32.5p    ps=18u
m12 ci     cn     vdd    vdd p w=11u  l=2.3636u ad=67p      pd=36u      as=55.22p   ps=23.98u
m13 cn     cp     vdd    vdd p w=10u  l=2.3636u ad=62p      pd=34u      as=50.2p    ps=21.8u
m14 vss    cn     ci     vss n w=6u   l=2.3636u ad=32.7931p pd=17.5862u as=42p      ps=26u
m15 w4     zn     vss    vss n w=6u   l=2.3636u ad=15p      pd=11u      as=32.7931p ps=17.5862u
m16 n4     cn     w4     vss n w=6u   l=2.3636u ad=24p      pd=14u      as=15p      ps=11u
m17 n2     ci     n4     vss n w=6u   l=2.3636u ad=24p      pd=14u      as=24p      ps=14u
m18 vss    n1     n2     vss n w=6u   l=2.3636u ad=32.7931p pd=17.5862u as=24p      ps=14u
m19 w5     n2     vss    vss n w=6u   l=2.3636u ad=15p      pd=11u      as=32.7931p ps=17.5862u
m20 n1     ci     w5     vss n w=6u   l=2.3636u ad=24p      pd=14u      as=15p      ps=11u
m21 w6     cn     n1     vss n w=6u   l=2.3636u ad=15p      pd=11u      as=24p      ps=14u
m22 vss    d      w6     vss n w=6u   l=2.3636u ad=32.7931p pd=17.5862u as=15p      ps=11u
m23 cn     cp     vss    vss n w=7u   l=2.3636u ad=49p      pd=28u      as=38.2586p ps=20.5172u
C0  cn     vdd    0.069f
C1  w4     n4     0.009f
C2  vss    vdd    0.021f
C3  n4     z      0.034f
C4  ci     n2     0.288f
C5  d      n1     0.048f
C6  cp     d      0.029f
C7  ci     z      0.006f
C8  n4     zn     0.202f
C9  n2     n1     0.327f
C10 d      cn     0.183f
C11 vss    d      0.028f
C12 cp     n2     0.003f
C13 w3     ci     0.006f
C14 d      vdd    0.023f
C15 ci     zn     0.107f
C16 n2     cn     0.162f
C17 vss    n2     0.087f
C18 n2     vdd    0.054f
C19 n1     zn     0.027f
C20 vss    z      0.026f
C21 w2     n1     0.004f
C22 n4     ci     0.218f
C23 z      vdd    0.078f
C24 cn     zn     0.094f
C25 vss    zn     0.047f
C26 n4     n1     0.044f
C27 d      n2     0.040f
C28 zn     vdd    0.031f
C29 n4     cn     0.018f
C30 ci     n1     0.435f
C31 vss    n4     0.152f
C32 w5     n1     0.009f
C33 cp     ci     0.091f
C34 n4     vdd    0.124f
C35 ci     cn     0.417f
C36 cp     n1     0.011f
C37 vss    ci     0.193f
C38 w1     n4     0.010f
C39 ci     vdd    0.164f
C40 n2     zn     0.037f
C41 n1     cn     0.124f
C42 vss    n1     0.202f
C43 cp     cn     0.228f
C44 n1     vdd    0.117f
C45 z      zn     0.134f
C46 cp     vss    0.020f
C47 vss    cn     0.095f
C48 cp     vdd    0.058f
C49 n4     n2     0.110f
C50 d      ci     0.349f
C51 cp     vss    0.030f
C53 n4     vss    0.032f
C54 d      vss    0.028f
C55 ci     vss    0.083f
C56 n2     vss    0.041f
C57 n1     vss    0.036f
C58 z      vss    0.007f
C59 cn     vss    0.109f
C60 zn     vss    0.052f
.ends
