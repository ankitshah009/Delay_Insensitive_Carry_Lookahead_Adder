magic
tech scmos
timestamp 1170759824
<< checkpaint >>
rect -22 -26 118 114
<< ab >>
rect 0 0 96 88
<< pwell >>
rect -4 -8 100 40
<< nwell >>
rect -4 40 100 96
<< polysilicon >>
rect 2 77 11 83
rect 9 74 11 77
rect 21 77 30 83
rect 34 77 43 83
rect 21 74 23 77
rect 41 74 43 77
rect 53 77 62 83
rect 66 82 75 83
rect 66 78 70 82
rect 74 78 75 82
rect 66 77 75 78
rect 53 74 55 77
rect 73 74 75 77
rect 85 82 94 83
rect 85 78 86 82
rect 90 78 94 82
rect 85 77 94 78
rect 85 74 87 77
rect 9 43 11 46
rect 21 43 23 46
rect 41 43 43 46
rect 53 43 55 46
rect 73 43 75 46
rect 85 43 87 46
rect 2 42 14 43
rect 2 38 6 42
rect 10 38 14 42
rect 2 37 14 38
rect 18 42 30 43
rect 18 38 22 42
rect 26 38 30 42
rect 18 37 30 38
rect 34 42 46 43
rect 34 38 41 42
rect 45 38 46 42
rect 34 37 46 38
rect 50 42 62 43
rect 50 38 51 42
rect 55 38 62 42
rect 50 37 62 38
rect 66 42 78 43
rect 66 38 70 42
rect 74 38 78 42
rect 66 37 78 38
rect 82 37 94 43
rect 9 34 11 37
rect 21 34 23 37
rect 41 34 43 37
rect 53 34 55 37
rect 73 34 75 37
rect 85 34 87 37
rect 9 11 11 14
rect 2 5 11 11
rect 21 11 23 14
rect 41 11 43 14
rect 21 5 30 11
rect 34 5 43 11
rect 53 11 55 14
rect 73 11 75 14
rect 53 5 62 11
rect 66 5 75 11
rect 85 11 87 14
rect 85 5 94 11
<< ndiffusion >>
rect 2 26 9 34
rect 2 22 3 26
rect 7 22 9 26
rect 2 19 9 22
rect 2 15 3 19
rect 7 15 9 19
rect 2 14 9 15
rect 11 29 21 34
rect 11 25 14 29
rect 18 25 21 29
rect 11 22 21 25
rect 11 18 14 22
rect 18 18 21 22
rect 11 14 21 18
rect 23 19 30 34
rect 23 15 25 19
rect 29 15 30 19
rect 23 14 30 15
rect 34 19 41 34
rect 34 15 35 19
rect 39 15 41 19
rect 34 14 41 15
rect 43 30 53 34
rect 43 26 46 30
rect 50 26 53 30
rect 43 23 53 26
rect 43 19 46 23
rect 50 19 53 23
rect 43 14 53 19
rect 55 19 62 34
rect 55 15 57 19
rect 61 15 62 19
rect 55 14 62 15
rect 66 19 73 34
rect 66 15 67 19
rect 71 15 73 19
rect 66 14 73 15
rect 75 33 85 34
rect 75 29 78 33
rect 82 29 85 33
rect 75 26 85 29
rect 75 22 78 26
rect 82 22 85 26
rect 75 14 85 22
rect 87 26 94 34
rect 87 22 89 26
rect 93 22 94 26
rect 87 19 94 22
rect 87 15 89 19
rect 93 15 94 19
rect 87 14 94 15
rect 13 2 19 14
rect 45 2 51 14
rect 77 2 83 14
<< pdiffusion >>
rect 13 74 19 86
rect 45 78 51 86
rect 45 74 46 78
rect 50 74 51 78
rect 77 74 83 86
rect 2 73 9 74
rect 2 69 3 73
rect 7 69 9 73
rect 2 66 9 69
rect 2 62 3 66
rect 7 62 9 66
rect 2 46 9 62
rect 11 59 21 74
rect 11 55 14 59
rect 18 55 21 59
rect 11 52 21 55
rect 11 48 14 52
rect 18 48 21 52
rect 11 46 21 48
rect 23 73 30 74
rect 23 69 25 73
rect 29 69 30 73
rect 23 66 30 69
rect 23 62 25 66
rect 29 62 30 66
rect 23 46 30 62
rect 34 61 41 74
rect 34 57 35 61
rect 39 57 41 61
rect 34 52 41 57
rect 34 48 35 52
rect 39 48 41 52
rect 34 46 41 48
rect 43 71 53 74
rect 43 67 46 71
rect 50 67 53 71
rect 43 46 53 67
rect 55 61 62 74
rect 55 57 57 61
rect 61 57 62 61
rect 55 54 62 57
rect 55 50 57 54
rect 61 50 62 54
rect 55 46 62 50
rect 66 70 73 74
rect 66 66 67 70
rect 71 66 73 70
rect 66 46 73 66
rect 75 58 85 74
rect 75 54 78 58
rect 82 54 85 58
rect 75 51 85 54
rect 75 47 78 51
rect 82 47 85 51
rect 75 46 85 47
rect 87 69 94 74
rect 87 65 89 69
rect 93 65 94 69
rect 87 62 94 65
rect 87 58 89 62
rect 93 58 94 62
rect 87 46 94 58
<< metal1 >>
rect -2 86 2 90
rect 10 86 22 90
rect 30 86 34 90
rect 42 86 54 90
rect 62 86 66 90
rect 74 86 86 90
rect 94 86 98 90
rect 3 82 7 86
rect 3 73 7 78
rect 3 66 7 69
rect 3 61 7 62
rect 25 82 29 86
rect 25 73 29 78
rect 25 66 29 69
rect 46 78 50 79
rect 69 78 70 82
rect 74 78 86 82
rect 90 78 91 82
rect 46 71 50 74
rect 50 67 67 70
rect 46 66 67 67
rect 71 69 93 70
rect 71 66 89 69
rect 25 61 29 62
rect 35 61 61 62
rect 14 59 18 60
rect 39 58 57 61
rect 35 55 39 57
rect 6 42 10 55
rect 14 52 39 55
rect 57 54 61 57
rect 18 51 35 52
rect 14 47 18 48
rect 35 47 39 48
rect 21 42 27 46
rect 21 38 22 42
rect 26 38 27 42
rect 40 38 41 42
rect 6 34 27 38
rect 45 34 51 54
rect 57 49 61 50
rect 70 42 74 63
rect 55 38 56 42
rect 61 34 74 38
rect 78 58 82 63
rect 89 62 93 65
rect 89 57 93 58
rect 78 51 82 54
rect 6 33 10 34
rect 78 33 82 47
rect 14 29 46 30
rect 3 26 7 27
rect 3 19 7 22
rect 18 26 46 29
rect 50 29 78 30
rect 50 26 82 29
rect 14 22 18 25
rect 46 23 50 26
rect 14 17 18 18
rect 25 19 29 20
rect 3 10 7 15
rect 3 2 7 6
rect 25 10 29 15
rect 25 2 29 6
rect 35 19 39 20
rect 46 17 50 19
rect 57 19 61 20
rect 35 10 39 15
rect 35 2 39 6
rect 57 10 61 15
rect 57 2 61 6
rect 67 19 71 20
rect 78 17 82 22
rect 89 26 93 27
rect 89 19 93 22
rect 67 10 71 15
rect 67 2 71 6
rect 89 10 93 15
rect 89 2 93 6
rect -2 -2 2 2
rect 10 -2 22 2
rect 30 -2 34 2
rect 42 -2 54 2
rect 62 -2 66 2
rect 74 -2 86 2
rect 94 -2 98 2
<< metal2 >>
rect -2 86 6 90
rect 10 86 22 90
rect 26 86 38 90
rect 42 86 54 90
rect 58 86 70 90
rect 74 86 86 90
rect 90 86 98 90
rect -2 82 98 86
rect -2 78 3 82
rect 7 78 25 82
rect 29 78 98 82
rect -2 76 98 78
rect -2 10 98 12
rect -2 6 3 10
rect 7 6 25 10
rect 29 6 35 10
rect 39 6 57 10
rect 61 6 67 10
rect 71 6 89 10
rect 93 6 98 10
rect -2 2 98 6
rect -2 -2 6 2
rect 10 -2 22 2
rect 26 -2 38 2
rect 42 -2 54 2
rect 58 -2 70 2
rect 74 -2 86 2
rect 90 -2 98 2
<< ntransistor >>
rect 9 14 11 34
rect 21 14 23 34
rect 41 14 43 34
rect 53 14 55 34
rect 73 14 75 34
rect 85 14 87 34
<< ptransistor >>
rect 9 46 11 74
rect 21 46 23 74
rect 41 46 43 74
rect 53 46 55 74
rect 73 46 75 74
rect 85 46 87 74
<< polycontact >>
rect 70 78 74 82
rect 86 78 90 82
rect 6 38 10 42
rect 22 38 26 42
rect 41 38 45 42
rect 51 38 55 42
rect 70 38 74 42
<< ndcontact >>
rect 3 22 7 26
rect 3 15 7 19
rect 14 25 18 29
rect 14 18 18 22
rect 25 15 29 19
rect 35 15 39 19
rect 46 26 50 30
rect 46 19 50 23
rect 57 15 61 19
rect 67 15 71 19
rect 78 29 82 33
rect 78 22 82 26
rect 89 22 93 26
rect 89 15 93 19
<< pdcontact >>
rect 46 74 50 78
rect 3 69 7 73
rect 3 62 7 66
rect 14 55 18 59
rect 14 48 18 52
rect 25 69 29 73
rect 25 62 29 66
rect 35 57 39 61
rect 35 48 39 52
rect 46 67 50 71
rect 57 57 61 61
rect 57 50 61 54
rect 67 66 71 70
rect 78 54 82 58
rect 78 47 82 51
rect 89 65 93 69
rect 89 58 93 62
<< m2contact >>
rect 6 86 10 90
rect 22 86 26 90
rect 38 86 42 90
rect 54 86 58 90
rect 70 86 74 90
rect 86 86 90 90
rect 3 78 7 82
rect 25 78 29 82
rect 3 6 7 10
rect 25 6 29 10
rect 35 6 39 10
rect 57 6 61 10
rect 67 6 71 10
rect 89 6 93 10
rect 6 -2 10 2
rect 22 -2 26 2
rect 38 -2 42 2
rect 54 -2 58 2
rect 70 -2 74 2
rect 86 -2 90 2
<< psubstratepcontact >>
rect 2 -2 6 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 90 -2 94 2
<< nsubstratencontact >>
rect 2 86 6 90
rect 26 86 30 90
rect 34 86 38 90
rect 58 86 62 90
rect 66 86 70 90
rect 90 86 94 90
<< psubstratepdiff >>
rect 0 2 7 3
rect 25 2 39 3
rect 57 2 71 3
rect 89 2 96 3
rect 0 -2 2 2
rect 6 -2 7 2
rect 0 -3 7 -2
rect 25 -2 26 2
rect 30 -2 34 2
rect 38 -2 39 2
rect 25 -3 39 -2
rect 57 -2 58 2
rect 62 -2 66 2
rect 70 -2 71 2
rect 57 -3 71 -2
rect 89 -2 90 2
rect 94 -2 96 2
rect 89 -3 96 -2
<< nsubstratendiff >>
rect 0 90 7 91
rect 0 86 2 90
rect 6 86 7 90
rect 25 90 39 91
rect 25 86 26 90
rect 30 86 34 90
rect 38 86 39 90
rect 57 90 71 91
rect 57 86 58 90
rect 62 86 66 90
rect 70 86 71 90
rect 89 90 96 91
rect 89 86 90 90
rect 94 86 96 90
rect 0 85 7 86
rect 25 85 39 86
rect 57 85 71 86
rect 89 85 96 86
<< labels >>
rlabel metal1 8 44 8 44 6 a
rlabel ndcontact 16 20 16 20 6 z
rlabel metal1 32 28 32 28 6 z
rlabel metal1 24 28 24 28 6 z
rlabel metal1 16 36 16 36 6 a
rlabel polycontact 24 40 24 40 6 a
rlabel metal1 40 28 40 28 6 z
rlabel metal1 56 28 56 28 6 z
rlabel metal1 48 24 48 24 6 z
rlabel metal1 48 44 48 44 6 b
rlabel metal1 72 28 72 28 6 z
rlabel metal1 64 28 64 28 6 z
rlabel metal1 64 36 64 36 6 c
rlabel metal1 72 52 72 52 6 c
rlabel metal1 80 40 80 40 6 z
rlabel metal2 48 6 48 6 6 vss
rlabel metal2 48 82 48 82 6 vdd
<< end >>
