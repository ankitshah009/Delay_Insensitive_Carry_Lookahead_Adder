.subckt iv1v5x6 a vdd vss z
*   SPICE3 file   created from iv1v5x6.ext -      technology: scmos
m00 vdd    a      z      vdd p w=28u  l=2.3636u ad=140p     pd=47.3333u as=130p     ps=47.3333u
m01 z      a      vdd    vdd p w=28u  l=2.3636u ad=130p     pd=47.3333u as=140p     ps=47.3333u
m02 vdd    a      z      vdd p w=28u  l=2.3636u ad=140p     pd=47.3333u as=130p     ps=47.3333u
m03 z      a      vss    vss n w=16u  l=2.3636u ad=64p      pd=24u      as=110.5p   ps=46u
m04 vss    a      z      vss n w=16u  l=2.3636u ad=110.5p   pd=46u      as=64p      ps=24u
C0  vss    z      0.151f
C1  vdd    a      0.028f
C2  vdd    z      0.090f
C3  vss    a      0.059f
C4  z      a      0.193f
C7  z      vss    0.006f
C8  a      vss    0.043f
.ends
