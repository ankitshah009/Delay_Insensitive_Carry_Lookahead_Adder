.subckt aoi21v0x1 a1 a2 b vdd vss z
*   SPICE3 file   created from aoi21v0x1.ext -      technology: scmos
m00 vdd    vdd    w1     vdd p w=28u  l=2.3636u ad=182.667p pd=56.6667u as=196p     ps=70u
m01 w2     a1     vdd    vdd p w=28u  l=2.3636u ad=182.667p pd=56.6667u as=182.667p ps=56.6667u
m02 w2     a2     vdd    vdd p w=28u  l=2.3636u ad=182.667p pd=56.6667u as=182.667p ps=56.6667u
m03 z      b      w2     vdd p w=28u  l=2.3636u ad=196p     pd=70u      as=182.667p ps=56.6667u
m04 vss    vdd    w3     vss n w=20u  l=2.3636u ad=137.333p pd=46u      as=140p     ps=54u
m05 w4     a1     vss    vss n w=20u  l=2.3636u ad=140p     pd=54u      as=137.333p ps=46u
m06 z      a2     w4     vss n w=20u  l=2.3636u ad=136p     pd=42u      as=140p     ps=54u
m07 vss    b      z      vss n w=20u  l=2.3636u ad=137.333p pd=46u      as=136p     ps=42u
C0  b      a1     0.035f
C1  w2     a2     0.029f
C2  vss    z      0.046f
C3  a2     a1     0.141f
C4  w2     vdd    0.195f
C5  w4     w2     0.026f
C6  vss    b      0.045f
C7  a1     vdd    0.075f
C8  z      b      0.222f
C9  vss    a2     0.011f
C10 w4     a1     0.023f
C11 z      a2     0.174f
C12 vss    vdd    0.010f
C13 w4     vss    0.076f
C14 z      vdd    0.018f
C15 b      a2     0.100f
C16 w4     z      0.040f
C17 w2     a1     0.018f
C18 b      vdd    0.022f
C19 w4     b      0.009f
C20 a2     vdd    0.059f
C21 w4     a2     0.023f
C22 w4     vdd    0.003f
C23 vss    a1     0.011f
C24 z      w2     0.078f
C25 z      a1     0.033f
C26 w4     vss    0.004f
C28 z      vss    0.006f
C29 b      vss    0.045f
C30 w2     vss    0.002f
C31 a2     vss    0.045f
C32 a1     vss    0.045f
.ends
