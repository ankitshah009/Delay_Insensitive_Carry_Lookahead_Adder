magic
tech scmos
timestamp 1179386035
<< checkpaint >>
rect -22 -25 46 105
<< ab >>
rect 0 0 24 80
<< pwell >>
rect -4 -7 28 36
<< nwell >>
rect -4 36 28 87
<< polysilicon >>
rect 9 61 11 65
rect 9 39 11 43
rect 9 38 15 39
rect 9 34 10 38
rect 14 34 15 38
rect 9 33 15 34
rect 9 28 11 33
rect 9 15 11 19
<< ndiffusion >>
rect 2 27 9 28
rect 2 23 3 27
rect 7 23 9 27
rect 2 22 9 23
rect 4 19 9 22
rect 11 19 20 28
rect 13 12 20 19
rect 13 8 14 12
rect 18 8 20 12
rect 13 7 20 8
<< pdiffusion >>
rect 13 72 20 73
rect 13 68 14 72
rect 18 68 20 72
rect 13 61 20 68
rect 4 56 9 61
rect 2 55 9 56
rect 2 51 3 55
rect 7 51 9 55
rect 2 48 9 51
rect 2 44 3 48
rect 7 44 9 48
rect 2 43 9 44
rect 11 43 20 61
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect -2 72 26 78
rect -2 68 14 72
rect 18 68 26 72
rect 2 57 14 63
rect 2 55 7 57
rect 2 51 3 55
rect 2 48 7 51
rect 2 44 3 48
rect 2 43 7 44
rect 2 28 6 43
rect 18 39 22 63
rect 10 38 22 39
rect 14 34 22 38
rect 10 33 22 34
rect 2 27 7 28
rect 2 23 3 27
rect 2 17 14 23
rect 18 17 22 33
rect -2 8 14 12
rect 18 8 26 12
rect -2 2 26 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
<< ntransistor >>
rect 9 19 11 28
<< ptransistor >>
rect 9 43 11 61
<< polycontact >>
rect 10 34 14 38
<< ndcontact >>
rect 3 23 7 27
rect 14 8 18 12
<< pdcontact >>
rect 14 68 18 72
rect 3 51 7 55
rect 3 44 7 48
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
<< psubstratepdiff >>
rect 0 2 24 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 24 2
rect 0 -3 24 -2
<< nsubstratendiff >>
rect 0 82 24 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 24 82
rect 0 77 24 78
<< labels >>
rlabel metal1 4 40 4 40 6 z
rlabel metal1 12 6 12 6 6 vss
rlabel metal1 12 20 12 20 6 z
rlabel polycontact 12 36 12 36 6 a
rlabel metal1 12 60 12 60 6 z
rlabel metal1 12 74 12 74 6 vdd
rlabel metal1 20 40 20 40 6 a
<< end >>
