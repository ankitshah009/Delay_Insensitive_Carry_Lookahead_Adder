.subckt nao22_x4 i0 i1 i2 nq vdd vss
*   SPICE3 file   created from nao22_x4.ext -      technology: scmos
m00 w1     i2     vdd    vdd p w=20u  l=2.3636u ad=100p     pd=30u      as=156.571p ps=48.5714u
m01 w2     i1     w1     vdd p w=20u  l=2.3636u ad=100p     pd=30u      as=100p     ps=30u
m02 vdd    i0     w2     vdd p w=20u  l=2.3636u ad=156.571p pd=48.5714u as=100p     ps=30u
m03 vdd    w1     w3     vdd p w=20u  l=2.3636u ad=156.571p pd=48.5714u as=160p     ps=56u
m04 nq     w3     vdd    vdd p w=40u  l=2.3636u ad=200p     pd=50u      as=313.143p ps=97.1429u
m05 vdd    w3     nq     vdd p w=40u  l=2.3636u ad=313.143p pd=97.1429u as=200p     ps=50u
m06 w4     i2     vss    vss n w=10u  l=2.3636u ad=60p      pd=25.3333u as=78p      ps=28u
m07 w1     i1     w4     vss n w=10u  l=2.3636u ad=74p      pd=28u      as=60p      ps=25.3333u
m08 w4     i0     w1     vss n w=10u  l=2.3636u ad=60p      pd=25.3333u as=74p      ps=28u
m09 vss    w1     w3     vss n w=10u  l=2.3636u ad=78p      pd=28u      as=80p      ps=36u
m10 nq     w3     vss    vss n w=20u  l=2.3636u ad=100p     pd=30u      as=156p     ps=56u
m11 vss    w3     nq     vss n w=20u  l=2.3636u ad=156p     pd=56u      as=100p     ps=30u
C0  w4     vss    0.218f
C1  w1     i2     0.356f
C2  w3     i1     0.041f
C3  vss    nq     0.099f
C4  w3     vdd    0.031f
C5  i0     i2     0.088f
C6  w4     w3     0.034f
C7  vss    w1     0.048f
C8  i1     vdd    0.017f
C9  w4     i1     0.017f
C10 w2     w1     0.019f
C11 nq     w3     0.217f
C12 vss    i0     0.028f
C13 w2     i0     0.004f
C14 w1     w3     0.345f
C15 vss    i2     0.055f
C16 nq     vdd    0.231f
C17 w1     i1     0.347f
C18 w3     i0     0.132f
C19 w4     nq     0.006f
C20 w3     i2     0.022f
C21 w1     vdd    0.415f
C22 i0     i1     0.357f
C23 w4     w1     0.117f
C24 i1     i2     0.152f
C25 i0     vdd    0.027f
C26 nq     w1     0.107f
C27 vss    w3     0.193f
C28 w4     i0     0.030f
C29 i2     vdd    0.074f
C30 vss    i1     0.011f
C31 nq     i0     0.044f
C32 w4     i2     0.039f
C33 w1     i0     0.203f
C34 w2     i1     0.016f
C35 vss    vdd    0.005f
C37 nq     vss    0.018f
C38 w1     vss    0.051f
C39 w3     vss    0.068f
C40 i0     vss    0.046f
C41 i1     vss    0.043f
C42 i2     vss    0.052f
.ends
