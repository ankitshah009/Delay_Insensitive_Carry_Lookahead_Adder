magic
tech scmos
timestamp 1179387289
<< checkpaint >>
rect -22 -25 110 105
<< ab >>
rect 0 0 88 80
<< pwell >>
rect -4 -7 92 36
<< nwell >>
rect -4 36 92 87
<< polysilicon >>
rect 9 70 11 74
rect 21 70 23 74
rect 28 70 30 74
rect 35 70 37 74
rect 42 70 44 74
rect 52 70 54 74
rect 59 70 61 74
rect 66 70 68 74
rect 73 70 75 74
rect 21 43 23 46
rect 18 42 24 43
rect 9 33 11 42
rect 18 38 19 42
rect 23 38 24 42
rect 18 37 24 38
rect 9 32 15 33
rect 9 28 10 32
rect 14 28 15 32
rect 9 27 15 28
rect 9 24 11 27
rect 21 22 23 37
rect 28 31 30 46
rect 35 37 37 46
rect 42 43 44 46
rect 52 43 54 46
rect 42 41 55 43
rect 49 38 55 41
rect 35 35 41 37
rect 39 31 41 35
rect 49 34 50 38
rect 54 34 55 38
rect 49 33 55 34
rect 27 30 33 31
rect 27 26 28 30
rect 32 26 33 30
rect 27 25 33 26
rect 39 30 45 31
rect 39 26 40 30
rect 44 26 45 30
rect 39 25 45 26
rect 31 22 33 25
rect 43 22 45 25
rect 53 22 55 33
rect 59 27 61 46
rect 66 37 68 46
rect 73 43 75 46
rect 73 42 82 43
rect 73 41 77 42
rect 76 38 77 41
rect 81 38 82 42
rect 76 37 82 38
rect 65 36 71 37
rect 65 32 66 36
rect 70 32 71 36
rect 65 31 71 32
rect 59 25 67 27
rect 65 23 67 25
rect 65 22 71 23
rect 65 18 66 22
rect 70 18 71 22
rect 65 17 71 18
rect 9 6 11 10
rect 21 10 23 15
rect 31 10 33 15
rect 43 10 45 15
rect 53 10 55 15
<< ndiffusion >>
rect 2 22 9 24
rect 2 18 3 22
rect 7 18 9 22
rect 2 17 9 18
rect 4 10 9 17
rect 11 22 19 24
rect 11 15 21 22
rect 23 21 31 22
rect 23 17 25 21
rect 29 17 31 21
rect 23 15 31 17
rect 33 15 43 22
rect 45 21 53 22
rect 45 17 47 21
rect 51 17 53 21
rect 45 15 53 17
rect 55 15 63 22
rect 11 12 19 15
rect 11 10 14 12
rect 13 8 14 10
rect 18 8 19 12
rect 35 12 41 15
rect 13 7 19 8
rect 35 8 36 12
rect 40 8 41 12
rect 57 12 63 15
rect 35 7 41 8
rect 57 8 58 12
rect 62 8 63 12
rect 57 7 63 8
<< pdiffusion >>
rect 4 55 9 70
rect 2 54 9 55
rect 2 50 3 54
rect 7 50 9 54
rect 2 47 9 50
rect 2 43 3 47
rect 7 43 9 47
rect 2 42 9 43
rect 11 69 21 70
rect 11 65 14 69
rect 18 65 21 69
rect 11 46 21 65
rect 23 46 28 70
rect 30 46 35 70
rect 37 46 42 70
rect 44 62 52 70
rect 44 58 46 62
rect 50 58 52 62
rect 44 46 52 58
rect 54 46 59 70
rect 61 46 66 70
rect 68 46 73 70
rect 75 69 82 70
rect 75 65 77 69
rect 81 65 82 69
rect 75 62 82 65
rect 75 58 77 62
rect 81 58 82 62
rect 75 46 82 58
rect 11 42 16 46
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect -2 69 90 78
rect -2 68 14 69
rect 13 65 14 68
rect 18 68 77 69
rect 18 65 19 68
rect 76 65 77 68
rect 81 68 90 69
rect 81 65 82 68
rect 2 55 6 63
rect 10 58 46 62
rect 50 58 51 62
rect 2 54 7 55
rect 2 50 3 54
rect 2 47 7 50
rect 2 43 3 47
rect 2 42 7 43
rect 2 23 6 42
rect 10 32 14 58
rect 58 54 62 63
rect 76 62 82 65
rect 76 58 77 62
rect 81 58 82 62
rect 18 50 79 54
rect 18 42 23 50
rect 18 38 19 42
rect 18 37 23 38
rect 29 42 70 46
rect 29 31 33 42
rect 41 34 50 38
rect 54 34 55 38
rect 66 36 70 42
rect 74 43 79 50
rect 74 42 82 43
rect 74 38 77 42
rect 81 38 82 42
rect 74 37 82 38
rect 74 33 79 37
rect 66 31 70 32
rect 14 28 22 31
rect 10 27 22 28
rect 2 22 14 23
rect 2 18 3 22
rect 7 18 14 22
rect 2 17 14 18
rect 18 21 22 27
rect 26 30 33 31
rect 26 26 28 30
rect 32 26 33 30
rect 39 26 40 30
rect 44 26 61 30
rect 26 25 33 26
rect 57 22 61 26
rect 18 17 25 21
rect 29 17 47 21
rect 51 17 52 21
rect 57 18 66 22
rect 70 18 71 22
rect -2 8 14 12
rect 18 8 36 12
rect 40 8 58 12
rect 62 8 90 12
rect -2 2 90 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
<< ntransistor >>
rect 9 10 11 24
rect 21 15 23 22
rect 31 15 33 22
rect 43 15 45 22
rect 53 15 55 22
<< ptransistor >>
rect 9 42 11 70
rect 21 46 23 70
rect 28 46 30 70
rect 35 46 37 70
rect 42 46 44 70
rect 52 46 54 70
rect 59 46 61 70
rect 66 46 68 70
rect 73 46 75 70
<< polycontact >>
rect 19 38 23 42
rect 10 28 14 32
rect 50 34 54 38
rect 28 26 32 30
rect 40 26 44 30
rect 77 38 81 42
rect 66 32 70 36
rect 66 18 70 22
<< ndcontact >>
rect 3 18 7 22
rect 25 17 29 21
rect 47 17 51 21
rect 14 8 18 12
rect 36 8 40 12
rect 58 8 62 12
<< pdcontact >>
rect 3 50 7 54
rect 3 43 7 47
rect 14 65 18 69
rect 46 58 50 62
rect 77 65 81 69
rect 77 58 81 62
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
<< psubstratepdiff >>
rect 0 2 88 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 88 2
rect 0 -3 88 -2
<< nsubstratendiff >>
rect 0 82 88 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 88 82
rect 0 77 88 78
<< labels >>
rlabel polycontact 12 30 12 30 6 zn
rlabel metal1 12 20 12 20 6 z
rlabel metal1 4 40 4 40 6 z
rlabel metal1 12 44 12 44 6 zn
rlabel metal1 28 28 28 28 6 b
rlabel metal1 20 44 20 44 6 a
rlabel metal1 28 52 28 52 6 a
rlabel metal1 44 6 44 6 6 vss
rlabel metal1 35 19 35 19 6 zn
rlabel metal1 44 28 44 28 6 c
rlabel metal1 36 44 36 44 6 b
rlabel metal1 44 36 44 36 6 d
rlabel metal1 44 44 44 44 6 b
rlabel metal1 44 52 44 52 6 a
rlabel metal1 36 52 36 52 6 a
rlabel metal1 30 60 30 60 6 zn
rlabel metal1 44 74 44 74 6 vdd
rlabel metal1 52 28 52 28 6 c
rlabel metal1 60 20 60 20 6 c
rlabel polycontact 68 20 68 20 6 c
rlabel polycontact 52 36 52 36 6 d
rlabel metal1 52 44 52 44 6 b
rlabel metal1 60 44 60 44 6 b
rlabel metal1 68 36 68 36 6 b
rlabel metal1 68 52 68 52 6 a
rlabel metal1 52 52 52 52 6 a
rlabel metal1 60 56 60 56 6 a
rlabel metal1 76 44 76 44 6 a
<< end >>
