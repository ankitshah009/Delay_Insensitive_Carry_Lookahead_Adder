magic
tech scmos
timestamp 1179385734
<< checkpaint >>
rect -22 -25 86 105
<< ab >>
rect 0 0 64 80
<< pwell >>
rect -4 -7 68 36
<< nwell >>
rect -4 36 68 87
<< polysilicon >>
rect 12 69 14 74
rect 22 69 24 74
rect 29 69 31 74
rect 39 69 41 74
rect 49 69 51 74
rect 12 39 14 42
rect 22 39 24 42
rect 9 38 24 39
rect 9 34 10 38
rect 14 34 24 38
rect 29 36 31 42
rect 39 39 41 42
rect 49 39 51 42
rect 9 33 24 34
rect 28 33 31 36
rect 35 38 41 39
rect 35 34 36 38
rect 40 34 41 38
rect 35 33 41 34
rect 48 38 55 39
rect 48 34 50 38
rect 54 34 55 38
rect 48 33 55 34
rect 9 28 11 33
rect 21 30 23 33
rect 28 30 30 33
rect 38 30 40 33
rect 48 30 50 33
rect 9 11 11 16
rect 21 13 23 18
rect 28 9 30 18
rect 38 13 40 18
rect 48 9 50 18
rect 28 7 50 9
<< ndiffusion >>
rect 13 28 21 30
rect 4 22 9 28
rect 2 21 9 22
rect 2 17 3 21
rect 7 17 9 21
rect 2 16 9 17
rect 11 18 21 28
rect 23 18 28 30
rect 30 29 38 30
rect 30 25 32 29
rect 36 25 38 29
rect 30 18 38 25
rect 40 23 48 30
rect 40 19 42 23
rect 46 19 48 23
rect 40 18 48 19
rect 50 23 58 30
rect 50 19 52 23
rect 56 19 58 23
rect 50 18 58 19
rect 11 16 19 18
rect 13 12 19 16
rect 13 8 14 12
rect 18 8 19 12
rect 13 7 19 8
<< pdiffusion >>
rect 7 63 12 69
rect 5 62 12 63
rect 5 58 6 62
rect 10 58 12 62
rect 5 55 12 58
rect 5 51 6 55
rect 10 51 12 55
rect 5 50 12 51
rect 7 42 12 50
rect 14 68 22 69
rect 14 64 16 68
rect 20 64 22 68
rect 14 61 22 64
rect 14 57 16 61
rect 20 57 22 61
rect 14 42 22 57
rect 24 42 29 69
rect 31 54 39 69
rect 31 50 33 54
rect 37 50 39 54
rect 31 47 39 50
rect 31 43 33 47
rect 37 43 39 47
rect 31 42 39 43
rect 41 63 49 69
rect 41 59 43 63
rect 47 59 49 63
rect 41 42 49 59
rect 51 68 58 69
rect 51 64 53 68
rect 57 64 58 68
rect 51 60 58 64
rect 51 56 53 60
rect 57 56 58 60
rect 51 42 58 56
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect -2 68 66 78
rect 15 64 16 68
rect 20 64 21 68
rect 6 62 10 63
rect 6 55 10 58
rect 15 61 21 64
rect 15 57 16 61
rect 20 57 21 61
rect 24 59 43 63
rect 47 59 48 63
rect 53 60 57 64
rect 24 54 28 59
rect 53 55 57 56
rect 10 51 28 54
rect 6 50 28 51
rect 33 54 38 55
rect 37 50 38 54
rect 33 47 38 50
rect 2 39 6 47
rect 18 43 33 46
rect 37 43 38 47
rect 18 42 38 43
rect 42 47 46 55
rect 42 42 55 47
rect 2 38 14 39
rect 2 34 10 38
rect 2 33 14 34
rect 18 30 22 42
rect 49 38 55 42
rect 33 34 36 38
rect 40 34 45 38
rect 49 34 50 38
rect 54 34 55 38
rect 41 30 45 34
rect 18 29 37 30
rect 18 25 32 29
rect 36 25 37 29
rect 41 26 55 30
rect 41 21 42 23
rect 2 17 3 21
rect 7 19 42 21
rect 46 19 47 23
rect 7 17 47 19
rect 51 19 52 23
rect 56 19 57 23
rect 51 12 57 19
rect -2 8 14 12
rect 18 8 66 12
rect -2 2 66 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
<< ntransistor >>
rect 9 16 11 28
rect 21 18 23 30
rect 28 18 30 30
rect 38 18 40 30
rect 48 18 50 30
<< ptransistor >>
rect 12 42 14 69
rect 22 42 24 69
rect 29 42 31 69
rect 39 42 41 69
rect 49 42 51 69
<< polycontact >>
rect 10 34 14 38
rect 36 34 40 38
rect 50 34 54 38
<< ndcontact >>
rect 3 17 7 21
rect 32 25 36 29
rect 42 19 46 23
rect 52 19 56 23
rect 14 8 18 12
<< pdcontact >>
rect 6 58 10 62
rect 6 51 10 55
rect 16 64 20 68
rect 16 57 20 61
rect 33 50 37 54
rect 33 43 37 47
rect 43 59 47 63
rect 53 64 57 68
rect 53 56 57 60
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
<< psubstratepdiff >>
rect 0 2 64 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 64 2
rect 0 -3 64 -2
<< nsubstratendiff >>
rect 0 82 64 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 64 82
rect 0 77 64 78
<< labels >>
rlabel metal1 4 40 4 40 6 a
rlabel metal1 8 56 8 56 6 n1
rlabel metal1 20 32 20 32 6 z
rlabel polycontact 12 36 12 36 6 a
rlabel metal1 32 6 32 6 6 vss
rlabel metal1 28 28 28 28 6 z
rlabel metal1 28 44 28 44 6 z
rlabel metal1 36 36 36 36 6 c
rlabel pdcontact 36 52 36 52 6 z
rlabel metal1 32 74 32 74 6 vdd
rlabel metal1 24 19 24 19 6 n3
rlabel metal1 44 28 44 28 6 c
rlabel metal1 44 52 44 52 6 b
rlabel metal1 36 61 36 61 6 n1
rlabel metal1 52 28 52 28 6 c
rlabel metal1 52 40 52 40 6 b
<< end >>
