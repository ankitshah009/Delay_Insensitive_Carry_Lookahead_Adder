magic
tech scmos
timestamp 1179387493
<< checkpaint >>
rect -22 -22 86 94
<< ab >>
rect 0 0 64 72
<< pwell >>
rect -4 -4 68 32
<< nwell >>
rect -4 32 68 76
<< polysilicon >>
rect 11 67 34 69
rect 11 61 13 67
rect 9 59 13 61
rect 22 59 24 63
rect 32 59 34 67
rect 42 66 44 70
rect 49 66 51 70
rect 9 56 11 59
rect 9 35 11 38
rect 22 35 24 41
rect 32 36 34 41
rect 42 35 44 38
rect 49 35 51 38
rect 9 34 18 35
rect 9 33 13 34
rect 12 30 13 33
rect 17 30 18 34
rect 12 29 18 30
rect 22 34 28 35
rect 22 30 23 34
rect 27 30 28 34
rect 22 29 28 30
rect 38 33 44 35
rect 48 34 54 35
rect 2 26 8 27
rect 2 22 3 26
rect 7 22 8 26
rect 15 22 17 29
rect 25 22 27 29
rect 38 27 40 33
rect 48 30 49 34
rect 53 30 54 34
rect 48 29 54 30
rect 48 27 50 29
rect 35 25 40 27
rect 45 25 50 27
rect 35 22 37 25
rect 45 22 47 25
rect 2 21 8 22
rect 4 5 6 21
rect 56 18 62 19
rect 56 14 57 18
rect 61 14 62 18
rect 56 13 62 14
rect 15 9 17 13
rect 25 9 27 13
rect 35 5 37 13
rect 45 9 47 13
rect 56 5 58 13
rect 4 3 58 5
<< ndiffusion >>
rect 10 19 15 22
rect 8 18 15 19
rect 8 14 9 18
rect 13 14 15 18
rect 8 13 15 14
rect 17 18 25 22
rect 17 14 19 18
rect 23 14 25 18
rect 17 13 25 14
rect 27 21 35 22
rect 27 17 29 21
rect 33 17 35 21
rect 27 13 35 17
rect 37 18 45 22
rect 37 14 39 18
rect 43 14 45 18
rect 37 13 45 14
rect 47 19 52 22
rect 47 18 54 19
rect 47 14 49 18
rect 53 14 54 18
rect 47 13 54 14
<< pdiffusion >>
rect 37 59 42 66
rect 15 58 22 59
rect 15 56 16 58
rect 4 51 9 56
rect 2 50 9 51
rect 2 46 3 50
rect 7 46 9 50
rect 2 43 9 46
rect 2 39 3 43
rect 7 39 9 43
rect 2 38 9 39
rect 11 54 16 56
rect 20 54 22 58
rect 11 41 22 54
rect 24 53 32 59
rect 24 49 26 53
rect 30 49 32 53
rect 24 46 32 49
rect 24 42 26 46
rect 30 42 32 46
rect 24 41 32 42
rect 34 50 42 59
rect 34 46 36 50
rect 40 46 42 50
rect 34 41 42 46
rect 11 38 16 41
rect 37 38 42 41
rect 44 38 49 66
rect 51 65 59 66
rect 51 61 53 65
rect 57 61 59 65
rect 51 58 59 61
rect 51 54 53 58
rect 57 54 59 58
rect 51 38 59 54
<< metal1 >>
rect -2 68 66 72
rect -2 64 4 68
rect 8 65 66 68
rect 8 64 53 65
rect 15 58 21 64
rect 15 54 16 58
rect 20 54 21 58
rect 52 61 53 64
rect 57 64 66 65
rect 57 61 58 64
rect 52 58 58 61
rect 52 54 53 58
rect 57 54 58 58
rect 26 53 30 54
rect 2 50 7 51
rect 2 46 3 50
rect 2 43 7 46
rect 18 43 22 51
rect 2 39 3 43
rect 2 38 7 39
rect 10 39 22 43
rect 26 46 30 49
rect 35 46 36 50
rect 40 46 62 50
rect 2 27 6 38
rect 10 37 17 39
rect 26 38 38 42
rect 13 34 17 37
rect 34 34 38 38
rect 13 29 17 30
rect 21 30 23 34
rect 27 30 31 34
rect 34 30 49 34
rect 53 30 54 34
rect 2 26 7 27
rect 21 26 25 30
rect 2 22 3 26
rect 17 22 25 26
rect 34 25 38 30
rect 58 26 62 46
rect 2 18 7 22
rect 29 21 38 25
rect 41 22 62 26
rect 2 14 9 18
rect 13 14 14 18
rect 18 14 19 18
rect 23 14 24 18
rect 41 18 45 22
rect 29 16 33 17
rect 38 14 39 18
rect 43 14 45 18
rect 48 14 49 18
rect 53 14 57 18
rect 61 14 62 18
rect 18 8 24 14
rect -2 0 66 8
<< ntransistor >>
rect 15 13 17 22
rect 25 13 27 22
rect 35 13 37 22
rect 45 13 47 22
<< ptransistor >>
rect 9 38 11 56
rect 22 41 24 59
rect 32 41 34 59
rect 42 38 44 66
rect 49 38 51 66
<< polycontact >>
rect 13 30 17 34
rect 23 30 27 34
rect 3 22 7 26
rect 49 30 53 34
rect 57 14 61 18
<< ndcontact >>
rect 9 14 13 18
rect 19 14 23 18
rect 29 17 33 21
rect 39 14 43 18
rect 49 14 53 18
<< pdcontact >>
rect 3 46 7 50
rect 3 39 7 43
rect 16 54 20 58
rect 26 49 30 53
rect 26 42 30 46
rect 36 46 40 50
rect 53 61 57 65
rect 53 54 57 58
<< nsubstratencontact >>
rect 4 64 8 68
<< nsubstratendiff >>
rect 3 68 9 69
rect 3 64 4 68
rect 8 64 9 68
rect 3 63 9 64
<< labels >>
rlabel polysilicon 5 15 5 15 6 bn
rlabel polycontact 59 16 59 16 6 bn
rlabel ptransistor 50 49 50 49 6 an
rlabel metal1 8 16 8 16 6 bn
rlabel metal1 12 40 12 40 6 b
rlabel metal1 4 32 4 32 6 bn
rlabel metal1 20 24 20 24 6 a
rlabel metal1 28 32 28 32 6 a
rlabel metal1 28 46 28 46 6 an
rlabel metal1 20 48 20 48 6 b
rlabel metal1 32 4 32 4 6 vss
rlabel ndcontact 31 20 31 20 6 an
rlabel metal1 44 24 44 24 6 z
rlabel metal1 44 48 44 48 6 z
rlabel metal1 32 68 32 68 6 vdd
rlabel metal1 55 16 55 16 6 bn
rlabel metal1 52 24 52 24 6 z
rlabel metal1 44 32 44 32 6 an
rlabel metal1 60 36 60 36 6 z
rlabel metal1 52 48 52 48 6 z
<< end >>
