magic
tech scmos
timestamp 1185039102
<< checkpaint >>
rect -22 -24 102 124
<< ab >>
rect 0 0 80 100
<< pwell >>
rect -2 -4 82 49
<< nwell >>
rect -2 49 82 104
<< polysilicon >>
rect 19 95 21 98
rect 27 95 29 98
rect 35 95 37 98
rect 43 95 45 98
rect 55 95 57 98
rect 67 95 69 98
rect 19 53 21 55
rect 17 52 23 53
rect 17 49 18 52
rect 11 48 18 49
rect 22 48 23 52
rect 11 47 23 48
rect 11 25 13 47
rect 27 43 29 55
rect 35 53 37 55
rect 43 53 45 55
rect 55 53 57 55
rect 67 53 69 55
rect 35 51 39 53
rect 43 51 49 53
rect 55 52 69 53
rect 55 51 58 52
rect 37 43 39 51
rect 47 43 49 51
rect 57 48 58 51
rect 62 51 69 52
rect 62 48 63 51
rect 57 47 63 48
rect 27 42 33 43
rect 27 39 28 42
rect 23 38 28 39
rect 32 38 33 42
rect 23 37 33 38
rect 37 42 43 43
rect 37 38 38 42
rect 42 38 43 42
rect 37 37 43 38
rect 47 42 53 43
rect 47 38 48 42
rect 52 38 53 42
rect 47 37 53 38
rect 23 25 25 37
rect 37 29 39 37
rect 47 29 49 37
rect 57 32 63 33
rect 57 29 58 32
rect 33 27 39 29
rect 45 27 49 29
rect 55 28 58 29
rect 62 29 63 32
rect 62 28 69 29
rect 55 27 69 28
rect 33 25 35 27
rect 45 25 47 27
rect 55 25 57 27
rect 67 25 69 27
rect 11 12 13 15
rect 23 12 25 15
rect 33 12 35 15
rect 45 12 47 15
rect 55 2 57 5
rect 67 2 69 5
<< ndiffusion >>
rect 3 15 11 25
rect 13 22 23 25
rect 13 18 16 22
rect 20 18 23 22
rect 13 15 23 18
rect 25 15 33 25
rect 35 22 45 25
rect 35 18 38 22
rect 42 18 45 22
rect 35 15 45 18
rect 47 15 55 25
rect 3 12 9 15
rect 3 8 4 12
rect 8 8 9 12
rect 3 7 9 8
rect 27 9 31 15
rect 49 9 55 15
rect 27 8 33 9
rect 27 4 28 8
rect 32 4 33 8
rect 27 3 33 4
rect 47 8 55 9
rect 47 4 48 8
rect 52 5 55 8
rect 57 22 67 25
rect 57 18 60 22
rect 64 18 67 22
rect 57 5 67 18
rect 69 12 77 25
rect 69 8 72 12
rect 76 8 77 12
rect 69 5 77 8
rect 52 4 53 5
rect 47 3 53 4
<< pdiffusion >>
rect 11 85 19 95
rect 7 82 19 85
rect 7 78 8 82
rect 12 78 19 82
rect 7 72 19 78
rect 7 68 8 72
rect 12 68 19 72
rect 7 62 19 68
rect 7 58 8 62
rect 12 58 19 62
rect 7 55 19 58
rect 21 55 27 95
rect 29 55 35 95
rect 37 55 43 95
rect 45 92 55 95
rect 45 88 48 92
rect 52 88 55 92
rect 45 55 55 88
rect 57 82 67 95
rect 57 78 60 82
rect 64 78 67 82
rect 57 72 67 78
rect 57 68 60 72
rect 64 68 67 72
rect 57 62 67 68
rect 57 58 60 62
rect 64 58 67 62
rect 57 55 67 58
rect 69 92 77 95
rect 69 88 72 92
rect 76 88 77 92
rect 69 82 77 88
rect 69 78 72 82
rect 76 78 77 82
rect 69 72 77 78
rect 69 68 72 72
rect 76 68 77 72
rect 69 55 77 68
<< metal1 >>
rect -2 92 82 101
rect -2 88 48 92
rect 52 88 72 92
rect 76 88 82 92
rect -2 87 82 88
rect 7 82 13 83
rect 59 82 65 83
rect 7 78 8 82
rect 12 78 13 82
rect 7 77 13 78
rect 8 73 12 77
rect 7 72 13 73
rect 7 68 8 72
rect 12 68 13 72
rect 7 67 13 68
rect 8 63 12 67
rect 7 62 13 63
rect 7 58 8 62
rect 12 58 13 62
rect 7 57 13 58
rect 8 23 12 57
rect 17 52 23 82
rect 17 48 18 52
rect 22 48 23 52
rect 17 28 23 48
rect 27 42 33 82
rect 27 38 28 42
rect 32 38 33 42
rect 27 28 33 38
rect 37 42 43 82
rect 37 38 38 42
rect 42 38 43 42
rect 37 28 43 38
rect 47 42 53 82
rect 57 78 60 82
rect 64 78 65 82
rect 57 77 65 78
rect 71 82 77 87
rect 71 78 72 82
rect 76 78 77 82
rect 57 73 63 77
rect 57 72 65 73
rect 57 68 60 72
rect 64 68 65 72
rect 57 67 65 68
rect 71 72 77 78
rect 71 68 72 72
rect 76 68 77 72
rect 71 67 77 68
rect 57 63 63 67
rect 57 62 73 63
rect 57 58 60 62
rect 64 58 73 62
rect 59 57 73 58
rect 57 52 63 53
rect 57 48 58 52
rect 62 48 63 52
rect 57 47 63 48
rect 47 38 48 42
rect 52 38 53 42
rect 47 37 53 38
rect 58 33 62 47
rect 57 32 63 33
rect 48 28 58 32
rect 62 28 63 32
rect 48 23 52 28
rect 57 27 63 28
rect 67 23 73 57
rect 8 22 21 23
rect 37 22 52 23
rect 8 18 16 22
rect 20 18 38 22
rect 42 18 52 22
rect 8 17 21 18
rect 37 17 52 18
rect 59 22 73 23
rect 59 18 60 22
rect 64 18 73 22
rect 59 17 72 18
rect -2 12 82 13
rect -2 8 4 12
rect 8 8 72 12
rect 76 8 82 12
rect -2 4 28 8
rect 32 4 48 8
rect 52 4 82 8
rect -2 -1 82 4
<< ntransistor >>
rect 11 15 13 25
rect 23 15 25 25
rect 33 15 35 25
rect 45 15 47 25
rect 55 5 57 25
rect 67 5 69 25
<< ptransistor >>
rect 19 55 21 95
rect 27 55 29 95
rect 35 55 37 95
rect 43 55 45 95
rect 55 55 57 95
rect 67 55 69 95
<< polycontact >>
rect 18 48 22 52
rect 58 48 62 52
rect 28 38 32 42
rect 38 38 42 42
rect 48 38 52 42
rect 58 28 62 32
<< ndcontact >>
rect 16 18 20 22
rect 38 18 42 22
rect 4 8 8 12
rect 28 4 32 8
rect 48 4 52 8
rect 60 18 64 22
rect 72 8 76 12
<< pdcontact >>
rect 8 78 12 82
rect 8 68 12 72
rect 8 58 12 62
rect 48 88 52 92
rect 60 78 64 82
rect 60 68 64 72
rect 60 58 64 62
rect 72 88 76 92
rect 72 78 76 82
rect 72 68 76 72
<< labels >>
rlabel metal1 20 55 20 55 6 i1
rlabel metal1 20 55 20 55 6 i1
rlabel metal1 30 55 30 55 6 i0
rlabel metal1 30 55 30 55 6 i0
rlabel metal1 40 6 40 6 6 vss
rlabel metal1 40 6 40 6 6 vss
rlabel metal1 40 55 40 55 6 i2
rlabel metal1 40 55 40 55 6 i2
rlabel metal1 60 70 60 70 6 q
rlabel metal1 50 60 50 60 6 i3
rlabel metal1 60 70 60 70 6 q
rlabel metal1 50 60 50 60 6 i3
rlabel metal1 40 94 40 94 6 vdd
rlabel metal1 40 94 40 94 6 vdd
rlabel metal1 70 40 70 40 6 q
rlabel metal1 70 40 70 40 6 q
<< end >>
