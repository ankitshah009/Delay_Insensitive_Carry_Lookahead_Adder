magic
tech scmos
timestamp 1185094785
<< checkpaint >>
rect -22 -22 92 122
<< ab >>
rect 0 0 70 100
<< pwell >>
rect -4 -4 74 48
<< nwell >>
rect -4 48 74 104
<< polysilicon >>
rect 15 94 17 98
rect 27 94 29 98
rect 35 94 37 98
rect 47 94 49 98
rect 55 94 57 98
rect 15 53 17 56
rect 15 52 23 53
rect 15 48 18 52
rect 22 48 23 52
rect 15 47 23 48
rect 27 47 29 56
rect 35 53 37 56
rect 47 53 49 56
rect 35 52 49 53
rect 35 51 38 52
rect 37 48 38 51
rect 42 51 49 52
rect 55 53 57 56
rect 55 52 63 53
rect 42 48 43 51
rect 37 47 43 48
rect 55 48 58 52
rect 62 48 63 52
rect 55 47 63 48
rect 15 38 17 47
rect 27 46 33 47
rect 27 42 28 46
rect 32 42 33 46
rect 27 41 33 42
rect 39 43 43 47
rect 39 41 53 43
rect 27 38 29 41
rect 39 38 41 41
rect 51 38 53 41
rect 39 17 41 22
rect 51 17 53 22
rect 15 2 17 6
rect 27 2 29 6
<< ndiffusion >>
rect 7 37 15 38
rect 7 33 8 37
rect 12 33 15 37
rect 7 29 15 33
rect 7 25 8 29
rect 12 25 15 29
rect 7 24 15 25
rect 10 6 15 24
rect 17 32 27 38
rect 17 28 20 32
rect 24 28 27 32
rect 17 22 27 28
rect 17 18 20 22
rect 24 18 27 22
rect 17 6 27 18
rect 29 22 39 38
rect 41 32 51 38
rect 41 28 44 32
rect 48 28 51 32
rect 41 22 51 28
rect 53 32 62 38
rect 53 28 56 32
rect 60 28 62 32
rect 53 22 62 28
rect 29 18 32 22
rect 36 18 37 22
rect 29 12 37 18
rect 29 8 32 12
rect 36 8 37 12
rect 29 6 37 8
<< pdiffusion >>
rect 10 70 15 94
rect 7 69 15 70
rect 7 65 8 69
rect 12 65 15 69
rect 7 61 15 65
rect 7 57 8 61
rect 12 57 15 61
rect 7 56 15 57
rect 17 92 27 94
rect 17 88 20 92
rect 24 88 27 92
rect 17 82 27 88
rect 17 78 20 82
rect 24 78 27 82
rect 17 56 27 78
rect 29 56 35 94
rect 37 82 47 94
rect 37 78 40 82
rect 44 78 47 82
rect 37 72 47 78
rect 37 68 40 72
rect 44 68 47 72
rect 37 56 47 68
rect 49 56 55 94
rect 57 92 66 94
rect 57 88 60 92
rect 64 88 66 92
rect 57 82 66 88
rect 57 78 60 82
rect 64 78 66 82
rect 57 56 66 78
<< metal1 >>
rect -2 92 72 100
rect -2 88 20 92
rect 24 88 60 92
rect 64 88 72 92
rect 20 82 24 88
rect 20 77 24 78
rect 38 82 44 83
rect 38 78 40 82
rect 38 73 44 78
rect 60 82 64 88
rect 60 77 64 78
rect 8 72 44 73
rect 8 69 40 72
rect 12 68 40 69
rect 12 67 44 68
rect 8 61 12 65
rect 48 63 52 73
rect 8 37 12 57
rect 18 58 33 63
rect 18 52 22 58
rect 18 37 22 48
rect 38 57 52 63
rect 38 52 42 57
rect 38 47 42 48
rect 58 52 63 63
rect 62 48 63 52
rect 27 46 33 47
rect 27 42 28 46
rect 32 42 33 46
rect 58 42 63 48
rect 27 38 63 42
rect 8 29 12 33
rect 56 32 60 33
rect 8 24 12 25
rect 19 28 20 32
rect 24 28 44 32
rect 48 28 49 32
rect 19 22 25 28
rect 19 18 20 22
rect 24 18 25 22
rect 32 22 36 23
rect 32 12 36 18
rect 56 12 60 28
rect -2 8 32 12
rect 36 8 72 12
rect -2 4 48 8
rect 52 4 58 8
rect 62 4 72 8
rect -2 0 72 4
<< ntransistor >>
rect 15 6 17 38
rect 27 6 29 38
rect 39 22 41 38
rect 51 22 53 38
<< ptransistor >>
rect 15 56 17 94
rect 27 56 29 94
rect 35 56 37 94
rect 47 56 49 94
rect 55 56 57 94
<< polycontact >>
rect 18 48 22 52
rect 38 48 42 52
rect 58 48 62 52
rect 28 42 32 46
<< ndcontact >>
rect 8 33 12 37
rect 8 25 12 29
rect 20 28 24 32
rect 20 18 24 22
rect 44 28 48 32
rect 56 28 60 32
rect 32 18 36 22
rect 32 8 36 12
<< pdcontact >>
rect 8 65 12 69
rect 8 57 12 61
rect 20 88 24 92
rect 20 78 24 82
rect 40 78 44 82
rect 40 68 44 72
rect 60 88 64 92
rect 60 78 64 82
<< psubstratepcontact >>
rect 48 4 52 8
rect 58 4 62 8
<< psubstratepdiff >>
rect 47 8 63 9
rect 47 4 48 8
rect 52 4 58 8
rect 62 4 63 8
rect 47 3 63 4
<< labels >>
rlabel metal1 22 25 22 25 6 n3
rlabel metal1 10 50 10 50 6 z
rlabel polycontact 20 50 20 50 6 b
rlabel metal1 20 70 20 70 6 z
rlabel metal1 35 6 35 6 6 vss
rlabel metal1 30 40 30 40 6 a1
rlabel metal1 30 60 30 60 6 b
rlabel metal1 30 70 30 70 6 z
rlabel metal1 35 94 35 94 6 vdd
rlabel metal1 34 30 34 30 6 n3
rlabel metal1 50 40 50 40 6 a1
rlabel metal1 40 40 40 40 6 a1
rlabel metal1 40 55 40 55 6 a2
rlabel metal1 40 75 40 75 6 z
rlabel metal1 50 65 50 65 6 a2
rlabel polycontact 60 50 60 50 6 a1
<< end >>
