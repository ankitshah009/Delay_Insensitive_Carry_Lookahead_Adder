magic
tech scmos
timestamp 1179385298
<< checkpaint >>
rect -22 -25 78 105
<< ab >>
rect 0 0 56 80
<< pwell >>
rect -4 -7 60 36
<< nwell >>
rect -4 36 60 87
<< polysilicon >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 41 70 43 74
rect 9 33 11 43
rect 19 40 21 43
rect 19 39 25 40
rect 19 35 20 39
rect 24 35 25 39
rect 19 34 25 35
rect 29 39 31 43
rect 29 38 35 39
rect 29 34 30 38
rect 34 34 35 38
rect 9 32 15 33
rect 9 28 10 32
rect 14 28 15 32
rect 9 27 15 28
rect 12 23 14 27
rect 20 23 22 34
rect 29 33 35 34
rect 30 23 32 33
rect 41 32 43 43
rect 41 31 47 32
rect 41 28 42 31
rect 38 27 42 28
rect 46 27 47 31
rect 38 26 47 27
rect 38 23 40 26
rect 12 6 14 11
rect 20 6 22 11
rect 30 6 32 11
rect 38 6 40 11
<< ndiffusion >>
rect 3 12 12 23
rect 3 8 5 12
rect 9 11 12 12
rect 14 11 20 23
rect 22 21 30 23
rect 22 17 24 21
rect 28 17 30 21
rect 22 11 30 17
rect 32 11 38 23
rect 40 16 48 23
rect 40 12 42 16
rect 46 12 48 16
rect 40 11 48 12
rect 9 8 10 11
rect 3 7 10 8
<< pdiffusion >>
rect 4 63 9 70
rect 2 62 9 63
rect 2 58 3 62
rect 7 58 9 62
rect 2 57 9 58
rect 4 43 9 57
rect 11 55 19 70
rect 11 51 13 55
rect 17 51 19 55
rect 11 43 19 51
rect 21 62 29 70
rect 21 58 23 62
rect 27 58 29 62
rect 21 43 29 58
rect 31 69 41 70
rect 31 65 34 69
rect 38 65 41 69
rect 31 43 41 65
rect 43 63 48 70
rect 43 62 50 63
rect 43 58 45 62
rect 49 58 50 62
rect 43 57 50 58
rect 43 43 48 57
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect -2 69 58 78
rect -2 68 34 69
rect 33 65 34 68
rect 38 68 58 69
rect 38 65 39 68
rect 2 58 3 62
rect 7 58 23 62
rect 27 58 45 62
rect 49 58 50 62
rect 2 51 13 55
rect 17 51 18 55
rect 2 23 6 51
rect 26 47 30 55
rect 10 32 14 47
rect 18 41 30 47
rect 34 50 47 54
rect 20 39 24 41
rect 20 34 24 35
rect 29 34 30 38
rect 34 33 38 50
rect 42 31 46 39
rect 14 28 22 31
rect 10 27 22 28
rect 18 25 22 27
rect 26 29 30 31
rect 26 27 42 29
rect 26 25 46 27
rect 2 21 14 23
rect 2 17 24 21
rect 28 17 29 21
rect 34 17 38 25
rect 42 16 46 17
rect -2 8 5 12
rect 9 8 58 12
rect -2 2 58 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
<< ntransistor >>
rect 12 11 14 23
rect 20 11 22 23
rect 30 11 32 23
rect 38 11 40 23
<< ptransistor >>
rect 9 43 11 70
rect 19 43 21 70
rect 29 43 31 70
rect 41 43 43 70
<< polycontact >>
rect 20 35 24 39
rect 30 34 34 38
rect 10 28 14 32
rect 42 27 46 31
<< ndcontact >>
rect 5 8 9 12
rect 24 17 28 21
rect 42 12 46 16
<< pdcontact >>
rect 3 58 7 62
rect 13 51 17 55
rect 23 58 27 62
rect 34 65 38 69
rect 45 58 49 62
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
<< psubstratepdiff >>
rect 0 2 56 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 56 2
rect 0 -3 56 -2
<< nsubstratendiff >>
rect 0 82 56 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 56 82
rect 0 77 56 78
<< labels >>
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 20 12 20 6 z
rlabel metal1 12 40 12 40 6 b1
rlabel metal1 28 6 28 6 6 vss
rlabel metal1 20 28 20 28 6 b1
rlabel metal1 28 28 28 28 6 a1
rlabel metal1 20 44 20 44 6 b2
rlabel metal1 28 48 28 48 6 b2
rlabel metal1 28 74 28 74 6 vdd
rlabel metal1 36 20 36 20 6 a1
rlabel metal1 44 32 44 32 6 a1
rlabel metal1 36 40 36 40 6 a2
rlabel metal1 44 52 44 52 6 a2
rlabel pdcontact 26 60 26 60 6 n3
<< end >>
