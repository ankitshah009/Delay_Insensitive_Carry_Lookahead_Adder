magic
tech scmos
timestamp 1179386365
<< checkpaint >>
rect -22 -25 70 105
<< ab >>
rect 0 0 48 80
<< pwell >>
rect -4 -7 52 36
<< nwell >>
rect -4 36 52 87
<< polysilicon >>
rect 9 66 11 71
rect 19 66 21 71
rect 9 39 11 42
rect 19 39 21 42
rect 9 38 15 39
rect 9 34 10 38
rect 14 34 15 38
rect 9 33 15 34
rect 19 38 32 39
rect 19 34 26 38
rect 30 34 32 38
rect 40 38 46 39
rect 40 35 41 38
rect 19 33 32 34
rect 13 30 15 33
rect 20 30 22 33
rect 30 30 32 33
rect 37 34 41 35
rect 45 34 46 38
rect 37 33 46 34
rect 37 30 39 33
rect 13 6 15 10
rect 20 6 22 10
rect 30 6 32 10
rect 37 6 39 10
<< ndiffusion >>
rect 5 15 13 30
rect 5 11 7 15
rect 11 11 13 15
rect 5 10 13 11
rect 15 10 20 30
rect 22 22 30 30
rect 22 18 24 22
rect 28 18 30 22
rect 22 10 30 18
rect 32 10 37 30
rect 39 22 46 30
rect 39 18 41 22
rect 45 18 46 22
rect 39 15 46 18
rect 39 11 41 15
rect 45 11 46 15
rect 39 10 46 11
<< pdiffusion >>
rect 2 65 9 66
rect 2 61 3 65
rect 7 61 9 65
rect 2 57 9 61
rect 2 53 3 57
rect 7 53 9 57
rect 2 42 9 53
rect 11 54 19 66
rect 11 50 13 54
rect 17 50 19 54
rect 11 47 19 50
rect 11 43 13 47
rect 17 43 19 47
rect 11 42 19 43
rect 21 65 29 66
rect 21 61 23 65
rect 27 61 29 65
rect 21 57 29 61
rect 21 53 23 57
rect 27 53 29 57
rect 21 42 29 53
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect -2 68 50 78
rect 3 65 7 68
rect 3 57 7 61
rect 23 65 27 68
rect 23 57 27 61
rect 3 52 7 53
rect 12 50 13 54
rect 17 50 18 54
rect 23 52 27 53
rect 12 47 18 50
rect 2 43 13 47
rect 17 43 18 47
rect 2 22 6 43
rect 25 42 39 46
rect 10 38 19 39
rect 14 34 19 38
rect 25 38 31 42
rect 25 34 26 38
rect 30 34 31 38
rect 40 34 41 38
rect 45 34 46 38
rect 10 33 19 34
rect 15 30 19 33
rect 40 30 46 34
rect 15 26 46 30
rect 2 18 24 22
rect 28 18 31 22
rect 40 18 41 22
rect 45 18 46 22
rect 40 15 46 18
rect 6 12 7 15
rect -2 11 7 12
rect 11 12 12 15
rect 40 12 41 15
rect 11 11 41 12
rect 45 12 46 15
rect 45 11 50 12
rect -2 2 50 11
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
<< ntransistor >>
rect 13 10 15 30
rect 20 10 22 30
rect 30 10 32 30
rect 37 10 39 30
<< ptransistor >>
rect 9 42 11 66
rect 19 42 21 66
<< polycontact >>
rect 10 34 14 38
rect 26 34 30 38
rect 41 34 45 38
<< ndcontact >>
rect 7 11 11 15
rect 24 18 28 22
rect 41 18 45 22
rect 41 11 45 15
<< pdcontact >>
rect 3 61 7 65
rect 3 53 7 57
rect 13 50 17 54
rect 13 43 17 47
rect 23 61 27 65
rect 23 53 27 57
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
<< psubstratepdiff >>
rect 0 2 48 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 48 2
rect 0 -3 48 -2
<< nsubstratendiff >>
rect 0 82 48 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 48 82
rect 0 77 48 78
<< labels >>
rlabel metal1 4 36 4 36 6 z
rlabel metal1 20 20 20 20 6 z
rlabel metal1 12 20 12 20 6 z
rlabel polycontact 12 36 12 36 6 a
rlabel metal1 20 28 20 28 6 a
rlabel metal1 24 6 24 6 6 vss
rlabel metal1 28 20 28 20 6 z
rlabel metal1 28 28 28 28 6 a
rlabel metal1 28 40 28 40 6 b
rlabel metal1 24 74 24 74 6 vdd
rlabel metal1 36 28 36 28 6 a
rlabel metal1 36 44 36 44 6 b
<< end >>
