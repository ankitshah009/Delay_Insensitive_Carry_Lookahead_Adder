.subckt nd2_x2 a b vdd vss z
*   SPICE3 file   created from nd2_x2.ext -      technology: scmos
m00 z      b      vdd    vdd p w=39u  l=2.3636u ad=195p     pd=49u      as=351p     ps=96u
m01 vdd    a      z      vdd p w=39u  l=2.3636u ad=351p     pd=96u      as=195p     ps=49u
m02 w1     b      z      vss n w=33u  l=2.3636u ad=99p      pd=39u      as=207p     ps=82u
m03 vss    a      w1     vss n w=33u  l=2.3636u ad=297p     pd=84u      as=99p      ps=39u
C0  vdd    b      0.034f
C1  vss    w1     0.011f
C2  vss    b      0.012f
C3  w1     a      0.004f
C4  z      vdd    0.177f
C5  z      b      0.183f
C6  vdd    a      0.008f
C7  a      b      0.194f
C8  vss    z      0.057f
C9  vss    a      0.062f
C10 z      a      0.077f
C12 z      vss    0.013f
C14 a      vss    0.024f
C15 b      vss    0.017f
.ends
