.subckt oa2ao222_x4 i0 i1 i2 i3 i4 q vdd vss
*   SPICE3 file   created from oa2ao222_x4.ext -      technology: scmos
m00 vdd    i0     w1     vdd p w=29u  l=2.3636u ad=206.783p pd=60.5217u as=193.123p ps=56.7391u
m01 w1     i1     vdd    vdd p w=29u  l=2.3636u ad=193.123p pd=56.7391u as=206.783p ps=60.5217u
m02 w2     i4     w1     vdd p w=40u  l=2.3636u ad=200p     pd=50u      as=266.377p ps=78.2609u
m03 w3     i2     w2     vdd p w=40u  l=2.3636u ad=160p     pd=48u      as=200p     ps=50u
m04 w1     i3     w3     vdd p w=40u  l=2.3636u ad=266.377p pd=78.2609u as=160p     ps=48u
m05 q      w2     vdd    vdd p w=40u  l=2.3636u ad=200p     pd=50u      as=285.217p ps=83.4783u
m06 vdd    w2     q      vdd p w=40u  l=2.3636u ad=285.217p pd=83.4783u as=200p     ps=50u
m07 w4     i0     vss    vss n w=18u  l=2.3636u ad=72p      pd=26u      as=162.439p ps=57.0732u
m08 w2     i1     w4     vss n w=18u  l=2.3636u ad=100.8p   pd=33.6u    as=72p      ps=26u
m09 w5     i4     w2     vss n w=12u  l=2.3636u ad=96p      pd=36u      as=67.2p    ps=22.4u
m10 vss    i2     w5     vss n w=12u  l=2.3636u ad=108.293p pd=38.0488u as=96p      ps=36u
m11 w5     i3     vss    vss n w=12u  l=2.3636u ad=96p      pd=36u      as=108.293p ps=38.0488u
m12 q      w2     vss    vss n w=20u  l=2.3636u ad=100p     pd=30u      as=180.488p ps=63.4146u
m13 vss    w2     q      vss n w=20u  l=2.3636u ad=180.488p pd=63.4146u as=100p     ps=30u
C0  vss    w2     0.112f
C1  w5     i2     0.033f
C2  w1     i1     0.036f
C3  q      vdd    0.313f
C4  i3     i4     0.052f
C5  w5     vss    0.261f
C6  q      i3     0.044f
C7  i1     i0     0.398f
C8  vss    i2     0.036f
C9  w1     vdd    0.508f
C10 w3     w2     0.016f
C11 i1     w2     0.109f
C12 i0     vdd    0.023f
C13 w1     i3     0.029f
C14 w3     i2     0.012f
C15 i1     i2     0.057f
C16 w1     i4     0.086f
C17 vdd    w2     0.211f
C18 q      w1     0.010f
C19 vss    i1     0.013f
C20 w4     i0     0.009f
C21 vdd    i2     0.012f
C22 i0     i4     0.094f
C23 w2     i3     0.169f
C24 vss    vdd    0.008f
C25 w5     i3     0.047f
C26 i3     i2     0.322f
C27 w2     i4     0.268f
C28 w1     i0     0.064f
C29 vss    i3     0.036f
C30 w3     vdd    0.019f
C31 q      w2     0.221f
C32 i2     i4     0.094f
C33 w5     q      0.012f
C34 w3     i3     0.004f
C35 i1     vdd    0.050f
C36 vss    i4     0.009f
C37 w1     w2     0.194f
C38 q      i2     0.031f
C39 vss    q      0.262f
C40 i0     w2     0.079f
C41 i1     i3     0.040f
C42 w1     i2     0.017f
C43 w5     i0     0.006f
C44 w4     i1     0.012f
C45 i1     i4     0.314f
C46 i0     i2     0.040f
C47 vdd    i3     0.017f
C48 w3     w1     0.016f
C49 w5     w2     0.087f
C50 vss    i0     0.063f
C51 vdd    i4     0.017f
C52 w2     i2     0.281f
C53 w5     vss    0.005f
C55 q      vss    0.010f
C56 i1     vss    0.024f
C57 i0     vss    0.023f
C59 w2     vss    0.056f
C60 i3     vss    0.023f
C61 i2     vss    0.024f
C62 i4     vss    0.028f
.ends
