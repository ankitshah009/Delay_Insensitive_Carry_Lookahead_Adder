magic
tech scmos
timestamp 1179385145
<< checkpaint >>
rect -22 -25 86 105
<< ab >>
rect 0 0 64 80
<< pwell >>
rect -4 -7 68 36
<< nwell >>
rect -4 36 68 87
<< polysilicon >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 41 70 43 74
rect 51 70 53 74
rect 9 34 11 42
rect 19 39 21 53
rect 29 47 31 53
rect 41 50 43 53
rect 41 49 47 50
rect 29 46 37 47
rect 29 42 31 46
rect 35 42 37 46
rect 41 45 42 49
rect 46 45 47 49
rect 41 44 47 45
rect 29 41 37 42
rect 19 38 25 39
rect 19 34 20 38
rect 24 35 25 38
rect 24 34 30 35
rect 9 33 15 34
rect 19 33 30 34
rect 9 29 10 33
rect 14 29 15 33
rect 28 30 30 33
rect 35 30 37 41
rect 42 30 44 44
rect 51 39 53 53
rect 49 38 62 39
rect 49 34 57 38
rect 61 34 62 38
rect 49 33 62 34
rect 49 30 51 33
rect 9 28 15 29
rect 9 25 11 28
rect 9 6 11 11
rect 28 6 30 10
rect 35 6 37 10
rect 42 6 44 10
rect 49 6 51 10
<< ndiffusion >>
rect 21 29 28 30
rect 21 25 22 29
rect 26 25 28 29
rect 4 23 9 25
rect 2 22 9 23
rect 2 18 3 22
rect 7 18 9 22
rect 2 17 9 18
rect 4 11 9 17
rect 11 20 17 25
rect 21 24 28 25
rect 11 12 19 20
rect 11 11 14 12
rect 13 8 14 11
rect 18 8 19 12
rect 23 10 28 24
rect 30 10 35 30
rect 37 10 42 30
rect 44 10 49 30
rect 51 22 58 30
rect 51 18 53 22
rect 57 18 58 22
rect 51 15 58 18
rect 51 11 53 15
rect 57 11 58 15
rect 51 10 58 11
rect 13 7 19 8
<< pdiffusion >>
rect 4 55 9 70
rect 2 54 9 55
rect 2 50 3 54
rect 7 50 9 54
rect 2 47 9 50
rect 2 43 3 47
rect 7 43 9 47
rect 2 42 9 43
rect 11 69 19 70
rect 11 65 13 69
rect 17 65 19 69
rect 11 62 19 65
rect 11 58 13 62
rect 17 58 19 62
rect 11 53 19 58
rect 21 62 29 70
rect 21 58 23 62
rect 27 58 29 62
rect 21 53 29 58
rect 31 69 41 70
rect 31 65 34 69
rect 38 65 41 69
rect 31 53 41 65
rect 43 62 51 70
rect 43 58 45 62
rect 49 58 51 62
rect 43 53 51 58
rect 53 69 60 70
rect 53 65 55 69
rect 59 65 60 69
rect 53 61 60 65
rect 53 57 55 61
rect 59 57 60 61
rect 53 53 60 57
rect 11 42 17 53
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect -2 69 66 78
rect -2 68 13 69
rect 12 65 13 68
rect 17 68 34 69
rect 17 65 18 68
rect 33 65 34 68
rect 38 68 55 69
rect 38 65 39 68
rect 59 68 66 69
rect 2 54 7 63
rect 12 62 18 65
rect 12 58 13 62
rect 17 58 18 62
rect 22 58 23 62
rect 27 58 45 62
rect 49 58 50 62
rect 55 61 59 65
rect 22 54 26 58
rect 55 56 59 57
rect 2 50 3 54
rect 2 47 7 50
rect 2 43 3 47
rect 2 42 7 43
rect 10 50 26 54
rect 2 23 6 42
rect 10 33 14 50
rect 34 46 38 55
rect 17 42 31 46
rect 35 42 38 46
rect 42 49 46 55
rect 46 45 54 47
rect 42 41 54 45
rect 17 34 20 38
rect 24 34 38 38
rect 14 29 27 30
rect 10 26 22 29
rect 21 25 22 26
rect 26 25 27 29
rect 2 22 14 23
rect 2 18 3 22
rect 7 18 14 22
rect 2 17 14 18
rect 34 17 38 34
rect 42 33 46 41
rect 58 38 62 39
rect 56 34 57 38
rect 61 34 62 38
rect 56 31 62 34
rect 50 29 62 31
rect 42 25 62 29
rect 42 17 46 25
rect 52 18 53 22
rect 57 18 58 22
rect 52 15 58 18
rect 52 12 53 15
rect -2 8 14 12
rect 18 11 53 12
rect 57 12 58 15
rect 57 11 66 12
rect 18 8 66 11
rect -2 2 66 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
<< ntransistor >>
rect 9 11 11 25
rect 28 10 30 30
rect 35 10 37 30
rect 42 10 44 30
rect 49 10 51 30
<< ptransistor >>
rect 9 42 11 70
rect 19 53 21 70
rect 29 53 31 70
rect 41 53 43 70
rect 51 53 53 70
<< polycontact >>
rect 31 42 35 46
rect 42 45 46 49
rect 20 34 24 38
rect 10 29 14 33
rect 57 34 61 38
<< ndcontact >>
rect 22 25 26 29
rect 3 18 7 22
rect 14 8 18 12
rect 53 18 57 22
rect 53 11 57 15
<< pdcontact >>
rect 3 50 7 54
rect 3 43 7 47
rect 13 65 17 69
rect 13 58 17 62
rect 23 58 27 62
rect 34 65 38 69
rect 45 58 49 62
rect 55 65 59 69
rect 55 57 59 61
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
<< psubstratepdiff >>
rect 0 2 64 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 64 2
rect 0 -3 64 -2
<< nsubstratendiff >>
rect 0 82 64 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 64 82
rect 0 77 64 78
<< labels >>
rlabel polycontact 12 31 12 31 6 zn
rlabel metal1 4 40 4 40 6 z
rlabel metal1 12 20 12 20 6 z
rlabel metal1 20 44 20 44 6 c
rlabel metal1 20 36 20 36 6 d
rlabel metal1 12 40 12 40 6 zn
rlabel metal1 32 6 32 6 6 vss
rlabel ndcontact 24 27 24 27 6 zn
rlabel metal1 36 24 36 24 6 d
rlabel metal1 28 36 28 36 6 d
rlabel metal1 28 44 28 44 6 c
rlabel metal1 36 52 36 52 6 c
rlabel metal1 32 74 32 74 6 vdd
rlabel metal1 44 20 44 20 6 a
rlabel metal1 44 44 44 44 6 b
rlabel metal1 36 60 36 60 6 zn
rlabel metal1 52 28 52 28 6 a
rlabel metal1 60 32 60 32 6 a
rlabel metal1 52 44 52 44 6 b
<< end >>
