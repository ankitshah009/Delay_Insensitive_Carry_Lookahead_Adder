.subckt noa22_x4 i0 i1 i2 nq vdd vss
*   SPICE3 file   created from noa22_x4.ext -      technology: scmos
m00 w1     i2     vdd    vdd p w=20u  l=2.3636u ad=120p     pd=38.6667u as=147.288p ps=44.7458u
m01 w2     i1     w1     vdd p w=20u  l=2.3636u ad=100p     pd=30u      as=120p     ps=38.6667u
m02 w1     i0     w2     vdd p w=20u  l=2.3636u ad=120p     pd=38.6667u as=100p     ps=30u
m03 vdd    w2     w3     vdd p w=20u  l=2.3636u ad=147.288p pd=44.7458u as=160p     ps=56u
m04 nq     w3     vdd    vdd p w=39u  l=2.3636u ad=195p     pd=49u      as=287.212p ps=87.2542u
m05 vdd    w3     nq     vdd p w=39u  l=2.3636u ad=287.212p pd=87.2542u as=195p     ps=49u
m06 w2     i2     vss    vss n w=10u  l=2.3636u ad=50p      pd=20u      as=85.2941p ps=31.7647u
m07 w4     i1     w2     vss n w=10u  l=2.3636u ad=50p      pd=20u      as=50p      ps=20u
m08 vss    i0     w4     vss n w=10u  l=2.3636u ad=85.2941p pd=31.7647u as=50p      ps=20u
m09 vss    w2     w3     vss n w=10u  l=2.3636u ad=85.2941p pd=31.7647u as=80p      ps=36u
m10 nq     w3     vss    vss n w=19u  l=2.3636u ad=95p      pd=29u      as=162.059p ps=60.3529u
m11 vss    w3     nq     vss n w=19u  l=2.3636u ad=162.059p pd=60.3529u as=95p      ps=29u
C0  w3     vdd    0.025f
C1  vss    i2     0.044f
C2  w2     i0     0.166f
C3  w1     i1     0.013f
C4  w2     i2     0.278f
C5  nq     w3     0.105f
C6  vss    vdd    0.004f
C7  w2     vdd    0.168f
C8  i0     i2     0.090f
C9  vss    nq     0.089f
C10 i0     vdd    0.007f
C11 i1     w3     0.066f
C12 nq     w2     0.076f
C13 i2     vdd    0.064f
C14 w2     w1     0.201f
C15 nq     i0     0.039f
C16 vss    i1     0.034f
C17 w2     i1     0.295f
C18 w1     i0     0.013f
C19 vss    w3     0.083f
C20 i0     i1     0.327f
C21 w2     w3     0.309f
C22 nq     vdd    0.165f
C23 w1     i2     0.024f
C24 i0     w3     0.132f
C25 w1     vdd    0.174f
C26 i1     i2     0.167f
C27 vss    w2     0.036f
C28 i1     vdd    0.008f
C29 i2     w3     0.033f
C30 nq     w1     0.004f
C31 vss    i0     0.046f
C32 w4     i1     0.018f
C34 nq     vss    0.012f
C35 w2     vss    0.048f
C36 i0     vss    0.037f
C37 i1     vss    0.043f
C38 i2     vss    0.044f
C39 w3     vss    0.071f
.ends
