magic
tech scmos
timestamp 1179386834
<< checkpaint >>
rect -22 -22 150 94
<< ab >>
rect 0 0 128 72
<< pwell >>
rect -4 -4 132 32
<< nwell >>
rect -4 32 132 76
<< polysilicon >>
rect 9 66 11 70
rect 16 66 18 70
rect 26 66 28 70
rect 33 66 35 70
rect 43 66 45 70
rect 50 66 52 70
rect 60 66 62 70
rect 67 66 69 70
rect 77 66 79 70
rect 84 66 86 70
rect 94 66 96 70
rect 101 66 103 70
rect 9 29 11 38
rect 16 35 18 38
rect 26 35 28 38
rect 33 35 35 38
rect 43 35 45 38
rect 50 35 52 38
rect 60 35 62 38
rect 67 35 69 38
rect 77 35 79 38
rect 84 35 86 38
rect 94 35 96 38
rect 16 34 29 35
rect 16 33 24 34
rect 23 30 24 33
rect 28 30 29 34
rect 33 34 45 35
rect 33 33 38 34
rect 23 29 29 30
rect 37 30 38 33
rect 42 30 45 34
rect 37 29 45 30
rect 49 34 63 35
rect 49 30 50 34
rect 54 30 63 34
rect 67 34 79 35
rect 67 33 74 34
rect 49 29 63 30
rect 9 28 19 29
rect 9 27 14 28
rect 13 24 14 27
rect 18 25 19 28
rect 39 26 41 29
rect 49 26 51 29
rect 61 26 63 29
rect 71 30 74 33
rect 78 30 79 34
rect 71 29 79 30
rect 83 34 96 35
rect 83 30 90 34
rect 94 30 96 34
rect 83 29 96 30
rect 101 35 103 38
rect 101 34 107 35
rect 101 30 102 34
rect 106 30 107 34
rect 101 29 107 30
rect 71 26 73 29
rect 83 26 85 29
rect 93 26 95 29
rect 105 26 107 29
rect 18 24 29 25
rect 13 23 29 24
rect 17 20 19 23
rect 27 20 29 23
rect 17 5 19 10
rect 27 5 29 10
rect 39 2 41 6
rect 49 2 51 6
rect 61 2 63 6
rect 71 2 73 6
rect 83 2 85 6
rect 93 2 95 6
rect 105 2 107 6
<< ndiffusion >>
rect 31 20 39 26
rect 8 10 17 20
rect 19 18 27 20
rect 19 14 21 18
rect 25 14 27 18
rect 19 10 27 14
rect 29 10 39 20
rect 8 8 15 10
rect 8 4 10 8
rect 14 4 15 8
rect 31 8 39 10
rect 8 3 15 4
rect 31 4 32 8
rect 36 6 39 8
rect 41 18 49 26
rect 41 14 43 18
rect 47 14 49 18
rect 41 6 49 14
rect 51 8 61 26
rect 51 6 54 8
rect 36 4 37 6
rect 31 3 37 4
rect 53 4 54 6
rect 58 6 61 8
rect 63 18 71 26
rect 63 14 65 18
rect 69 14 71 18
rect 63 6 71 14
rect 73 8 83 26
rect 73 6 76 8
rect 58 4 59 6
rect 53 3 59 4
rect 75 4 76 6
rect 80 6 83 8
rect 85 18 93 26
rect 85 14 87 18
rect 91 14 93 18
rect 85 6 93 14
rect 95 8 105 26
rect 95 6 98 8
rect 80 4 81 6
rect 75 3 81 4
rect 97 4 98 6
rect 102 6 105 8
rect 107 25 114 26
rect 107 21 109 25
rect 113 21 114 25
rect 107 18 114 21
rect 107 14 109 18
rect 113 14 114 18
rect 107 13 114 14
rect 107 6 112 13
rect 102 4 103 6
rect 97 3 103 4
<< pdiffusion >>
rect 2 65 9 66
rect 2 61 3 65
rect 7 61 9 65
rect 2 58 9 61
rect 2 54 3 58
rect 7 54 9 58
rect 2 38 9 54
rect 11 38 16 66
rect 18 58 26 66
rect 18 54 20 58
rect 24 54 26 58
rect 18 50 26 54
rect 18 46 20 50
rect 24 46 26 50
rect 18 38 26 46
rect 28 38 33 66
rect 35 65 43 66
rect 35 61 37 65
rect 41 61 43 65
rect 35 58 43 61
rect 35 54 37 58
rect 41 54 43 58
rect 35 38 43 54
rect 45 38 50 66
rect 52 57 60 66
rect 52 53 54 57
rect 58 53 60 57
rect 52 50 60 53
rect 52 46 54 50
rect 58 46 60 50
rect 52 38 60 46
rect 62 38 67 66
rect 69 65 77 66
rect 69 61 71 65
rect 75 61 77 65
rect 69 58 77 61
rect 69 54 71 58
rect 75 54 77 58
rect 69 38 77 54
rect 79 38 84 66
rect 86 58 94 66
rect 86 54 88 58
rect 92 54 94 58
rect 86 50 94 54
rect 86 46 88 50
rect 92 46 94 50
rect 86 38 94 46
rect 96 38 101 66
rect 103 65 110 66
rect 103 61 105 65
rect 109 61 110 65
rect 103 58 110 61
rect 103 54 105 58
rect 109 54 110 58
rect 103 38 110 54
<< metal1 >>
rect -2 68 130 72
rect -2 65 115 68
rect -2 64 3 65
rect 2 61 3 64
rect 7 64 37 65
rect 7 61 8 64
rect 2 58 8 61
rect 36 61 37 64
rect 41 64 71 65
rect 41 61 42 64
rect 2 54 3 58
rect 7 54 8 58
rect 18 58 24 59
rect 18 54 20 58
rect 36 58 42 61
rect 70 61 71 64
rect 75 64 105 65
rect 75 61 76 64
rect 70 58 76 61
rect 104 61 105 64
rect 109 64 115 65
rect 119 64 130 68
rect 109 61 110 64
rect 36 54 37 58
rect 41 54 42 58
rect 54 57 58 58
rect 18 50 24 54
rect 70 54 71 58
rect 75 54 76 58
rect 88 58 94 59
rect 92 54 94 58
rect 104 58 110 61
rect 104 54 105 58
rect 109 54 110 58
rect 54 50 58 53
rect 88 50 94 54
rect 2 46 20 50
rect 24 46 54 50
rect 58 46 88 50
rect 92 46 94 50
rect 2 18 6 46
rect 27 38 103 42
rect 27 34 31 38
rect 49 34 55 38
rect 89 34 95 38
rect 23 30 24 34
rect 28 30 31 34
rect 37 30 38 34
rect 42 30 43 34
rect 49 30 50 34
rect 54 30 55 34
rect 73 30 74 34
rect 78 30 79 34
rect 89 30 90 34
rect 94 30 95 34
rect 99 30 102 34
rect 106 30 111 34
rect 14 28 18 29
rect 37 26 43 30
rect 73 26 79 30
rect 99 26 103 30
rect 18 24 103 26
rect 14 22 103 24
rect 109 25 113 26
rect 109 18 113 21
rect 2 14 21 18
rect 25 14 43 18
rect 47 14 65 18
rect 69 14 87 18
rect 91 14 109 18
rect 113 14 119 18
rect -2 4 10 8
rect 14 4 32 8
rect 36 4 54 8
rect 58 4 76 8
rect 80 4 98 8
rect 102 4 120 8
rect 124 4 130 8
rect -2 0 130 4
<< ntransistor >>
rect 17 10 19 20
rect 27 10 29 20
rect 39 6 41 26
rect 49 6 51 26
rect 61 6 63 26
rect 71 6 73 26
rect 83 6 85 26
rect 93 6 95 26
rect 105 6 107 26
<< ptransistor >>
rect 9 38 11 66
rect 16 38 18 66
rect 26 38 28 66
rect 33 38 35 66
rect 43 38 45 66
rect 50 38 52 66
rect 60 38 62 66
rect 67 38 69 66
rect 77 38 79 66
rect 84 38 86 66
rect 94 38 96 66
rect 101 38 103 66
<< polycontact >>
rect 24 30 28 34
rect 38 30 42 34
rect 50 30 54 34
rect 14 24 18 28
rect 74 30 78 34
rect 90 30 94 34
rect 102 30 106 34
<< ndcontact >>
rect 21 14 25 18
rect 10 4 14 8
rect 32 4 36 8
rect 43 14 47 18
rect 54 4 58 8
rect 65 14 69 18
rect 76 4 80 8
rect 87 14 91 18
rect 98 4 102 8
rect 109 21 113 25
rect 109 14 113 18
<< pdcontact >>
rect 3 61 7 65
rect 3 54 7 58
rect 20 54 24 58
rect 20 46 24 50
rect 37 61 41 65
rect 37 54 41 58
rect 54 53 58 57
rect 54 46 58 50
rect 71 61 75 65
rect 71 54 75 58
rect 88 54 92 58
rect 88 46 92 50
rect 105 61 109 65
rect 105 54 109 58
<< psubstratepcontact >>
rect 120 4 124 8
<< nsubstratencontact >>
rect 115 64 119 68
<< psubstratepdiff >>
rect 119 8 125 24
rect 119 4 120 8
rect 124 4 125 8
rect 119 3 125 4
<< nsubstratendiff >>
rect 114 68 120 69
rect 114 64 115 68
rect 119 64 120 68
rect 114 40 120 64
<< labels >>
rlabel metal1 20 16 20 16 6 z
rlabel metal1 12 16 12 16 6 z
rlabel metal1 20 24 20 24 6 a
rlabel metal1 4 32 4 32 6 z
rlabel metal1 20 52 20 52 6 z
rlabel metal1 12 48 12 48 6 z
rlabel ndcontact 44 16 44 16 6 z
rlabel metal1 36 16 36 16 6 z
rlabel metal1 28 16 28 16 6 z
rlabel metal1 44 24 44 24 6 a
rlabel metal1 36 24 36 24 6 a
rlabel metal1 28 24 28 24 6 a
rlabel metal1 28 32 28 32 6 b
rlabel metal1 44 40 44 40 6 b
rlabel metal1 36 40 36 40 6 b
rlabel metal1 44 48 44 48 6 z
rlabel metal1 36 48 36 48 6 z
rlabel metal1 28 48 28 48 6 z
rlabel metal1 64 4 64 4 6 vss
rlabel ndcontact 68 16 68 16 6 z
rlabel metal1 60 16 60 16 6 z
rlabel metal1 52 16 52 16 6 z
rlabel metal1 52 24 52 24 6 a
rlabel metal1 68 24 68 24 6 a
rlabel metal1 60 24 60 24 6 a
rlabel metal1 52 36 52 36 6 b
rlabel metal1 68 40 68 40 6 b
rlabel metal1 60 40 60 40 6 b
rlabel metal1 52 48 52 48 6 z
rlabel metal1 68 48 68 48 6 z
rlabel metal1 60 48 60 48 6 z
rlabel metal1 64 68 64 68 6 vdd
rlabel metal1 92 16 92 16 6 z
rlabel metal1 84 16 84 16 6 z
rlabel metal1 100 16 100 16 6 z
rlabel metal1 76 16 76 16 6 z
rlabel metal1 92 24 92 24 6 a
rlabel metal1 84 24 84 24 6 a
rlabel metal1 100 24 100 24 6 a
rlabel metal1 76 28 76 28 6 a
rlabel metal1 76 40 76 40 6 b
rlabel metal1 84 40 84 40 6 b
rlabel metal1 100 40 100 40 6 b
rlabel metal1 92 36 92 36 6 b
rlabel metal1 76 48 76 48 6 z
rlabel metal1 84 48 84 48 6 z
rlabel metal1 92 56 92 56 6 z
rlabel metal1 116 16 116 16 6 z
rlabel metal1 108 16 108 16 6 z
rlabel metal1 108 32 108 32 6 a
<< end >>
