magic
tech scmos
timestamp 1185039025
<< checkpaint >>
rect -22 -24 172 124
<< ab >>
rect 0 0 150 100
<< pwell >>
rect -2 -4 152 49
<< nwell >>
rect -2 49 152 104
<< polysilicon >>
rect 25 95 27 98
rect 37 95 39 98
rect 49 95 51 98
rect 57 95 59 98
rect 69 95 71 98
rect 81 95 83 98
rect 89 95 91 98
rect 113 95 115 98
rect 125 95 127 98
rect 13 69 15 72
rect 13 53 15 55
rect 5 52 15 53
rect 5 48 6 52
rect 10 48 15 52
rect 5 47 15 48
rect 13 37 15 47
rect 25 53 27 75
rect 37 73 39 75
rect 31 72 39 73
rect 31 68 32 72
rect 36 68 39 72
rect 31 67 39 68
rect 25 52 33 53
rect 25 48 28 52
rect 32 48 33 52
rect 25 47 33 48
rect 13 26 15 29
rect 25 23 27 47
rect 37 41 39 67
rect 49 63 51 75
rect 45 62 51 63
rect 45 58 46 62
rect 50 58 51 62
rect 45 57 51 58
rect 47 52 53 53
rect 47 48 48 52
rect 52 51 53 52
rect 57 51 59 75
rect 69 73 71 75
rect 81 73 83 75
rect 52 49 59 51
rect 52 48 53 49
rect 47 47 53 48
rect 37 39 51 41
rect 31 32 39 33
rect 31 28 32 32
rect 36 28 39 32
rect 31 27 39 28
rect 37 23 39 27
rect 49 23 51 39
rect 57 23 59 49
rect 67 71 71 73
rect 77 71 83 73
rect 67 33 69 71
rect 77 53 79 71
rect 89 63 91 75
rect 101 69 103 72
rect 83 62 91 63
rect 83 58 84 62
rect 88 58 91 62
rect 83 57 91 58
rect 137 75 139 78
rect 73 52 79 53
rect 73 48 74 52
rect 78 51 79 52
rect 101 51 103 55
rect 78 49 103 51
rect 78 48 79 49
rect 73 47 79 48
rect 77 39 79 47
rect 63 32 69 33
rect 63 28 64 32
rect 68 28 69 32
rect 63 27 69 28
rect 73 37 79 39
rect 83 42 91 43
rect 83 38 84 42
rect 88 38 91 42
rect 83 37 91 38
rect 101 37 103 49
rect 113 43 115 55
rect 125 43 127 55
rect 137 53 139 55
rect 131 52 139 53
rect 131 48 132 52
rect 136 51 139 52
rect 136 48 137 51
rect 131 47 137 48
rect 141 44 147 45
rect 141 43 142 44
rect 113 41 142 43
rect 73 23 75 37
rect 79 32 85 33
rect 79 28 80 32
rect 84 28 85 32
rect 79 27 85 28
rect 69 21 75 23
rect 69 19 71 21
rect 81 19 83 27
rect 89 19 91 37
rect 101 26 103 29
rect 113 27 115 41
rect 125 27 127 41
rect 141 40 142 41
rect 146 40 147 44
rect 141 39 147 40
rect 131 34 137 35
rect 131 30 132 34
rect 136 31 137 34
rect 136 30 139 31
rect 131 29 139 30
rect 137 27 139 29
rect 25 8 27 11
rect 37 8 39 11
rect 49 8 51 11
rect 57 8 59 11
rect 137 14 139 17
rect 69 4 71 7
rect 81 4 83 7
rect 89 4 91 7
rect 113 4 115 7
rect 125 4 127 7
<< ndiffusion >>
rect 5 29 13 37
rect 15 34 23 37
rect 15 30 18 34
rect 22 30 23 34
rect 15 29 23 30
rect 5 22 11 29
rect 41 32 47 33
rect 41 28 42 32
rect 46 28 47 32
rect 41 23 47 28
rect 5 18 6 22
rect 10 18 11 22
rect 5 17 11 18
rect 17 22 25 23
rect 17 18 18 22
rect 22 18 25 22
rect 17 11 25 18
rect 27 11 37 23
rect 39 11 49 23
rect 51 11 57 23
rect 59 22 67 23
rect 59 18 62 22
rect 66 19 67 22
rect 93 36 101 37
rect 93 32 94 36
rect 98 32 101 36
rect 93 29 101 32
rect 103 29 111 37
rect 105 27 111 29
rect 117 32 123 33
rect 117 28 118 32
rect 122 28 123 32
rect 117 27 123 28
rect 93 22 99 23
rect 93 19 94 22
rect 66 18 69 19
rect 59 11 69 18
rect 61 7 69 11
rect 71 12 81 19
rect 71 8 74 12
rect 78 8 81 12
rect 71 7 81 8
rect 83 7 89 19
rect 91 18 94 19
rect 98 18 99 22
rect 91 7 99 18
rect 105 12 113 27
rect 105 8 106 12
rect 110 8 113 12
rect 105 7 113 8
rect 115 7 125 27
rect 127 17 137 27
rect 139 24 147 27
rect 139 20 142 24
rect 146 20 147 24
rect 139 17 147 20
rect 127 12 135 17
rect 127 8 130 12
rect 134 8 135 12
rect 127 7 135 8
<< pdiffusion >>
rect 5 82 11 83
rect 5 78 6 82
rect 10 78 11 82
rect 5 69 11 78
rect 17 82 25 95
rect 17 78 18 82
rect 22 78 25 82
rect 17 75 25 78
rect 27 75 37 95
rect 39 75 49 95
rect 51 75 57 95
rect 59 82 69 95
rect 59 78 62 82
rect 66 78 69 82
rect 59 75 69 78
rect 71 92 81 95
rect 71 88 74 92
rect 78 88 81 92
rect 71 75 81 88
rect 83 75 89 95
rect 91 82 99 95
rect 91 78 94 82
rect 98 78 99 82
rect 91 75 99 78
rect 105 94 113 95
rect 105 90 106 94
rect 110 90 113 94
rect 5 55 13 69
rect 15 62 23 69
rect 15 58 18 62
rect 22 58 23 62
rect 15 55 23 58
rect 41 72 47 75
rect 41 68 42 72
rect 46 68 47 72
rect 41 67 47 68
rect 105 69 113 90
rect 93 62 101 69
rect 93 58 94 62
rect 98 58 101 62
rect 93 55 101 58
rect 103 55 113 69
rect 115 82 125 95
rect 115 78 118 82
rect 122 78 125 82
rect 115 72 125 78
rect 115 68 118 72
rect 122 68 125 72
rect 115 62 125 68
rect 115 58 118 62
rect 122 58 125 62
rect 115 55 125 58
rect 127 94 135 95
rect 127 90 130 94
rect 134 90 135 94
rect 127 82 135 90
rect 127 78 130 82
rect 134 78 135 82
rect 127 75 135 78
rect 127 72 137 75
rect 127 68 130 72
rect 134 68 137 72
rect 127 62 137 68
rect 127 58 130 62
rect 134 58 137 62
rect 127 55 137 58
rect 139 72 147 75
rect 139 68 142 72
rect 146 68 147 72
rect 139 62 147 68
rect 139 58 142 62
rect 146 58 147 62
rect 139 55 147 58
<< metal1 >>
rect -2 96 152 101
rect -2 94 142 96
rect -2 92 106 94
rect -2 88 74 92
rect 78 90 106 92
rect 110 90 130 94
rect 134 92 142 94
rect 146 92 152 96
rect 134 90 152 92
rect 78 88 152 90
rect -2 87 152 88
rect 5 82 11 87
rect 5 78 6 82
rect 10 78 11 82
rect 5 77 11 78
rect 17 82 67 83
rect 17 78 18 82
rect 22 78 62 82
rect 66 78 67 82
rect 17 77 67 78
rect 93 82 99 83
rect 93 78 94 82
rect 98 78 99 82
rect 93 73 99 78
rect 117 82 123 83
rect 117 78 118 82
rect 122 78 123 82
rect 31 72 37 73
rect 7 68 32 72
rect 36 68 37 72
rect 7 53 13 68
rect 31 67 37 68
rect 41 72 112 73
rect 117 72 123 78
rect 41 68 42 72
rect 46 68 113 72
rect 41 67 113 68
rect 5 52 13 53
rect 5 48 6 52
rect 10 48 13 52
rect 5 47 13 48
rect 7 28 13 47
rect 17 62 51 63
rect 17 58 18 62
rect 22 58 46 62
rect 50 58 51 62
rect 17 57 51 58
rect 17 34 23 57
rect 27 52 33 53
rect 27 48 28 52
rect 32 48 33 52
rect 27 40 33 48
rect 38 52 53 53
rect 38 48 48 52
rect 52 48 53 52
rect 38 47 53 48
rect 57 43 63 67
rect 78 62 89 63
rect 52 42 63 43
rect 17 30 18 34
rect 22 33 23 34
rect 51 38 63 42
rect 67 53 73 62
rect 78 58 84 62
rect 88 58 89 62
rect 78 57 89 58
rect 93 62 102 63
rect 93 58 94 62
rect 98 58 103 62
rect 93 57 103 58
rect 83 53 89 57
rect 67 52 79 53
rect 67 48 74 52
rect 78 48 79 52
rect 67 47 79 48
rect 83 47 92 53
rect 67 38 73 47
rect 83 43 89 47
rect 78 42 89 43
rect 78 38 84 42
rect 88 38 89 42
rect 97 38 103 57
rect 51 37 62 38
rect 78 37 89 38
rect 94 37 103 38
rect 51 33 57 37
rect 93 36 103 37
rect 93 33 94 36
rect 22 32 37 33
rect 22 30 32 32
rect 17 29 32 30
rect 18 28 32 29
rect 36 28 37 32
rect 18 27 37 28
rect 41 32 57 33
rect 41 28 42 32
rect 46 28 57 32
rect 63 32 94 33
rect 98 33 103 36
rect 98 32 102 33
rect 63 28 64 32
rect 68 28 80 32
rect 84 28 99 32
rect 41 27 56 28
rect 63 27 98 28
rect 107 23 113 67
rect 117 68 118 72
rect 122 68 123 72
rect 117 62 123 68
rect 117 58 118 62
rect 122 58 123 62
rect 117 32 123 58
rect 129 82 135 87
rect 129 78 130 82
rect 134 78 135 82
rect 129 72 135 78
rect 129 68 130 72
rect 134 68 135 72
rect 129 62 135 68
rect 129 58 130 62
rect 134 58 135 62
rect 129 57 135 58
rect 141 72 147 73
rect 141 68 142 72
rect 146 68 147 72
rect 141 62 147 68
rect 141 58 142 62
rect 146 58 147 62
rect 117 28 118 32
rect 122 28 123 32
rect 117 27 123 28
rect 131 52 137 53
rect 131 48 132 52
rect 136 48 137 52
rect 131 34 137 48
rect 131 30 132 34
rect 136 30 137 34
rect 131 23 137 30
rect 5 22 11 23
rect 5 18 6 22
rect 10 18 11 22
rect 5 13 11 18
rect 17 22 67 23
rect 17 18 18 22
rect 22 18 62 22
rect 66 18 67 22
rect 17 17 67 18
rect 93 22 137 23
rect 93 18 94 22
rect 98 18 137 22
rect 141 44 147 58
rect 141 40 142 44
rect 146 40 147 44
rect 141 24 147 40
rect 141 20 142 24
rect 146 20 147 24
rect 141 19 147 20
rect 93 17 136 18
rect -2 12 152 13
rect -2 8 74 12
rect 78 8 106 12
rect 110 8 130 12
rect 134 8 152 12
rect -2 -1 152 8
<< ntransistor >>
rect 13 29 15 37
rect 25 11 27 23
rect 37 11 39 23
rect 49 11 51 23
rect 57 11 59 23
rect 101 29 103 37
rect 69 7 71 19
rect 81 7 83 19
rect 89 7 91 19
rect 113 7 115 27
rect 125 7 127 27
rect 137 17 139 27
<< ptransistor >>
rect 25 75 27 95
rect 37 75 39 95
rect 49 75 51 95
rect 57 75 59 95
rect 69 75 71 95
rect 81 75 83 95
rect 89 75 91 95
rect 13 55 15 69
rect 101 55 103 69
rect 113 55 115 95
rect 125 55 127 95
rect 137 55 139 75
<< polycontact >>
rect 6 48 10 52
rect 32 68 36 72
rect 28 48 32 52
rect 46 58 50 62
rect 48 48 52 52
rect 32 28 36 32
rect 84 58 88 62
rect 74 48 78 52
rect 64 28 68 32
rect 84 38 88 42
rect 132 48 136 52
rect 80 28 84 32
rect 142 40 146 44
rect 132 30 136 34
<< ndcontact >>
rect 18 30 22 34
rect 42 28 46 32
rect 6 18 10 22
rect 18 18 22 22
rect 62 18 66 22
rect 94 32 98 36
rect 118 28 122 32
rect 74 8 78 12
rect 94 18 98 22
rect 106 8 110 12
rect 142 20 146 24
rect 130 8 134 12
<< pdcontact >>
rect 6 78 10 82
rect 18 78 22 82
rect 62 78 66 82
rect 74 88 78 92
rect 94 78 98 82
rect 106 90 110 94
rect 18 58 22 62
rect 42 68 46 72
rect 94 58 98 62
rect 118 78 122 82
rect 118 68 122 72
rect 118 58 122 62
rect 130 90 134 94
rect 130 78 134 82
rect 130 68 134 72
rect 130 58 134 62
rect 142 68 146 72
rect 142 58 146 62
<< nsubstratencontact >>
rect 142 92 146 96
<< nsubstratendiff >>
rect 141 96 147 97
rect 141 92 142 96
rect 146 92 147 96
rect 141 85 147 92
<< labels >>
rlabel metal1 10 50 10 50 6 cmd1
rlabel metal1 10 50 10 50 6 cmd1
rlabel polycontact 30 50 30 50 6 i2
rlabel polycontact 30 50 30 50 6 i2
rlabel polycontact 50 50 50 50 6 i1
rlabel polycontact 50 50 50 50 6 i1
rlabel metal1 75 6 75 6 6 vss
rlabel metal1 75 6 75 6 6 vss
rlabel metal1 80 40 80 40 6 i0
rlabel metal1 80 40 80 40 6 i0
rlabel metal1 70 50 70 50 6 cmd0
rlabel metal1 70 50 70 50 6 cmd0
rlabel metal1 80 60 80 60 6 i0
rlabel metal1 80 60 80 60 6 i0
rlabel metal1 75 94 75 94 6 vdd
rlabel metal1 75 94 75 94 6 vdd
rlabel metal1 90 50 90 50 6 i0
rlabel metal1 90 50 90 50 6 i0
rlabel metal1 120 55 120 55 6 nq
rlabel metal1 120 55 120 55 6 nq
<< end >>
