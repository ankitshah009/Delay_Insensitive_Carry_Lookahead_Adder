magic
tech scmos
timestamp 1179387053
<< checkpaint >>
rect -22 -22 174 94
<< ab >>
rect 0 0 152 72
<< pwell >>
rect -4 -4 156 32
<< nwell >>
rect -4 32 156 76
<< polysilicon >>
rect 9 66 11 70
rect 19 66 21 70
rect 29 66 31 70
rect 39 66 41 70
rect 46 66 48 70
rect 56 66 58 70
rect 63 66 65 70
rect 73 66 75 70
rect 80 66 82 70
rect 90 66 92 70
rect 97 66 99 70
rect 107 66 109 70
rect 114 66 116 70
rect 124 58 126 63
rect 131 58 133 63
rect 9 35 11 38
rect 19 35 21 38
rect 29 35 31 38
rect 39 35 41 38
rect 46 35 48 38
rect 56 35 58 38
rect 9 34 31 35
rect 9 33 19 34
rect 9 26 11 33
rect 18 30 19 33
rect 23 30 26 34
rect 30 30 31 34
rect 18 29 31 30
rect 36 34 42 35
rect 36 30 37 34
rect 41 30 42 34
rect 46 33 58 35
rect 63 35 65 38
rect 73 35 75 38
rect 63 34 75 35
rect 63 33 67 34
rect 36 29 42 30
rect 19 26 21 29
rect 29 26 31 29
rect 40 20 42 25
rect 50 24 52 33
rect 66 30 67 33
rect 71 33 75 34
rect 80 35 82 38
rect 90 35 92 38
rect 80 34 92 35
rect 71 30 72 33
rect 66 29 72 30
rect 80 30 81 34
rect 85 33 92 34
rect 97 35 99 38
rect 107 35 109 38
rect 114 35 116 38
rect 124 35 126 38
rect 131 35 133 38
rect 97 34 109 35
rect 85 30 86 33
rect 80 29 86 30
rect 97 30 104 34
rect 108 30 109 34
rect 97 29 109 30
rect 113 34 126 35
rect 113 30 114 34
rect 118 33 126 34
rect 130 34 136 35
rect 118 30 119 33
rect 113 29 119 30
rect 130 30 131 34
rect 135 31 136 34
rect 135 30 142 31
rect 130 29 142 30
rect 60 24 62 29
rect 70 26 72 29
rect 83 26 85 29
rect 93 27 105 29
rect 70 8 72 12
rect 93 24 95 27
rect 103 24 105 27
rect 113 26 115 29
rect 130 26 132 29
rect 140 26 142 29
rect 9 2 11 7
rect 19 2 21 7
rect 29 4 31 7
rect 40 4 42 7
rect 29 2 42 4
rect 50 4 52 7
rect 60 4 62 7
rect 83 4 85 10
rect 130 11 132 16
rect 140 11 142 16
rect 50 2 85 4
rect 93 2 95 6
rect 103 2 105 6
rect 113 2 115 6
<< ndiffusion >>
rect 4 18 9 26
rect 2 17 9 18
rect 2 13 3 17
rect 7 13 9 17
rect 2 12 9 13
rect 4 7 9 12
rect 11 25 19 26
rect 11 21 13 25
rect 17 21 19 25
rect 11 7 19 21
rect 21 17 29 26
rect 21 13 23 17
rect 27 13 29 17
rect 21 7 29 13
rect 31 25 38 26
rect 31 21 33 25
rect 37 21 38 25
rect 31 20 38 21
rect 65 24 70 26
rect 45 20 50 24
rect 31 7 40 20
rect 42 19 50 20
rect 42 15 44 19
rect 48 15 50 19
rect 42 7 50 15
rect 52 12 60 24
rect 52 8 54 12
rect 58 8 60 12
rect 52 7 60 8
rect 62 22 70 24
rect 62 18 64 22
rect 68 18 70 22
rect 62 12 70 18
rect 72 17 83 26
rect 72 13 76 17
rect 80 13 83 17
rect 72 12 83 13
rect 62 7 67 12
rect 78 10 83 12
rect 85 24 90 26
rect 108 24 113 26
rect 85 22 93 24
rect 85 18 87 22
rect 91 18 93 22
rect 85 10 93 18
rect 88 6 93 10
rect 95 11 103 24
rect 95 7 97 11
rect 101 7 103 11
rect 95 6 103 7
rect 105 18 113 24
rect 105 14 107 18
rect 111 14 113 18
rect 105 6 113 14
rect 115 16 130 26
rect 132 22 140 26
rect 132 18 134 22
rect 138 18 140 22
rect 132 16 140 18
rect 142 21 149 26
rect 142 17 144 21
rect 148 17 149 21
rect 142 16 149 17
rect 115 11 128 16
rect 115 7 121 11
rect 125 7 128 11
rect 115 6 128 7
<< pdiffusion >>
rect 4 51 9 66
rect 2 50 9 51
rect 2 46 3 50
rect 7 46 9 50
rect 2 43 9 46
rect 2 39 3 43
rect 7 39 9 43
rect 2 38 9 39
rect 11 65 19 66
rect 11 61 13 65
rect 17 61 19 65
rect 11 58 19 61
rect 11 54 13 58
rect 17 54 19 58
rect 11 38 19 54
rect 21 57 29 66
rect 21 53 23 57
rect 27 53 29 57
rect 21 50 29 53
rect 21 46 23 50
rect 27 46 29 50
rect 21 38 29 46
rect 31 65 39 66
rect 31 61 33 65
rect 37 61 39 65
rect 31 58 39 61
rect 31 54 33 58
rect 37 54 39 58
rect 31 38 39 54
rect 41 38 46 66
rect 48 57 56 66
rect 48 53 50 57
rect 54 53 56 57
rect 48 50 56 53
rect 48 46 50 50
rect 54 46 56 50
rect 48 38 56 46
rect 58 38 63 66
rect 65 65 73 66
rect 65 61 67 65
rect 71 61 73 65
rect 65 58 73 61
rect 65 54 67 58
rect 71 54 73 58
rect 65 38 73 54
rect 75 38 80 66
rect 82 57 90 66
rect 82 53 84 57
rect 88 53 90 57
rect 82 50 90 53
rect 82 46 84 50
rect 88 46 90 50
rect 82 38 90 46
rect 92 38 97 66
rect 99 65 107 66
rect 99 61 101 65
rect 105 61 107 65
rect 99 58 107 61
rect 99 54 101 58
rect 105 54 107 58
rect 99 38 107 54
rect 109 38 114 66
rect 116 58 121 66
rect 116 57 124 58
rect 116 53 118 57
rect 122 53 124 57
rect 116 50 124 53
rect 116 46 118 50
rect 122 46 124 50
rect 116 38 124 46
rect 126 38 131 58
rect 133 57 140 58
rect 133 53 135 57
rect 139 53 140 57
rect 133 50 140 53
rect 133 46 135 50
rect 139 46 140 50
rect 133 38 140 46
<< metal1 >>
rect -2 68 154 72
rect -2 65 142 68
rect -2 64 13 65
rect 12 61 13 64
rect 17 64 33 65
rect 17 61 18 64
rect 12 58 18 61
rect 32 61 33 64
rect 37 64 67 65
rect 37 61 38 64
rect 32 58 38 61
rect 66 61 67 64
rect 71 64 101 65
rect 71 61 72 64
rect 12 54 13 58
rect 17 54 18 58
rect 23 57 27 58
rect 32 54 33 58
rect 37 54 38 58
rect 50 57 54 59
rect 23 50 27 53
rect 66 58 72 61
rect 100 61 101 64
rect 105 64 142 65
rect 146 64 154 68
rect 105 61 106 64
rect 66 54 67 58
rect 71 54 72 58
rect 82 57 88 59
rect 50 50 54 53
rect 82 53 84 57
rect 100 58 106 61
rect 100 54 101 58
rect 105 54 106 58
rect 118 57 123 58
rect 82 50 88 53
rect 122 53 123 57
rect 118 50 123 53
rect 134 57 140 64
rect 134 53 135 57
rect 139 53 140 57
rect 134 50 140 53
rect 2 46 3 50
rect 7 46 23 50
rect 27 46 50 50
rect 54 46 84 50
rect 88 46 118 50
rect 122 46 127 50
rect 134 46 135 50
rect 139 46 140 50
rect 2 43 7 46
rect 2 39 3 43
rect 2 38 7 39
rect 25 38 39 42
rect 68 38 135 42
rect 2 26 6 38
rect 25 34 31 38
rect 68 34 72 38
rect 103 34 109 38
rect 130 34 135 38
rect 17 30 19 34
rect 23 30 26 34
rect 30 30 31 34
rect 36 30 37 34
rect 41 30 67 34
rect 71 30 72 34
rect 80 30 81 34
rect 85 30 99 34
rect 103 30 104 34
rect 108 30 109 34
rect 113 30 114 34
rect 118 30 119 34
rect 95 26 99 30
rect 113 26 119 30
rect 130 30 131 34
rect 130 29 135 30
rect 2 25 39 26
rect 2 21 13 25
rect 17 21 33 25
rect 37 21 39 25
rect 44 22 91 25
rect 95 22 119 26
rect 134 22 138 23
rect 44 21 64 22
rect 44 19 48 21
rect 2 13 3 17
rect 7 13 23 17
rect 27 15 44 17
rect 68 21 87 22
rect 64 17 68 18
rect 27 13 48 15
rect 75 13 76 17
rect 80 13 81 17
rect 87 14 107 18
rect 111 14 138 18
rect 144 21 148 22
rect 54 12 58 13
rect 75 8 81 13
rect 96 8 97 11
rect -2 7 97 8
rect 101 8 102 11
rect 120 8 121 11
rect 101 7 121 8
rect 125 8 126 11
rect 144 8 148 17
rect 125 7 133 8
rect -2 4 133 7
rect 137 4 144 8
rect 148 4 154 8
rect -2 0 154 4
<< ntransistor >>
rect 9 7 11 26
rect 19 7 21 26
rect 29 7 31 26
rect 40 7 42 20
rect 50 7 52 24
rect 60 7 62 24
rect 70 12 72 26
rect 83 10 85 26
rect 93 6 95 24
rect 103 6 105 24
rect 113 6 115 26
rect 130 16 132 26
rect 140 16 142 26
<< ptransistor >>
rect 9 38 11 66
rect 19 38 21 66
rect 29 38 31 66
rect 39 38 41 66
rect 46 38 48 66
rect 56 38 58 66
rect 63 38 65 66
rect 73 38 75 66
rect 80 38 82 66
rect 90 38 92 66
rect 97 38 99 66
rect 107 38 109 66
rect 114 38 116 66
rect 124 38 126 58
rect 131 38 133 58
<< polycontact >>
rect 19 30 23 34
rect 26 30 30 34
rect 37 30 41 34
rect 67 30 71 34
rect 81 30 85 34
rect 104 30 108 34
rect 114 30 118 34
rect 131 30 135 34
<< ndcontact >>
rect 3 13 7 17
rect 13 21 17 25
rect 23 13 27 17
rect 33 21 37 25
rect 44 15 48 19
rect 54 8 58 12
rect 64 18 68 22
rect 76 13 80 17
rect 87 18 91 22
rect 97 7 101 11
rect 107 14 111 18
rect 134 18 138 22
rect 144 17 148 21
rect 121 7 125 11
<< pdcontact >>
rect 3 46 7 50
rect 3 39 7 43
rect 13 61 17 65
rect 13 54 17 58
rect 23 53 27 57
rect 23 46 27 50
rect 33 61 37 65
rect 33 54 37 58
rect 50 53 54 57
rect 50 46 54 50
rect 67 61 71 65
rect 67 54 71 58
rect 84 53 88 57
rect 84 46 88 50
rect 101 61 105 65
rect 101 54 105 58
rect 118 53 122 57
rect 118 46 122 50
rect 135 53 139 57
rect 135 46 139 50
<< psubstratepcontact >>
rect 133 4 137 8
rect 144 4 148 8
<< nsubstratencontact >>
rect 142 64 146 68
<< psubstratepdiff >>
rect 132 8 149 9
rect 132 4 133 8
rect 137 4 144 8
rect 148 4 149 8
rect 132 3 149 4
<< nsubstratendiff >>
rect 139 68 149 69
rect 139 64 142 68
rect 146 64 149 68
rect 139 63 149 64
<< labels >>
rlabel metal1 20 24 20 24 6 z
rlabel metal1 12 24 12 24 6 z
rlabel metal1 4 32 4 32 6 z
rlabel polycontact 20 32 20 32 6 b
rlabel metal1 20 48 20 48 6 z
rlabel metal1 12 48 12 48 6 z
rlabel metal1 46 19 46 19 6 n1
rlabel ndcontact 25 15 25 15 6 n1
rlabel metal1 28 24 28 24 6 z
rlabel ndcontact 36 24 36 24 6 z
rlabel metal1 52 32 52 32 6 a1
rlabel metal1 44 32 44 32 6 a1
rlabel metal1 28 36 28 36 6 b
rlabel metal1 36 40 36 40 6 b
rlabel metal1 28 48 28 48 6 z
rlabel metal1 52 52 52 52 6 z
rlabel metal1 44 48 44 48 6 z
rlabel metal1 36 48 36 48 6 z
rlabel metal1 76 4 76 4 6 vss
rlabel ndcontact 89 19 89 19 6 n1
rlabel metal1 67 23 67 23 6 n1
rlabel polycontact 84 32 84 32 6 a2
rlabel polycontact 68 32 68 32 6 a1
rlabel metal1 60 32 60 32 6 a1
rlabel metal1 84 40 84 40 6 a1
rlabel metal1 76 40 76 40 6 a1
rlabel metal1 60 48 60 48 6 z
rlabel metal1 84 52 84 52 6 z
rlabel metal1 76 48 76 48 6 z
rlabel metal1 68 48 68 48 6 z
rlabel metal1 76 68 76 68 6 vdd
rlabel metal1 108 24 108 24 6 a2
rlabel metal1 100 24 100 24 6 a2
rlabel metal1 116 28 116 28 6 a2
rlabel metal1 92 32 92 32 6 a2
rlabel metal1 92 40 92 40 6 a1
rlabel metal1 116 40 116 40 6 a1
rlabel metal1 108 40 108 40 6 a1
rlabel metal1 100 40 100 40 6 a1
rlabel metal1 92 48 92 48 6 z
rlabel metal1 116 48 116 48 6 z
rlabel metal1 108 48 108 48 6 z
rlabel metal1 100 48 100 48 6 z
rlabel metal1 136 18 136 18 6 n1
rlabel metal1 112 16 112 16 6 n1
rlabel metal1 124 40 124 40 6 a1
rlabel metal1 132 36 132 36 6 a1
rlabel metal1 124 48 124 48 6 z
<< end >>
