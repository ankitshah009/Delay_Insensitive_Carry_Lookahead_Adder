magic
tech scmos
timestamp 1180640197
<< checkpaint >>
rect -24 -26 94 126
<< ab >>
rect 0 0 70 100
<< pwell >>
rect -4 -6 74 49
<< nwell >>
rect -4 49 74 106
<< polysilicon >>
rect 11 83 13 88
rect 23 83 25 88
rect 35 83 37 88
rect 57 83 64 84
rect 57 79 59 83
rect 63 79 64 83
rect 57 78 64 79
rect 57 75 59 78
rect 11 47 13 63
rect 23 54 25 63
rect 35 60 37 63
rect 35 58 47 60
rect 23 53 41 54
rect 23 52 36 53
rect 23 51 27 52
rect 11 46 21 47
rect 11 44 16 46
rect 13 42 16 44
rect 20 42 21 46
rect 13 41 21 42
rect 13 26 15 41
rect 25 31 27 51
rect 35 49 36 52
rect 40 49 41 53
rect 35 48 41 49
rect 45 43 47 58
rect 45 42 51 43
rect 45 38 46 42
rect 50 38 51 42
rect 45 37 51 38
rect 21 29 27 31
rect 21 26 23 29
rect 33 26 35 31
rect 45 26 47 37
rect 57 26 59 55
rect 13 12 15 17
rect 21 12 23 17
rect 33 5 35 17
rect 45 12 47 17
rect 57 5 59 17
rect 33 3 59 5
<< ndiffusion >>
rect 4 22 13 26
rect 4 18 6 22
rect 10 18 13 22
rect 4 17 13 18
rect 15 17 21 26
rect 23 22 33 26
rect 23 18 26 22
rect 30 18 33 22
rect 23 17 33 18
rect 35 22 45 26
rect 35 18 38 22
rect 42 18 45 22
rect 35 17 45 18
rect 47 17 57 26
rect 59 23 64 26
rect 59 22 67 23
rect 59 18 62 22
rect 66 18 67 22
rect 59 17 67 18
rect 49 12 55 17
rect 49 8 50 12
rect 54 8 55 12
rect 49 7 55 8
<< pdiffusion >>
rect 39 92 55 93
rect 39 88 40 92
rect 44 88 50 92
rect 54 88 55 92
rect 39 83 55 88
rect 3 82 11 83
rect 3 78 4 82
rect 8 78 11 82
rect 3 77 11 78
rect 6 63 11 77
rect 13 72 23 83
rect 13 68 16 72
rect 20 68 23 72
rect 13 63 23 68
rect 25 72 35 83
rect 25 68 28 72
rect 32 68 35 72
rect 25 63 35 68
rect 37 82 55 83
rect 37 78 50 82
rect 54 78 55 82
rect 37 75 55 78
rect 37 63 57 75
rect 50 55 57 63
rect 59 61 64 75
rect 59 60 67 61
rect 59 56 62 60
rect 66 56 67 60
rect 59 55 67 56
<< metal1 >>
rect -2 92 72 100
rect -2 88 40 92
rect 44 88 50 92
rect 54 88 72 92
rect 50 82 54 88
rect 3 78 4 82
rect 8 78 40 82
rect 8 72 23 73
rect 8 68 16 72
rect 20 68 23 72
rect 28 72 32 73
rect 8 33 12 68
rect 28 47 32 68
rect 36 53 40 78
rect 50 77 54 78
rect 58 79 59 83
rect 63 79 64 83
rect 58 73 64 79
rect 48 67 64 73
rect 48 57 52 67
rect 62 60 66 61
rect 62 52 66 56
rect 40 49 66 52
rect 36 48 66 49
rect 16 46 32 47
rect 20 42 32 46
rect 16 41 32 42
rect 8 27 22 33
rect 28 32 32 41
rect 37 42 52 43
rect 37 38 46 42
rect 50 38 52 42
rect 28 28 42 32
rect 6 22 10 23
rect 6 12 10 18
rect 18 22 22 27
rect 38 22 42 28
rect 18 18 26 22
rect 30 18 33 22
rect 18 17 33 18
rect 38 17 42 18
rect 48 17 52 38
rect 62 22 66 48
rect 62 17 66 18
rect -2 8 50 12
rect 54 8 72 12
rect -2 0 72 8
<< ntransistor >>
rect 13 17 15 26
rect 21 17 23 26
rect 33 17 35 26
rect 45 17 47 26
rect 57 17 59 26
<< ptransistor >>
rect 11 63 13 83
rect 23 63 25 83
rect 35 63 37 83
rect 57 55 59 75
<< polycontact >>
rect 59 79 63 83
rect 16 42 20 46
rect 36 49 40 53
rect 46 38 50 42
<< ndcontact >>
rect 6 18 10 22
rect 26 18 30 22
rect 38 18 42 22
rect 62 18 66 22
rect 50 8 54 12
<< pdcontact >>
rect 40 88 44 92
rect 50 88 54 92
rect 4 78 8 82
rect 16 68 20 72
rect 28 68 32 72
rect 50 78 54 82
rect 62 56 66 60
<< psubstratepcontact >>
rect 9 4 13 8
rect 18 4 22 8
<< nsubstratencontact >>
rect 8 92 12 96
rect 18 92 22 96
<< psubstratepdiff >>
rect 8 8 23 9
rect 8 4 9 8
rect 13 4 18 8
rect 22 4 23 8
rect 8 3 23 4
<< nsubstratendiff >>
rect 7 96 23 97
rect 7 92 8 96
rect 12 92 18 96
rect 22 92 23 96
rect 7 91 23 92
<< labels >>
rlabel polycontact 38 51 38 51 6 bn
rlabel metal1 10 50 10 50 6 z
rlabel metal1 10 50 10 50 6 z
rlabel metal1 30 20 30 20 6 z
rlabel metal1 30 20 30 20 6 z
rlabel metal1 20 25 20 25 6 z
rlabel metal1 20 25 20 25 6 z
rlabel metal1 24 44 24 44 6 an
rlabel metal1 30 50 30 50 6 an
rlabel metal1 20 70 20 70 6 z
rlabel metal1 20 70 20 70 6 z
rlabel metal1 35 6 35 6 6 vss
rlabel metal1 35 6 35 6 6 vss
rlabel metal1 40 24 40 24 6 an
rlabel metal1 50 30 50 30 6 a
rlabel metal1 40 40 40 40 6 a
rlabel metal1 50 30 50 30 6 a
rlabel metal1 40 40 40 40 6 a
rlabel metal1 50 65 50 65 6 b
rlabel metal1 50 65 50 65 6 b
rlabel metal1 38 65 38 65 6 bn
rlabel metal1 35 94 35 94 6 vdd
rlabel metal1 35 94 35 94 6 vdd
rlabel metal1 21 80 21 80 6 bn
rlabel metal1 64 39 64 39 6 bn
rlabel metal1 60 75 60 75 6 b
rlabel metal1 60 75 60 75 6 b
<< end >>
