magic
tech scmos
timestamp 1180640070
<< checkpaint >>
rect -24 -26 74 126
<< ab >>
rect 0 0 50 100
<< pwell >>
rect -4 -6 54 49
<< nwell >>
rect -4 49 54 106
<< polysilicon >>
rect 13 83 15 88
rect 25 83 27 88
rect 37 83 39 88
rect 13 53 15 71
rect 25 63 27 71
rect 25 62 33 63
rect 25 58 28 62
rect 32 58 33 62
rect 25 57 33 58
rect 13 52 23 53
rect 13 51 18 52
rect 17 48 18 51
rect 22 48 23 52
rect 17 47 23 48
rect 21 39 23 47
rect 29 39 31 57
rect 37 48 39 71
rect 37 47 43 48
rect 37 43 38 47
rect 42 43 43 47
rect 37 42 43 43
rect 37 39 39 42
rect 21 22 23 27
rect 29 22 31 27
rect 37 22 39 27
<< ndiffusion >>
rect 16 33 21 39
rect 13 32 21 33
rect 13 28 14 32
rect 18 28 21 32
rect 13 27 21 28
rect 23 27 29 39
rect 31 27 37 39
rect 39 32 47 39
rect 39 28 42 32
rect 46 28 47 32
rect 39 27 47 28
<< pdiffusion >>
rect 41 92 47 93
rect 41 88 42 92
rect 46 88 47 92
rect 41 83 47 88
rect 8 77 13 83
rect 5 76 13 77
rect 5 72 6 76
rect 10 72 13 76
rect 5 71 13 72
rect 15 82 25 83
rect 15 78 18 82
rect 22 78 25 82
rect 15 71 25 78
rect 27 76 37 83
rect 27 72 30 76
rect 34 72 37 76
rect 27 71 37 72
rect 39 71 47 83
<< metal1 >>
rect -2 92 52 100
rect -2 88 42 92
rect 46 88 52 92
rect 18 82 22 88
rect 18 77 22 78
rect 6 76 12 77
rect 10 72 12 76
rect 30 76 34 77
rect 6 68 34 72
rect 8 32 12 68
rect 38 63 42 83
rect 18 53 22 63
rect 28 62 42 63
rect 32 58 42 62
rect 28 57 42 58
rect 18 52 32 53
rect 22 48 32 52
rect 18 47 32 48
rect 38 47 42 53
rect 18 37 22 47
rect 28 37 42 43
rect 8 28 14 32
rect 18 28 23 32
rect 8 27 23 28
rect 28 27 32 37
rect 42 32 46 33
rect 42 12 46 28
rect -2 0 52 12
<< ntransistor >>
rect 21 27 23 39
rect 29 27 31 39
rect 37 27 39 39
<< ptransistor >>
rect 13 71 15 83
rect 25 71 27 83
rect 37 71 39 83
<< polycontact >>
rect 28 58 32 62
rect 18 48 22 52
rect 38 43 42 47
<< ndcontact >>
rect 14 28 18 32
rect 42 28 46 32
<< pdcontact >>
rect 42 88 46 92
rect 6 72 10 76
rect 18 78 22 82
rect 30 72 34 76
<< psubstratepcontact >>
rect 8 4 12 8
rect 18 4 22 8
<< nsubstratencontact >>
rect 8 92 12 96
rect 18 92 22 96
<< psubstratepdiff >>
rect 7 8 23 9
rect 7 4 8 8
rect 12 4 18 8
rect 22 4 23 8
rect 7 3 23 4
<< nsubstratendiff >>
rect 7 96 23 97
rect 7 92 8 96
rect 12 92 18 96
rect 22 92 23 96
rect 7 91 23 92
<< labels >>
rlabel metal1 10 50 10 50 6 z
rlabel metal1 10 50 10 50 6 z
rlabel metal1 25 6 25 6 6 vss
rlabel metal1 25 6 25 6 6 vss
rlabel metal1 20 30 20 30 6 z
rlabel metal1 20 30 20 30 6 z
rlabel polycontact 20 50 20 50 6 c
rlabel polycontact 20 50 20 50 6 c
rlabel metal1 20 70 20 70 6 z
rlabel metal1 20 70 20 70 6 z
rlabel metal1 25 94 25 94 6 vdd
rlabel metal1 25 94 25 94 6 vdd
rlabel metal1 30 35 30 35 6 a
rlabel metal1 30 35 30 35 6 a
rlabel metal1 30 50 30 50 6 c
rlabel metal1 30 50 30 50 6 c
rlabel polycontact 30 60 30 60 6 b
rlabel polycontact 30 60 30 60 6 b
rlabel metal1 30 70 30 70 6 z
rlabel metal1 30 70 30 70 6 z
rlabel polycontact 40 45 40 45 6 a
rlabel polycontact 40 45 40 45 6 a
rlabel metal1 40 70 40 70 6 b
rlabel metal1 40 70 40 70 6 b
<< end >>
