magic
tech scmos
timestamp 1179385384
<< checkpaint >>
rect -22 -22 166 94
<< ab >>
rect 0 0 144 72
<< pwell >>
rect -4 -4 148 32
<< nwell >>
rect -4 32 148 76
<< polysilicon >>
rect 9 66 11 70
rect 19 66 21 70
rect 29 66 31 70
rect 39 66 41 70
rect 49 66 51 70
rect 59 66 61 70
rect 69 66 71 70
rect 79 66 81 70
rect 89 66 91 70
rect 99 66 101 70
rect 109 66 111 70
rect 119 66 121 70
rect 9 35 11 38
rect 19 35 21 38
rect 29 35 31 38
rect 9 34 31 35
rect 9 30 10 34
rect 14 33 31 34
rect 14 30 21 33
rect 9 29 21 30
rect 19 23 21 29
rect 29 23 31 33
rect 39 35 41 38
rect 49 35 51 38
rect 59 35 61 38
rect 39 34 61 35
rect 39 30 44 34
rect 48 30 56 34
rect 60 30 61 34
rect 39 29 61 30
rect 39 26 41 29
rect 49 26 51 29
rect 59 26 61 29
rect 69 35 71 38
rect 79 35 81 38
rect 89 35 91 38
rect 69 34 91 35
rect 69 30 76 34
rect 80 30 84 34
rect 88 30 91 34
rect 69 29 91 30
rect 69 26 71 29
rect 79 26 81 29
rect 89 26 91 29
rect 99 35 101 38
rect 109 35 111 38
rect 119 35 121 38
rect 99 34 121 35
rect 99 33 109 34
rect 99 26 101 33
rect 108 30 109 33
rect 113 30 116 34
rect 120 30 121 34
rect 108 29 121 30
rect 109 26 111 29
rect 119 26 121 29
rect 19 7 21 12
rect 29 7 31 12
rect 39 3 41 8
rect 49 3 51 8
rect 59 3 61 8
rect 69 3 71 8
rect 79 3 81 8
rect 89 3 91 8
rect 99 3 101 8
rect 109 3 111 8
rect 119 3 121 8
<< ndiffusion >>
rect 34 23 39 26
rect 12 22 19 23
rect 12 18 13 22
rect 17 18 19 22
rect 12 17 19 18
rect 14 12 19 17
rect 21 17 29 23
rect 21 13 23 17
rect 27 13 29 17
rect 21 12 29 13
rect 31 22 39 23
rect 31 18 33 22
rect 37 18 39 22
rect 31 12 39 18
rect 34 8 39 12
rect 41 17 49 26
rect 41 13 43 17
rect 47 13 49 17
rect 41 8 49 13
rect 51 25 59 26
rect 51 21 53 25
rect 57 21 59 25
rect 51 8 59 21
rect 61 24 69 26
rect 61 20 63 24
rect 67 20 69 24
rect 61 17 69 20
rect 61 13 63 17
rect 67 13 69 17
rect 61 8 69 13
rect 71 25 79 26
rect 71 21 73 25
rect 77 21 79 25
rect 71 8 79 21
rect 81 17 89 26
rect 81 13 83 17
rect 87 13 89 17
rect 81 8 89 13
rect 91 25 99 26
rect 91 21 93 25
rect 97 21 99 25
rect 91 18 99 21
rect 91 14 93 18
rect 97 14 99 18
rect 91 8 99 14
rect 101 13 109 26
rect 101 9 103 13
rect 107 9 109 13
rect 101 8 109 9
rect 111 24 119 26
rect 111 20 113 24
rect 117 20 119 24
rect 111 17 119 20
rect 111 13 113 17
rect 117 13 119 17
rect 111 8 119 13
rect 121 21 128 26
rect 121 17 123 21
rect 127 17 128 21
rect 121 13 128 17
rect 121 9 123 13
rect 127 9 128 13
rect 121 8 128 9
<< pdiffusion >>
rect 4 51 9 66
rect 2 50 9 51
rect 2 46 3 50
rect 7 46 9 50
rect 2 43 9 46
rect 2 39 3 43
rect 7 39 9 43
rect 2 38 9 39
rect 11 58 19 66
rect 11 54 13 58
rect 17 54 19 58
rect 11 51 19 54
rect 11 47 13 51
rect 17 47 19 51
rect 11 38 19 47
rect 21 50 29 66
rect 21 46 23 50
rect 27 46 29 50
rect 21 43 29 46
rect 21 39 23 43
rect 27 39 29 43
rect 21 38 29 39
rect 31 58 39 66
rect 31 54 33 58
rect 37 54 39 58
rect 31 51 39 54
rect 31 47 33 51
rect 37 47 39 51
rect 31 38 39 47
rect 41 65 49 66
rect 41 61 43 65
rect 47 61 49 65
rect 41 58 49 61
rect 41 54 43 58
rect 47 54 49 58
rect 41 38 49 54
rect 51 50 59 66
rect 51 46 53 50
rect 57 46 59 50
rect 51 43 59 46
rect 51 39 53 43
rect 57 39 59 43
rect 51 38 59 39
rect 61 65 69 66
rect 61 61 63 65
rect 67 61 69 65
rect 61 58 69 61
rect 61 54 63 58
rect 67 54 69 58
rect 61 38 69 54
rect 71 50 79 66
rect 71 46 73 50
rect 77 46 79 50
rect 71 43 79 46
rect 71 39 73 43
rect 77 39 79 43
rect 71 38 79 39
rect 81 65 89 66
rect 81 61 83 65
rect 87 61 89 65
rect 81 58 89 61
rect 81 54 83 58
rect 87 54 89 58
rect 81 38 89 54
rect 91 50 99 66
rect 91 46 93 50
rect 97 46 99 50
rect 91 43 99 46
rect 91 39 93 43
rect 97 39 99 43
rect 91 38 99 39
rect 101 65 109 66
rect 101 61 103 65
rect 107 61 109 65
rect 101 58 109 61
rect 101 54 103 58
rect 107 54 109 58
rect 101 38 109 54
rect 111 58 119 66
rect 111 54 113 58
rect 117 54 119 58
rect 111 51 119 54
rect 111 47 113 51
rect 117 47 119 51
rect 111 38 119 47
rect 121 65 128 66
rect 121 61 123 65
rect 127 61 128 65
rect 121 58 128 61
rect 121 54 123 58
rect 127 54 128 58
rect 121 38 128 54
<< metal1 >>
rect -2 68 146 72
rect -2 65 133 68
rect -2 64 43 65
rect 42 61 43 64
rect 47 64 63 65
rect 47 61 48 64
rect 2 50 7 59
rect 42 58 48 61
rect 2 46 3 50
rect 12 54 13 58
rect 17 54 33 58
rect 37 54 38 58
rect 42 54 43 58
rect 47 54 48 58
rect 62 61 63 64
rect 67 64 83 65
rect 67 61 68 64
rect 62 58 68 61
rect 62 54 63 58
rect 67 54 68 58
rect 82 61 83 64
rect 87 64 103 65
rect 87 61 88 64
rect 82 58 88 61
rect 82 54 83 58
rect 87 54 88 58
rect 102 61 103 64
rect 107 64 123 65
rect 107 61 108 64
rect 102 58 108 61
rect 122 61 123 64
rect 127 64 133 65
rect 137 64 146 68
rect 127 61 128 64
rect 102 54 103 58
rect 107 54 108 58
rect 113 58 117 59
rect 122 58 128 61
rect 122 54 123 58
rect 127 54 128 58
rect 12 51 18 54
rect 12 47 13 51
rect 17 47 18 51
rect 32 51 38 54
rect 2 43 7 46
rect 2 39 3 43
rect 22 46 23 50
rect 27 46 28 50
rect 32 47 33 51
rect 37 50 38 51
rect 113 51 117 54
rect 37 47 53 50
rect 32 46 53 47
rect 57 46 73 50
rect 77 46 93 50
rect 97 47 113 50
rect 97 46 117 47
rect 22 43 28 46
rect 22 42 23 43
rect 7 39 23 42
rect 27 42 28 43
rect 53 43 57 46
rect 27 39 30 42
rect 2 38 30 39
rect 2 30 10 34
rect 14 30 15 34
rect 2 13 6 30
rect 26 26 30 38
rect 41 34 47 42
rect 53 38 57 39
rect 73 43 77 46
rect 93 43 97 46
rect 73 38 77 39
rect 81 34 87 42
rect 93 38 97 39
rect 122 34 126 51
rect 41 30 44 34
rect 48 30 56 34
rect 60 30 63 34
rect 73 30 76 34
rect 80 30 84 34
rect 88 30 95 34
rect 105 30 109 34
rect 113 30 116 34
rect 120 30 126 34
rect 13 25 58 26
rect 13 22 53 25
rect 37 21 53 22
rect 57 21 58 25
rect 63 24 67 25
rect 37 18 38 21
rect 13 17 17 18
rect 23 17 27 18
rect 33 13 38 18
rect 72 21 73 25
rect 77 21 93 25
rect 97 24 117 25
rect 97 21 113 24
rect 63 17 67 20
rect 93 18 97 21
rect 42 13 43 17
rect 47 13 63 17
rect 67 13 83 17
rect 87 13 88 17
rect 113 17 117 20
rect 93 13 97 14
rect 103 13 107 14
rect 23 8 27 13
rect 113 12 117 13
rect 123 21 127 22
rect 123 13 127 17
rect 103 8 107 9
rect 123 8 127 9
rect -2 4 4 8
rect 8 4 133 8
rect 137 4 146 8
rect -2 0 146 4
<< ntransistor >>
rect 19 12 21 23
rect 29 12 31 23
rect 39 8 41 26
rect 49 8 51 26
rect 59 8 61 26
rect 69 8 71 26
rect 79 8 81 26
rect 89 8 91 26
rect 99 8 101 26
rect 109 8 111 26
rect 119 8 121 26
<< ptransistor >>
rect 9 38 11 66
rect 19 38 21 66
rect 29 38 31 66
rect 39 38 41 66
rect 49 38 51 66
rect 59 38 61 66
rect 69 38 71 66
rect 79 38 81 66
rect 89 38 91 66
rect 99 38 101 66
rect 109 38 111 66
rect 119 38 121 66
<< polycontact >>
rect 10 30 14 34
rect 44 30 48 34
rect 56 30 60 34
rect 76 30 80 34
rect 84 30 88 34
rect 109 30 113 34
rect 116 30 120 34
<< ndcontact >>
rect 13 18 17 22
rect 23 13 27 17
rect 33 18 37 22
rect 43 13 47 17
rect 53 21 57 25
rect 63 20 67 24
rect 63 13 67 17
rect 73 21 77 25
rect 83 13 87 17
rect 93 21 97 25
rect 93 14 97 18
rect 103 9 107 13
rect 113 20 117 24
rect 113 13 117 17
rect 123 17 127 21
rect 123 9 127 13
<< pdcontact >>
rect 3 46 7 50
rect 3 39 7 43
rect 13 54 17 58
rect 13 47 17 51
rect 23 46 27 50
rect 23 39 27 43
rect 33 54 37 58
rect 33 47 37 51
rect 43 61 47 65
rect 43 54 47 58
rect 53 46 57 50
rect 53 39 57 43
rect 63 61 67 65
rect 63 54 67 58
rect 73 46 77 50
rect 73 39 77 43
rect 83 61 87 65
rect 83 54 87 58
rect 93 46 97 50
rect 93 39 97 43
rect 103 61 107 65
rect 103 54 107 58
rect 113 54 117 58
rect 113 47 117 51
rect 123 61 127 65
rect 123 54 127 58
<< psubstratepcontact >>
rect 4 4 8 8
rect 133 4 137 8
<< nsubstratencontact >>
rect 133 64 137 68
<< psubstratepdiff >>
rect 3 8 9 13
rect 3 4 4 8
rect 8 4 9 8
rect 132 8 138 24
rect 3 3 9 4
rect 132 4 133 8
rect 137 4 138 8
rect 132 3 138 4
<< nsubstratendiff >>
rect 132 68 138 69
rect 132 64 133 68
rect 137 64 138 68
rect 132 40 138 64
<< labels >>
rlabel metal1 20 24 20 24 6 z
rlabel metal1 4 20 4 20 6 b
rlabel polycontact 12 32 12 32 6 b
rlabel metal1 12 40 12 40 6 z
rlabel metal1 20 40 20 40 6 z
rlabel metal1 4 52 4 52 6 z
rlabel metal1 15 52 15 52 6 n3
rlabel metal1 44 24 44 24 6 z
rlabel metal1 52 24 52 24 6 z
rlabel ndcontact 36 20 36 20 6 z
rlabel metal1 52 32 52 32 6 a3
rlabel metal1 28 28 28 28 6 z
rlabel metal1 44 36 44 36 6 a3
rlabel metal1 35 52 35 52 6 n3
rlabel metal1 25 56 25 56 6 n3
rlabel metal1 72 4 72 4 6 vss
rlabel metal1 65 19 65 19 6 n2
rlabel metal1 76 32 76 32 6 a2
rlabel metal1 60 32 60 32 6 a3
rlabel metal1 84 36 84 36 6 a2
rlabel metal1 75 44 75 44 6 n3
rlabel metal1 55 44 55 44 6 n3
rlabel metal1 72 68 72 68 6 vdd
rlabel metal1 95 19 95 19 6 n1
rlabel ndcontact 65 15 65 15 6 n2
rlabel metal1 108 32 108 32 6 a1
rlabel metal1 92 32 92 32 6 a2
rlabel metal1 95 44 95 44 6 n3
rlabel metal1 115 18 115 18 6 n1
rlabel ndcontact 94 23 94 23 6 n1
rlabel metal1 116 32 116 32 6 a1
rlabel metal1 124 44 124 44 6 a1
rlabel metal1 115 52 115 52 6 n3
<< end >>
