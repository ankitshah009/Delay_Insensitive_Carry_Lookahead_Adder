magic
tech scmos
timestamp 1179387697
<< checkpaint >>
rect -22 -25 94 105
<< ab >>
rect 0 0 72 80
<< pwell >>
rect -4 -7 76 36
<< nwell >>
rect -4 36 76 87
<< polysilicon >>
rect 29 72 53 74
rect 9 63 11 68
rect 19 63 21 68
rect 29 63 31 72
rect 41 60 43 65
rect 51 63 53 72
rect 51 62 57 63
rect 9 44 11 47
rect 9 43 15 44
rect 9 39 10 43
rect 14 39 15 43
rect 9 38 15 39
rect 19 39 21 47
rect 19 38 25 39
rect 10 28 12 38
rect 19 34 20 38
rect 24 34 25 38
rect 17 32 25 34
rect 17 28 19 32
rect 29 30 31 47
rect 51 58 52 62
rect 56 58 57 62
rect 51 57 57 58
rect 57 46 63 47
rect 41 41 43 44
rect 57 42 58 46
rect 62 42 63 46
rect 57 41 63 42
rect 39 39 63 41
rect 39 30 41 39
rect 49 30 51 35
rect 59 30 61 39
rect 10 12 12 17
rect 17 12 19 17
rect 29 14 31 24
rect 39 18 41 22
rect 49 14 51 22
rect 59 19 61 24
rect 29 12 51 14
<< ndiffusion >>
rect 24 28 29 30
rect 5 23 10 28
rect 3 22 10 23
rect 3 18 4 22
rect 8 18 10 22
rect 3 17 10 18
rect 12 17 17 28
rect 19 24 29 28
rect 31 29 39 30
rect 31 25 33 29
rect 37 25 39 29
rect 31 24 39 25
rect 19 17 27 24
rect 21 12 27 17
rect 34 22 39 24
rect 41 28 49 30
rect 41 24 43 28
rect 47 24 49 28
rect 41 22 49 24
rect 51 29 59 30
rect 51 25 53 29
rect 57 25 59 29
rect 51 24 59 25
rect 61 29 68 30
rect 61 25 63 29
rect 67 25 68 29
rect 61 24 68 25
rect 51 22 56 24
rect 21 8 22 12
rect 26 8 27 12
rect 21 7 27 8
<< pdiffusion >>
rect 33 69 39 70
rect 33 65 34 69
rect 38 65 39 69
rect 33 63 39 65
rect 2 62 9 63
rect 2 58 3 62
rect 7 58 9 62
rect 2 57 9 58
rect 4 47 9 57
rect 11 54 19 63
rect 11 50 13 54
rect 17 50 19 54
rect 11 47 19 50
rect 21 52 29 63
rect 21 48 23 52
rect 27 48 29 52
rect 21 47 29 48
rect 31 60 39 63
rect 31 47 41 60
rect 33 44 41 47
rect 43 50 48 60
rect 43 49 50 50
rect 43 45 45 49
rect 49 45 50 49
rect 43 44 50 45
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect -2 69 74 78
rect -2 68 34 69
rect 33 65 34 68
rect 38 68 74 69
rect 38 65 39 68
rect 2 58 3 62
rect 7 58 37 62
rect 49 58 52 62
rect 56 58 63 62
rect 2 50 13 54
rect 17 50 18 54
rect 23 52 27 53
rect 2 22 6 50
rect 23 46 27 48
rect 11 44 27 46
rect 10 43 27 44
rect 14 42 27 43
rect 14 39 15 42
rect 10 38 15 39
rect 33 38 37 58
rect 57 50 63 58
rect 45 49 49 50
rect 45 38 49 45
rect 57 42 58 46
rect 62 42 70 46
rect 11 30 15 38
rect 19 34 20 38
rect 24 34 57 38
rect 11 29 38 30
rect 53 29 57 34
rect 66 33 70 42
rect 11 26 33 29
rect 32 25 33 26
rect 37 25 38 29
rect 43 28 47 29
rect 53 24 57 25
rect 63 29 67 30
rect 43 22 47 24
rect 2 18 4 22
rect 8 18 47 22
rect 63 12 67 25
rect -2 8 22 12
rect 26 8 74 12
rect -2 2 74 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
<< ntransistor >>
rect 10 17 12 28
rect 17 17 19 28
rect 29 24 31 30
rect 39 22 41 30
rect 49 22 51 30
rect 59 24 61 30
<< ptransistor >>
rect 9 47 11 63
rect 19 47 21 63
rect 29 47 31 63
rect 41 44 43 60
<< polycontact >>
rect 10 39 14 43
rect 20 34 24 38
rect 52 58 56 62
rect 58 42 62 46
<< ndcontact >>
rect 4 18 8 22
rect 33 25 37 29
rect 43 24 47 28
rect 53 25 57 29
rect 63 25 67 29
rect 22 8 26 12
<< pdcontact >>
rect 34 65 38 69
rect 3 58 7 62
rect 13 50 17 54
rect 23 48 27 52
rect 45 45 49 49
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
<< psubstratepdiff >>
rect 0 2 72 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 72 2
rect 0 -3 72 -2
<< nsubstratendiff >>
rect 0 82 72 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 72 82
rect 0 77 72 78
<< labels >>
rlabel polycontact 22 35 22 35 6 an
rlabel polysilicon 11 28 11 28 6 bn
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 20 12 20 6 z
rlabel metal1 20 20 20 20 6 z
rlabel metal1 13 36 13 36 6 bn
rlabel metal1 25 47 25 47 6 bn
rlabel metal1 12 52 12 52 6 z
rlabel metal1 36 6 36 6 6 vss
rlabel metal1 28 20 28 20 6 z
rlabel metal1 24 28 24 28 6 bn
rlabel metal1 36 20 36 20 6 z
rlabel metal1 19 60 19 60 6 an
rlabel metal1 36 74 36 74 6 vdd
rlabel metal1 44 20 44 20 6 z
rlabel metal1 55 31 55 31 6 an
rlabel metal1 38 36 38 36 6 an
rlabel metal1 47 42 47 42 6 an
rlabel metal1 52 60 52 60 6 b
rlabel polycontact 60 44 60 44 6 a
rlabel metal1 68 36 68 36 6 a
rlabel metal1 60 56 60 56 6 b
<< end >>
