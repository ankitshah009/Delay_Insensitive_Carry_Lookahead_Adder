.subckt nts_x2 cmd i nq vdd vss
*   SPICE3 file   created from nts_x2.ext -      technology: scmos
m00 w1     i      vdd    vdd p w=39u  l=2.3636u ad=195p     pd=49.6364u as=388.408p ps=82.7755u
m01 nq     w2     w1     vdd p w=38u  l=2.3636u ad=190p     pd=48u      as=190p     ps=48.3636u
m02 w3     w2     nq     vdd p w=38u  l=2.3636u ad=190p     pd=48.3636u as=190p     ps=48u
m03 vdd    i      w3     vdd p w=39u  l=2.3636u ad=388.408p pd=82.7755u as=195p     ps=49.6364u
m04 w2     cmd    vdd    vdd p w=20u  l=2.3636u ad=160p     pd=56u      as=199.184p ps=42.449u
m05 w4     i      vss    vss n w=19u  l=2.3636u ad=95p      pd=29.7838u as=188.417p ps=50.6667u
m06 nq     cmd    w4     vss n w=18u  l=2.3636u ad=90p      pd=28u      as=90p      ps=28.2162u
m07 w5     cmd    nq     vss n w=18u  l=2.3636u ad=90p      pd=28.2162u as=90p      ps=28u
m08 vss    i      w5     vss n w=19u  l=2.3636u ad=188.417p pd=50.6667u as=95p      ps=29.7838u
m09 w2     cmd    vss    vss n w=10u  l=2.3636u ad=80p      pd=36u      as=99.1667p ps=26.6667u
C0  vdd    w2     0.262f
C1  w1     i      0.055f
C2  w2     i      0.171f
C3  cmd    nq     0.090f
C4  w4     i      0.016f
C5  cmd    vdd    0.045f
C6  vss    w2     0.028f
C7  cmd    i      0.195f
C8  nq     vdd    0.083f
C9  w3     w2     0.061f
C10 w4     vss    0.019f
C11 nq     i      0.339f
C12 vss    cmd    0.094f
C13 vdd    i      0.113f
C14 vss    nq     0.052f
C15 vss    vdd    0.004f
C16 vss    i      0.052f
C17 w3     vdd    0.019f
C18 cmd    w2     0.278f
C19 w5     vss    0.019f
C20 nq     w2     0.229f
C21 w1     vdd    0.019f
C23 cmd    vss    0.066f
C24 nq     vss    0.013f
C26 w2     vss    0.042f
C27 i      vss    0.064f
.ends
