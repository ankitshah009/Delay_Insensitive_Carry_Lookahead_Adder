magic
tech scmos
timestamp 1179387239
<< checkpaint >>
rect -22 -25 102 105
<< ab >>
rect 0 0 80 80
<< pwell >>
rect -4 -7 84 36
<< nwell >>
rect -4 36 84 87
<< polysilicon >>
rect 31 70 33 74
rect 38 70 40 74
rect 45 70 47 74
rect 55 70 57 74
rect 62 70 64 74
rect 69 70 71 74
rect 9 61 11 65
rect 19 63 21 68
rect 9 39 11 42
rect 19 39 21 42
rect 31 39 33 42
rect 9 38 21 39
rect 9 34 16 38
rect 20 34 21 38
rect 9 33 21 34
rect 28 38 34 39
rect 28 34 29 38
rect 33 34 34 38
rect 28 33 34 34
rect 9 30 11 33
rect 29 22 31 33
rect 38 31 40 42
rect 45 39 47 42
rect 55 39 57 42
rect 45 38 57 39
rect 45 37 52 38
rect 51 34 52 37
rect 56 34 57 38
rect 51 33 57 34
rect 38 30 47 31
rect 38 26 42 30
rect 46 26 47 30
rect 38 25 47 26
rect 39 22 41 25
rect 52 22 54 33
rect 62 31 64 42
rect 69 39 71 42
rect 69 38 78 39
rect 69 37 73 38
rect 72 34 73 37
rect 77 34 78 38
rect 72 33 78 34
rect 62 30 68 31
rect 62 26 63 30
rect 67 26 68 30
rect 62 25 68 26
rect 9 6 11 10
rect 29 7 31 12
rect 39 7 41 12
rect 52 7 54 12
<< ndiffusion >>
rect 2 29 9 30
rect 2 25 3 29
rect 7 25 9 29
rect 2 22 9 25
rect 2 18 3 22
rect 7 18 9 22
rect 2 17 9 18
rect 4 10 9 17
rect 11 23 27 30
rect 11 19 13 23
rect 17 22 27 23
rect 17 19 29 22
rect 11 17 29 19
rect 11 15 23 17
rect 11 11 13 15
rect 17 13 23 15
rect 27 13 29 17
rect 17 12 29 13
rect 31 21 39 22
rect 31 17 33 21
rect 37 17 39 21
rect 31 12 39 17
rect 41 12 52 22
rect 54 21 61 22
rect 54 17 56 21
rect 60 17 61 21
rect 54 16 61 17
rect 54 12 59 16
rect 17 11 27 12
rect 11 10 27 11
rect 43 8 44 12
rect 48 8 50 12
rect 43 7 50 8
<< pdiffusion >>
rect 23 69 31 70
rect 23 65 24 69
rect 28 65 31 69
rect 23 63 31 65
rect 14 61 19 63
rect 2 60 9 61
rect 2 56 3 60
rect 7 56 9 60
rect 2 53 9 56
rect 2 49 3 53
rect 7 49 9 53
rect 2 42 9 49
rect 11 54 19 61
rect 11 50 13 54
rect 17 50 19 54
rect 11 47 19 50
rect 11 43 13 47
rect 17 43 19 47
rect 11 42 19 43
rect 21 62 31 63
rect 21 58 24 62
rect 28 58 31 62
rect 21 42 31 58
rect 33 42 38 70
rect 40 42 45 70
rect 47 62 55 70
rect 47 58 49 62
rect 53 58 55 62
rect 47 55 55 58
rect 47 51 49 55
rect 53 51 55 55
rect 47 42 55 51
rect 57 42 62 70
rect 64 42 69 70
rect 71 69 78 70
rect 71 65 73 69
rect 77 65 78 69
rect 71 61 78 65
rect 71 57 73 61
rect 77 57 78 61
rect 71 42 78 57
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect -2 69 82 78
rect -2 68 24 69
rect 2 60 8 68
rect 2 56 3 60
rect 7 56 8 60
rect 23 65 24 68
rect 28 68 73 69
rect 28 65 29 68
rect 23 62 29 65
rect 77 68 82 69
rect 23 58 24 62
rect 28 58 29 62
rect 49 62 53 63
rect 2 53 8 56
rect 49 55 53 58
rect 73 61 77 65
rect 73 56 77 57
rect 2 49 3 53
rect 7 49 8 53
rect 13 54 17 55
rect 13 47 17 50
rect 2 43 13 46
rect 2 42 17 43
rect 21 51 49 54
rect 21 50 53 51
rect 2 30 6 42
rect 21 38 25 50
rect 58 46 62 55
rect 33 42 78 46
rect 15 34 16 38
rect 20 34 25 38
rect 28 34 29 38
rect 33 34 39 42
rect 72 38 78 42
rect 49 34 52 38
rect 56 34 63 38
rect 72 34 73 38
rect 77 34 78 38
rect 2 29 7 30
rect 2 25 3 29
rect 21 29 25 34
rect 74 33 78 34
rect 21 25 36 29
rect 41 26 42 30
rect 46 26 63 30
rect 67 26 70 30
rect 2 22 7 25
rect 2 18 3 22
rect 2 17 7 18
rect 13 23 17 24
rect 13 15 17 19
rect 32 21 36 25
rect -2 11 13 12
rect 23 17 27 18
rect 32 17 33 21
rect 37 17 56 21
rect 60 17 61 21
rect 66 17 70 26
rect 23 12 27 13
rect 17 11 44 12
rect -2 8 44 11
rect 48 8 82 12
rect -2 2 82 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
<< ntransistor >>
rect 9 10 11 30
rect 29 12 31 22
rect 39 12 41 22
rect 52 12 54 22
<< ptransistor >>
rect 9 42 11 61
rect 19 42 21 63
rect 31 42 33 70
rect 38 42 40 70
rect 45 42 47 70
rect 55 42 57 70
rect 62 42 64 70
rect 69 42 71 70
<< polycontact >>
rect 16 34 20 38
rect 29 34 33 38
rect 52 34 56 38
rect 42 26 46 30
rect 73 34 77 38
rect 63 26 67 30
<< ndcontact >>
rect 3 25 7 29
rect 3 18 7 22
rect 13 19 17 23
rect 13 11 17 15
rect 23 13 27 17
rect 33 17 37 21
rect 56 17 60 21
rect 44 8 48 12
<< pdcontact >>
rect 24 65 28 69
rect 3 56 7 60
rect 3 49 7 53
rect 13 50 17 54
rect 13 43 17 47
rect 24 58 28 62
rect 49 58 53 62
rect 49 51 53 55
rect 73 65 77 69
rect 73 57 77 61
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
<< psubstratepdiff >>
rect 0 2 80 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 80 2
rect 0 -3 80 -2
<< nsubstratendiff >>
rect 0 82 80 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 80 82
rect 0 77 80 78
<< labels >>
rlabel polysilicon 15 36 15 36 6 zn
rlabel ndcontact 4 28 4 28 6 z
rlabel metal1 12 44 12 44 6 z
rlabel metal1 20 36 20 36 6 zn
rlabel metal1 40 6 40 6 6 vss
rlabel polycontact 44 28 44 28 6 b
rlabel metal1 44 44 44 44 6 a
rlabel metal1 36 40 36 40 6 a
rlabel metal1 40 74 40 74 6 vdd
rlabel metal1 52 28 52 28 6 b
rlabel metal1 46 19 46 19 6 zn
rlabel metal1 60 28 60 28 6 b
rlabel metal1 52 36 52 36 6 c
rlabel metal1 52 44 52 44 6 a
rlabel metal1 60 36 60 36 6 c
rlabel metal1 60 48 60 48 6 a
rlabel metal1 51 56 51 56 6 zn
rlabel metal1 68 20 68 20 6 b
rlabel metal1 68 44 68 44 6 a
rlabel polycontact 76 36 76 36 6 a
<< end >>
