magic
tech scmos
timestamp 1179387018
<< checkpaint >>
rect -22 -25 62 105
<< ab >>
rect 0 0 40 80
<< pwell >>
rect -4 -7 44 36
<< nwell >>
rect -4 36 44 87
<< polysilicon >>
rect 12 70 14 74
rect 22 70 24 74
rect 29 70 31 74
rect 12 50 14 56
rect 9 49 15 50
rect 9 45 10 49
rect 14 45 15 49
rect 9 44 15 45
rect 9 22 11 44
rect 22 40 24 43
rect 17 39 24 40
rect 17 35 18 39
rect 22 35 24 39
rect 17 34 24 35
rect 29 39 31 43
rect 29 38 38 39
rect 29 34 33 38
rect 37 34 38 38
rect 19 22 21 34
rect 29 33 38 34
rect 29 22 31 33
rect 9 6 11 10
rect 19 6 21 10
rect 29 6 31 10
<< ndiffusion >>
rect 2 21 9 22
rect 2 17 3 21
rect 7 17 9 21
rect 2 16 9 17
rect 4 10 9 16
rect 11 21 19 22
rect 11 17 13 21
rect 17 17 19 21
rect 11 10 19 17
rect 21 15 29 22
rect 21 11 23 15
rect 27 11 29 15
rect 21 10 29 11
rect 31 21 38 22
rect 31 17 33 21
rect 37 17 38 21
rect 31 16 38 17
rect 31 10 36 16
<< pdiffusion >>
rect 4 69 12 70
rect 4 65 6 69
rect 10 65 12 69
rect 4 56 12 65
rect 14 62 22 70
rect 14 58 16 62
rect 20 58 22 62
rect 14 56 22 58
rect 17 43 22 56
rect 24 43 29 70
rect 31 69 38 70
rect 31 65 33 69
rect 37 65 38 69
rect 31 62 38 65
rect 31 58 33 62
rect 37 58 38 62
rect 31 43 38 58
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect -2 69 42 78
rect -2 68 6 69
rect 5 65 6 68
rect 10 68 33 69
rect 10 65 11 68
rect 32 65 33 68
rect 37 68 42 69
rect 37 65 38 68
rect 32 62 38 65
rect 2 58 16 62
rect 20 58 23 62
rect 32 58 33 62
rect 37 58 38 62
rect 2 22 6 58
rect 10 49 14 50
rect 25 47 31 54
rect 10 30 14 45
rect 18 42 31 47
rect 18 39 22 42
rect 18 34 22 35
rect 25 34 33 38
rect 37 34 38 38
rect 10 26 23 30
rect 34 25 38 34
rect 2 21 8 22
rect 2 17 3 21
rect 7 17 8 21
rect 12 21 38 22
rect 12 17 13 21
rect 17 18 33 21
rect 17 17 18 18
rect 32 17 33 18
rect 37 17 38 21
rect 22 12 23 15
rect -2 11 23 12
rect 27 12 28 15
rect 27 11 42 12
rect -2 2 42 11
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
<< ntransistor >>
rect 9 10 11 22
rect 19 10 21 22
rect 29 10 31 22
<< ptransistor >>
rect 12 56 14 70
rect 22 43 24 70
rect 29 43 31 70
<< polycontact >>
rect 10 45 14 49
rect 18 35 22 39
rect 33 34 37 38
<< ndcontact >>
rect 3 17 7 21
rect 13 17 17 21
rect 23 11 27 15
rect 33 17 37 21
<< pdcontact >>
rect 6 65 10 69
rect 16 58 20 62
rect 33 65 37 69
rect 33 58 37 62
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
<< psubstratepdiff >>
rect 0 2 40 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 40 2
rect 0 -3 40 -2
<< nsubstratendiff >>
rect 0 82 40 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 40 82
rect 0 77 40 78
<< labels >>
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 40 12 40 6 b
rlabel metal1 12 60 12 60 6 z
rlabel metal1 20 6 20 6 6 vss
rlabel metal1 20 28 20 28 6 b
rlabel metal1 28 36 28 36 6 a1
rlabel metal1 20 44 20 44 6 a2
rlabel metal1 28 48 28 48 6 a2
rlabel metal1 20 60 20 60 6 z
rlabel metal1 20 74 20 74 6 vdd
rlabel metal1 25 20 25 20 6 n1
rlabel metal1 36 28 36 28 6 a1
<< end >>
