magic
tech scmos
timestamp 1170759777
<< checkpaint >>
rect -22 -26 54 114
<< ab >>
rect 0 0 32 88
<< pwell >>
rect -4 -8 36 40
<< nwell >>
rect -4 40 36 96
<< polysilicon >>
rect 2 82 11 83
rect 2 78 6 82
rect 10 78 11 82
rect 2 77 11 78
rect 9 74 11 77
rect 21 82 30 83
rect 21 78 23 82
rect 27 78 30 82
rect 21 77 30 78
rect 21 74 23 77
rect 9 43 11 46
rect 21 43 23 46
rect 2 37 14 43
rect 18 37 30 43
rect 9 34 11 37
rect 21 34 23 37
rect 9 11 11 14
rect 2 5 11 11
rect 21 11 23 14
rect 21 5 30 11
<< ndiffusion >>
rect 2 14 9 34
rect 11 26 21 34
rect 11 22 14 26
rect 18 22 21 26
rect 11 19 21 22
rect 11 15 14 19
rect 18 15 21 19
rect 11 14 21 15
rect 23 33 30 34
rect 23 29 25 33
rect 29 29 30 33
rect 23 26 30 29
rect 23 22 25 26
rect 29 22 30 26
rect 23 14 30 22
rect 13 2 19 14
<< pdiffusion >>
rect 13 75 19 86
rect 13 74 14 75
rect 2 46 9 74
rect 11 71 14 74
rect 18 74 19 75
rect 18 71 21 74
rect 11 46 21 71
rect 23 58 30 74
rect 23 54 25 58
rect 29 54 30 58
rect 23 51 30 54
rect 23 47 25 51
rect 29 47 30 51
rect 23 46 30 47
<< metal1 >>
rect -2 86 2 90
rect 10 86 22 90
rect 30 86 34 90
rect 6 82 10 86
rect 6 77 10 78
rect 14 82 18 86
rect 14 75 18 78
rect 14 70 18 71
rect 22 78 23 82
rect 27 78 28 82
rect 22 66 28 78
rect 14 62 28 66
rect 14 41 18 62
rect 24 55 25 58
rect 22 54 25 55
rect 29 54 30 58
rect 22 51 30 54
rect 22 47 25 51
rect 29 47 30 51
rect 22 33 26 47
rect 22 29 25 33
rect 29 29 30 33
rect 14 26 18 27
rect 14 19 18 22
rect 22 26 30 29
rect 22 22 25 26
rect 29 22 30 26
rect 22 17 26 22
rect 14 10 18 15
rect 14 2 18 6
rect -2 -2 2 2
rect 10 -2 22 2
rect 30 -2 34 2
<< metal2 >>
rect -2 86 6 90
rect 10 86 22 90
rect 26 86 34 90
rect -2 82 34 86
rect -2 78 14 82
rect 18 78 34 82
rect -2 76 34 78
rect -2 10 34 12
rect -2 6 14 10
rect 18 6 34 10
rect -2 2 34 6
rect -2 -2 6 2
rect 10 -2 22 2
rect 26 -2 34 2
<< ntransistor >>
rect 9 14 11 34
rect 21 14 23 34
<< ptransistor >>
rect 9 46 11 74
rect 21 46 23 74
<< polycontact >>
rect 6 78 10 82
rect 23 78 27 82
<< ndcontact >>
rect 14 22 18 26
rect 14 15 18 19
rect 25 29 29 33
rect 25 22 29 26
<< pdcontact >>
rect 14 71 18 75
rect 25 54 29 58
rect 25 47 29 51
<< m2contact >>
rect 6 86 10 90
rect 22 86 26 90
rect 14 78 18 82
rect 14 6 18 10
rect 6 -2 10 2
rect 22 -2 26 2
<< psubstratepcontact >>
rect 2 -2 6 2
rect 26 -2 30 2
<< nsubstratencontact >>
rect 2 86 6 90
rect 26 86 30 90
<< psubstratepdiff >>
rect 0 2 7 3
rect 25 2 32 3
rect 0 -2 2 2
rect 6 -2 7 2
rect 0 -3 7 -2
rect 25 -2 26 2
rect 30 -2 32 2
rect 25 -3 32 -2
<< nsubstratendiff >>
rect 0 90 7 91
rect 0 86 2 90
rect 6 86 7 90
rect 25 90 32 91
rect 25 86 26 90
rect 30 86 32 90
rect 0 85 7 86
rect 25 85 32 86
<< labels >>
rlabel metal1 16 52 16 52 6 a
rlabel metal1 24 36 24 36 6 z
rlabel metal1 24 68 24 68 6 a
rlabel metal2 16 6 16 6 6 vss
rlabel metal2 16 6 16 6 6 vss
rlabel metal2 16 82 16 82 6 vdd
<< end >>
