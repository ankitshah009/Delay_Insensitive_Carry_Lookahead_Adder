magic
tech scmos
timestamp 1179386345
<< checkpaint >>
rect -22 -22 54 94
<< ab >>
rect 0 0 32 72
<< pwell >>
rect -4 -4 36 32
<< nwell >>
rect -4 32 36 76
<< polysilicon >>
rect 10 56 16 57
rect 10 52 11 56
rect 15 52 16 56
rect 10 51 16 52
rect 10 48 12 51
rect 20 48 22 53
rect 10 35 12 38
rect 20 35 22 38
rect 9 32 12 35
rect 16 34 23 35
rect 9 26 11 32
rect 16 30 18 34
rect 22 30 23 34
rect 16 29 23 30
rect 16 26 18 29
rect 9 4 11 9
rect 16 4 18 9
<< ndiffusion >>
rect 2 25 9 26
rect 2 21 3 25
rect 7 21 9 25
rect 2 18 9 21
rect 2 14 3 18
rect 7 14 9 18
rect 2 13 9 14
rect 4 9 9 13
rect 11 9 16 26
rect 18 14 26 26
rect 18 10 20 14
rect 24 10 26 14
rect 18 9 26 10
<< pdiffusion >>
rect 2 66 8 67
rect 2 62 3 66
rect 7 62 8 66
rect 2 48 8 62
rect 24 50 30 51
rect 24 48 25 50
rect 2 38 10 48
rect 12 43 20 48
rect 12 39 14 43
rect 18 39 20 43
rect 12 38 20 39
rect 22 46 25 48
rect 29 46 30 50
rect 22 38 30 46
<< metal1 >>
rect -2 68 34 72
rect -2 66 16 68
rect -2 64 3 66
rect 2 62 3 64
rect 7 64 16 66
rect 20 64 24 68
rect 28 64 34 68
rect 7 62 8 64
rect 9 56 23 58
rect 9 52 11 56
rect 15 54 23 56
rect 9 46 15 52
rect 26 50 30 64
rect 24 46 25 50
rect 29 46 30 50
rect 13 42 14 43
rect 2 39 14 42
rect 18 39 19 43
rect 2 38 19 39
rect 2 26 6 38
rect 17 30 18 34
rect 22 30 23 34
rect 17 27 23 30
rect 2 25 7 26
rect 2 21 3 25
rect 17 21 30 27
rect 2 18 7 21
rect 2 14 3 18
rect 2 13 7 14
rect 20 14 24 15
rect 20 8 24 10
rect -2 0 34 8
<< ntransistor >>
rect 9 9 11 26
rect 16 9 18 26
<< ptransistor >>
rect 10 38 12 48
rect 20 38 22 48
<< polycontact >>
rect 11 52 15 56
rect 18 30 22 34
<< ndcontact >>
rect 3 21 7 25
rect 3 14 7 18
rect 20 10 24 14
<< pdcontact >>
rect 3 62 7 66
rect 14 39 18 43
rect 25 46 29 50
<< nsubstratencontact >>
rect 16 64 20 68
rect 24 64 28 68
<< nsubstratendiff >>
rect 15 68 29 69
rect 15 64 16 68
rect 20 64 24 68
rect 28 64 29 68
rect 15 63 29 64
<< labels >>
rlabel ndcontact 4 24 4 24 6 z
rlabel metal1 12 40 12 40 6 z
rlabel metal1 12 52 12 52 6 b
rlabel metal1 16 4 16 4 6 vss
rlabel metal1 20 28 20 28 6 a
rlabel metal1 20 56 20 56 6 b
rlabel metal1 16 68 16 68 6 vdd
rlabel metal1 28 24 28 24 6 a
<< end >>
