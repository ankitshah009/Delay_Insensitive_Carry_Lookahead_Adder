magic
tech scmos
timestamp 1179386445
<< checkpaint >>
rect -22 -25 54 105
<< ab >>
rect 0 0 32 80
<< pwell >>
rect -4 -7 36 36
<< nwell >>
rect -4 36 36 87
<< polysilicon >>
rect 10 62 16 63
rect 10 58 11 62
rect 15 58 16 62
rect 10 57 16 58
rect 10 54 12 57
rect 20 54 22 59
rect 10 39 12 42
rect 20 39 22 42
rect 9 36 12 39
rect 16 38 23 39
rect 9 30 11 36
rect 16 34 18 38
rect 22 34 23 38
rect 16 33 23 34
rect 16 30 18 33
rect 9 17 11 22
rect 16 17 18 22
<< ndiffusion >>
rect 2 29 9 30
rect 2 25 3 29
rect 7 25 9 29
rect 2 24 9 25
rect 4 22 9 24
rect 11 22 16 30
rect 18 22 27 30
rect 20 18 21 22
rect 25 18 27 22
rect 20 17 27 18
<< pdiffusion >>
rect 2 70 8 71
rect 2 66 3 70
rect 7 66 8 70
rect 2 54 8 66
rect 2 42 10 54
rect 12 47 20 54
rect 12 43 14 47
rect 18 43 20 47
rect 12 42 20 43
rect 22 53 30 54
rect 22 49 25 53
rect 29 49 30 53
rect 22 42 30 49
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect -2 70 34 78
rect -2 68 3 70
rect 2 66 3 68
rect 7 68 34 70
rect 7 66 8 68
rect 9 58 11 62
rect 15 58 23 62
rect 9 50 15 58
rect 26 53 30 68
rect 24 49 25 53
rect 29 49 30 53
rect 13 46 14 47
rect 2 43 14 46
rect 18 43 19 47
rect 2 42 19 43
rect 2 30 6 42
rect 17 34 18 38
rect 22 34 23 38
rect 17 31 23 34
rect 2 29 7 30
rect 2 25 3 29
rect 17 25 30 31
rect 2 24 7 25
rect 20 18 21 22
rect 25 18 26 22
rect 20 12 26 18
rect -2 2 34 12
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
<< ntransistor >>
rect 9 22 11 30
rect 16 22 18 30
<< ptransistor >>
rect 10 42 12 54
rect 20 42 22 54
<< polycontact >>
rect 11 58 15 62
rect 18 34 22 38
<< ndcontact >>
rect 3 25 7 29
rect 21 18 25 22
<< pdcontact >>
rect 3 66 7 70
rect 14 43 18 47
rect 25 49 29 53
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
<< psubstratepdiff >>
rect 0 2 32 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 32 2
rect 0 -3 32 -2
<< nsubstratendiff >>
rect 0 82 32 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 32 82
rect 0 77 32 78
<< labels >>
rlabel metal1 4 32 4 32 6 z
rlabel metal1 12 44 12 44 6 z
rlabel metal1 12 56 12 56 6 b
rlabel metal1 16 6 16 6 6 vss
rlabel metal1 20 32 20 32 6 a
rlabel metal1 20 60 20 60 6 b
rlabel metal1 16 74 16 74 6 vdd
rlabel metal1 28 28 28 28 6 a
<< end >>
