.subckt nr2av1x05 a b vdd vss z
*   SPICE3 file   created from nr2av1x05.ext -      technology: scmos
m00 w1     b      z      vdd p w=15u  l=2.3636u ad=37.5p    pd=20u      as=87p      ps=44u
m01 vdd    an     w1     vdd p w=15u  l=2.3636u ad=96.6667p pd=30u      as=37.5p    ps=20u
m02 an     a      vdd    vdd p w=12u  l=2.3636u ad=72p      pd=38u      as=77.3333p ps=24u
m03 an     a      vss    vss n w=6u   l=2.3636u ad=42p      pd=26u      as=62.7273p ps=26.7273u
m04 z      b      vss    vss n w=8u   l=2.3636u ad=32p      pd=16u      as=83.6364p ps=35.6364u
m05 vss    an     z      vss n w=8u   l=2.3636u ad=83.6364p pd=35.6364u as=32p      ps=16u
C0  w1     b      0.006f
C1  z      an     0.088f
C2  a      vdd    0.039f
C3  an     b      0.171f
C4  z      vdd    0.097f
C5  b      vdd    0.059f
C6  a      z      0.041f
C7  vss    an     0.084f
C8  vss    vdd    0.006f
C9  a      b      0.140f
C10 z      b      0.173f
C11 an     vdd    0.049f
C12 vss    a      0.022f
C13 vss    z      0.184f
C14 w1     z      0.003f
C15 a      an     0.241f
C16 vss    b      0.017f
C18 a      vss    0.030f
C19 z      vss    0.020f
C20 an     vss    0.030f
C21 b      vss    0.025f
.ends
