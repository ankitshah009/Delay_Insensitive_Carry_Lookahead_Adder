magic
tech scmos
timestamp 1180600683
<< checkpaint >>
rect -22 -22 102 122
<< ab >>
rect 0 0 80 100
<< pwell >>
rect -4 -4 84 48
<< nwell >>
rect -4 48 84 104
<< polysilicon >>
rect 45 94 47 98
rect 57 94 59 98
rect 11 83 13 87
rect 23 83 25 87
rect 35 83 37 87
rect 11 43 13 63
rect 23 53 25 63
rect 17 52 25 53
rect 17 48 18 52
rect 22 48 25 52
rect 17 47 25 48
rect 7 42 15 43
rect 7 38 8 42
rect 12 38 15 42
rect 7 37 15 38
rect 13 34 15 37
rect 21 34 23 47
rect 35 43 37 63
rect 67 83 73 84
rect 67 79 68 83
rect 72 79 73 83
rect 67 78 73 79
rect 67 75 69 78
rect 45 43 47 55
rect 57 43 59 55
rect 27 42 37 43
rect 27 38 28 42
rect 32 41 37 42
rect 43 42 63 43
rect 32 38 33 41
rect 27 37 33 38
rect 43 38 58 42
rect 62 38 63 42
rect 43 37 63 38
rect 29 34 31 37
rect 43 25 45 37
rect 55 25 57 37
rect 67 25 69 55
rect 13 11 15 15
rect 21 11 23 15
rect 29 11 31 15
rect 67 11 69 15
rect 43 2 45 6
rect 55 2 57 6
<< ndiffusion >>
rect 5 22 13 34
rect 5 18 6 22
rect 10 18 13 22
rect 5 15 13 18
rect 15 15 21 34
rect 23 15 29 34
rect 31 25 41 34
rect 31 15 43 25
rect 33 12 43 15
rect 33 8 36 12
rect 40 8 43 12
rect 33 6 43 8
rect 45 22 55 25
rect 45 18 48 22
rect 52 18 55 22
rect 45 6 55 18
rect 57 15 67 25
rect 69 22 77 25
rect 69 18 72 22
rect 76 18 77 22
rect 69 15 77 18
rect 57 12 65 15
rect 57 8 60 12
rect 64 8 65 12
rect 57 6 65 8
<< pdiffusion >>
rect 37 94 43 95
rect 61 94 67 95
rect 15 92 21 93
rect 15 88 16 92
rect 20 88 21 92
rect 37 90 38 94
rect 42 90 45 94
rect 37 89 45 90
rect 15 83 21 88
rect 39 83 45 89
rect 3 82 11 83
rect 3 78 4 82
rect 8 78 11 82
rect 3 63 11 78
rect 13 63 23 83
rect 25 82 35 83
rect 25 78 28 82
rect 32 78 35 82
rect 25 63 35 78
rect 37 63 45 83
rect 39 55 45 63
rect 47 72 57 94
rect 47 68 50 72
rect 54 68 57 72
rect 47 62 57 68
rect 47 58 50 62
rect 54 58 57 62
rect 47 55 57 58
rect 59 90 62 94
rect 66 90 67 94
rect 59 89 67 90
rect 59 75 65 89
rect 59 55 67 75
rect 69 72 77 75
rect 69 68 72 72
rect 76 68 77 72
rect 69 62 77 68
rect 69 58 72 62
rect 76 58 77 62
rect 69 55 77 58
<< metal1 >>
rect -2 94 82 100
rect -2 92 38 94
rect -2 88 16 92
rect 20 90 38 92
rect 42 90 62 94
rect 66 90 82 94
rect 20 88 82 90
rect 67 82 68 83
rect 3 78 4 82
rect 8 78 28 82
rect 32 79 68 82
rect 72 79 73 83
rect 32 78 72 79
rect 8 42 12 73
rect 8 27 12 38
rect 18 52 22 73
rect 18 27 22 48
rect 28 42 32 73
rect 28 27 32 38
rect 38 22 42 78
rect 5 18 6 22
rect 10 18 42 22
rect 48 72 52 73
rect 72 72 76 73
rect 48 68 50 72
rect 54 68 55 72
rect 48 62 52 68
rect 72 62 76 68
rect 48 58 50 62
rect 54 58 55 62
rect 48 22 52 58
rect 72 42 76 58
rect 57 38 58 42
rect 62 38 76 42
rect 48 17 52 18
rect 72 22 76 38
rect 72 17 76 18
rect -2 8 36 12
rect 40 8 60 12
rect 64 8 82 12
rect -2 4 4 8
rect 8 4 12 8
rect 16 4 20 8
rect 24 4 82 8
rect -2 0 82 4
<< ntransistor >>
rect 13 15 15 34
rect 21 15 23 34
rect 29 15 31 34
rect 43 6 45 25
rect 55 6 57 25
rect 67 15 69 25
<< ptransistor >>
rect 11 63 13 83
rect 23 63 25 83
rect 35 63 37 83
rect 45 55 47 94
rect 57 55 59 94
rect 67 55 69 75
<< polycontact >>
rect 18 48 22 52
rect 8 38 12 42
rect 68 79 72 83
rect 28 38 32 42
rect 58 38 62 42
<< ndcontact >>
rect 6 18 10 22
rect 36 8 40 12
rect 48 18 52 22
rect 72 18 76 22
rect 60 8 64 12
<< pdcontact >>
rect 16 88 20 92
rect 38 90 42 94
rect 4 78 8 82
rect 28 78 32 82
rect 50 68 54 72
rect 50 58 54 62
rect 62 90 66 94
rect 72 68 76 72
rect 72 58 76 62
<< psubstratepcontact >>
rect 4 4 8 8
rect 12 4 16 8
rect 20 4 24 8
<< psubstratepdiff >>
rect 3 8 25 9
rect 3 4 4 8
rect 8 4 12 8
rect 16 4 20 8
rect 24 4 25 8
rect 3 3 25 4
<< labels >>
rlabel metal1 10 50 10 50 6 i0
rlabel metal1 30 50 30 50 6 i1
rlabel polycontact 20 50 20 50 6 i2
rlabel metal1 40 6 40 6 6 vss
rlabel metal1 50 45 50 45 6 nq
rlabel metal1 40 94 40 94 6 vdd
<< end >>
