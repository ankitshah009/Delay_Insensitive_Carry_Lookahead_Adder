magic
tech scmos
timestamp 1180600641
<< checkpaint >>
rect -22 -22 102 122
<< ab >>
rect 0 0 80 100
<< pwell >>
rect -4 -4 84 48
<< nwell >>
rect -4 48 84 104
<< polysilicon >>
rect 11 94 13 98
rect 23 94 25 98
rect 35 94 37 98
rect 47 94 49 98
rect 59 94 61 98
rect 11 53 13 56
rect 11 52 19 53
rect 11 48 14 52
rect 18 48 19 52
rect 11 47 19 48
rect 23 43 25 55
rect 35 43 37 55
rect 47 43 49 55
rect 59 43 61 55
rect 3 42 61 43
rect 3 38 4 42
rect 8 38 61 42
rect 3 37 61 38
rect 11 32 19 33
rect 11 28 14 32
rect 18 28 19 32
rect 11 27 19 28
rect 11 24 13 27
rect 23 25 25 37
rect 35 25 37 37
rect 47 25 49 37
rect 59 25 61 37
rect 11 2 13 6
rect 23 2 25 6
rect 35 2 37 6
rect 47 2 49 6
rect 59 2 61 6
<< ndiffusion >>
rect 18 24 23 25
rect 3 22 11 24
rect 3 18 4 22
rect 8 18 11 22
rect 3 6 11 18
rect 13 12 23 24
rect 13 8 16 12
rect 20 8 23 12
rect 13 6 23 8
rect 25 22 35 25
rect 25 18 28 22
rect 32 18 35 22
rect 25 6 35 18
rect 37 22 47 25
rect 37 18 40 22
rect 44 18 47 22
rect 37 12 47 18
rect 37 8 40 12
rect 44 8 47 12
rect 37 6 47 8
rect 49 22 59 25
rect 49 18 52 22
rect 56 18 59 22
rect 49 6 59 18
rect 61 22 69 25
rect 61 18 64 22
rect 68 18 69 22
rect 61 12 69 18
rect 61 8 64 12
rect 68 8 69 12
rect 61 6 69 8
<< pdiffusion >>
rect 3 82 11 94
rect 3 78 4 82
rect 8 78 11 82
rect 3 72 11 78
rect 3 68 4 72
rect 8 68 11 72
rect 3 62 11 68
rect 3 58 4 62
rect 8 58 11 62
rect 3 56 11 58
rect 13 92 23 94
rect 13 88 16 92
rect 20 88 23 92
rect 13 56 23 88
rect 18 55 23 56
rect 25 82 35 94
rect 25 78 28 82
rect 32 78 35 82
rect 25 72 35 78
rect 25 68 28 72
rect 32 68 35 72
rect 25 62 35 68
rect 25 58 28 62
rect 32 58 35 62
rect 25 55 35 58
rect 37 92 47 94
rect 37 88 40 92
rect 44 88 47 92
rect 37 82 47 88
rect 37 78 40 82
rect 44 78 47 82
rect 37 72 47 78
rect 37 68 40 72
rect 44 68 47 72
rect 37 62 47 68
rect 37 58 40 62
rect 44 58 47 62
rect 37 55 47 58
rect 49 82 59 94
rect 49 78 52 82
rect 56 78 59 82
rect 49 72 59 78
rect 49 68 52 72
rect 56 68 59 72
rect 49 62 59 68
rect 49 58 52 62
rect 56 58 59 62
rect 49 55 59 58
rect 61 92 69 94
rect 61 88 64 92
rect 68 88 69 92
rect 61 82 69 88
rect 61 78 64 82
rect 68 78 69 82
rect 61 77 69 78
rect 61 55 66 77
<< metal1 >>
rect -2 92 82 100
rect -2 88 16 92
rect 20 88 40 92
rect 44 88 64 92
rect 68 88 82 92
rect 4 82 8 83
rect 4 72 8 78
rect 4 62 8 68
rect 4 42 8 58
rect 13 48 14 52
rect 4 22 8 38
rect 13 28 14 32
rect 4 17 8 18
rect 18 17 22 83
rect 28 82 32 83
rect 28 72 32 78
rect 28 62 32 68
rect 28 42 32 58
rect 40 82 44 88
rect 40 72 44 78
rect 40 62 44 68
rect 40 57 44 58
rect 52 82 56 83
rect 52 72 56 78
rect 52 62 56 68
rect 64 82 68 88
rect 64 70 68 78
rect 72 70 76 71
rect 64 66 72 70
rect 52 42 56 58
rect 72 60 76 66
rect 72 55 76 56
rect 28 38 56 42
rect 28 22 32 38
rect 28 17 32 18
rect 40 22 44 23
rect 40 12 44 18
rect 52 22 56 38
rect 52 17 56 18
rect 64 36 68 37
rect 68 32 72 36
rect 76 32 77 36
rect 64 22 68 32
rect 64 12 68 18
rect -2 8 16 12
rect 20 8 40 12
rect 44 8 64 12
rect 68 8 82 12
rect -2 0 82 8
<< ntransistor >>
rect 11 6 13 24
rect 23 6 25 25
rect 35 6 37 25
rect 47 6 49 25
rect 59 6 61 25
<< ptransistor >>
rect 11 56 13 94
rect 23 55 25 94
rect 35 55 37 94
rect 47 55 49 94
rect 59 55 61 94
<< polycontact >>
rect 14 48 18 52
rect 4 38 8 42
rect 14 28 18 32
<< ndcontact >>
rect 4 18 8 22
rect 16 8 20 12
rect 28 18 32 22
rect 40 18 44 22
rect 40 8 44 12
rect 52 18 56 22
rect 64 18 68 22
rect 64 8 68 12
<< pdcontact >>
rect 4 78 8 82
rect 4 68 8 72
rect 4 58 8 62
rect 16 88 20 92
rect 28 78 32 82
rect 28 68 32 72
rect 28 58 32 62
rect 40 88 44 92
rect 40 78 44 82
rect 40 68 44 72
rect 40 58 44 62
rect 52 78 56 82
rect 52 68 56 72
rect 52 58 56 62
rect 64 88 68 92
rect 64 78 68 82
<< psubstratepcontact >>
rect 64 32 68 36
rect 72 32 76 36
<< nsubstratencontact >>
rect 72 66 76 70
rect 72 56 76 60
<< psubstratepdiff >>
rect 63 36 77 37
rect 63 32 64 36
rect 68 32 72 36
rect 76 32 77 36
rect 63 31 77 32
<< nsubstratendiff >>
rect 71 70 77 71
rect 71 66 72 70
rect 76 66 77 70
rect 71 60 77 66
rect 71 56 72 60
rect 76 56 77 60
rect 71 55 77 56
<< labels >>
rlabel metal1 30 50 30 50 6 q
rlabel metal1 20 50 20 50 6 i
rlabel metal1 40 6 40 6 6 vss
rlabel metal1 40 40 40 40 6 q
rlabel metal1 50 40 50 40 6 q
rlabel metal1 40 94 40 94 6 vdd
<< end >>
