magic
tech scmos
timestamp 1185039008
<< checkpaint >>
rect -22 -24 122 124
<< ab >>
rect 0 0 100 100
<< pwell >>
rect -2 -4 102 49
<< nwell >>
rect -2 49 102 104
<< polysilicon >>
rect 13 85 15 88
rect 25 85 27 88
rect 37 85 39 88
rect 73 95 75 98
rect 85 95 87 98
rect 61 75 63 78
rect 13 43 15 65
rect 7 42 15 43
rect 7 38 8 42
rect 12 38 15 42
rect 7 37 15 38
rect 13 25 15 37
rect 25 43 27 65
rect 37 43 39 65
rect 61 53 63 55
rect 61 52 69 53
rect 61 48 64 52
rect 68 48 69 52
rect 61 47 69 48
rect 25 42 33 43
rect 25 38 28 42
rect 32 38 33 42
rect 25 37 33 38
rect 37 42 43 43
rect 37 38 38 42
rect 42 38 43 42
rect 37 37 43 38
rect 25 25 27 37
rect 37 25 39 37
rect 61 25 63 47
rect 73 43 75 55
rect 85 43 87 55
rect 67 42 87 43
rect 67 38 68 42
rect 72 38 87 42
rect 67 37 87 38
rect 73 25 75 37
rect 85 25 87 37
rect 13 12 15 15
rect 25 12 27 15
rect 37 12 39 15
rect 61 12 63 15
rect 73 2 75 5
rect 85 2 87 5
<< ndiffusion >>
rect 29 32 35 33
rect 29 28 30 32
rect 34 28 35 32
rect 29 25 35 28
rect 5 15 13 25
rect 15 22 25 25
rect 15 18 18 22
rect 22 18 25 22
rect 15 15 25 18
rect 27 15 37 25
rect 39 22 47 25
rect 39 18 42 22
rect 46 18 47 22
rect 39 15 47 18
rect 53 22 61 25
rect 53 18 54 22
rect 58 18 61 22
rect 53 15 61 18
rect 63 15 73 25
rect 5 12 11 15
rect 65 12 73 15
rect 5 8 6 12
rect 10 8 11 12
rect 5 7 11 8
rect 65 8 66 12
rect 70 8 73 12
rect 65 5 73 8
rect 75 22 85 25
rect 75 18 78 22
rect 82 18 85 22
rect 75 5 85 18
rect 87 22 95 25
rect 87 18 90 22
rect 94 18 95 22
rect 87 12 95 18
rect 87 8 90 12
rect 94 8 95 12
rect 87 5 95 8
<< pdiffusion >>
rect 5 92 11 93
rect 5 88 6 92
rect 10 88 11 92
rect 41 92 47 93
rect 41 88 42 92
rect 46 88 47 92
rect 5 85 11 88
rect 41 85 47 88
rect 65 92 73 95
rect 65 88 66 92
rect 70 88 73 92
rect 5 65 13 85
rect 15 82 25 85
rect 15 78 18 82
rect 22 78 25 82
rect 15 72 25 78
rect 15 68 18 72
rect 22 68 25 72
rect 15 65 25 68
rect 27 65 37 85
rect 39 65 47 85
rect 65 82 73 88
rect 65 78 66 82
rect 70 78 73 82
rect 65 75 73 78
rect 53 62 61 75
rect 53 58 54 62
rect 58 58 61 62
rect 53 55 61 58
rect 63 55 73 75
rect 75 82 85 95
rect 75 78 78 82
rect 82 78 85 82
rect 75 72 85 78
rect 75 68 78 72
rect 82 68 85 72
rect 75 62 85 68
rect 75 58 78 62
rect 82 58 85 62
rect 75 55 85 58
rect 87 92 95 95
rect 87 88 90 92
rect 94 88 95 92
rect 87 82 95 88
rect 87 78 90 82
rect 94 78 95 82
rect 87 72 95 78
rect 87 68 90 72
rect 94 68 95 72
rect 87 62 95 68
rect 87 58 90 62
rect 94 58 95 62
rect 87 55 95 58
<< metal1 >>
rect -2 96 102 101
rect -2 92 18 96
rect 22 92 30 96
rect 34 92 54 96
rect 58 92 102 96
rect -2 88 6 92
rect 10 88 42 92
rect 46 88 66 92
rect 70 88 90 92
rect 94 88 102 92
rect -2 87 102 88
rect 17 82 23 83
rect 65 82 71 87
rect 7 42 13 82
rect 17 78 18 82
rect 22 78 58 82
rect 17 77 23 78
rect 18 73 22 77
rect 17 72 23 73
rect 54 72 58 78
rect 65 78 66 82
rect 70 78 71 82
rect 65 77 71 78
rect 77 82 83 83
rect 77 78 78 82
rect 82 78 83 82
rect 77 72 83 78
rect 17 68 18 72
rect 22 68 23 72
rect 17 67 23 68
rect 7 38 8 42
rect 12 38 13 42
rect 7 18 13 38
rect 18 32 22 67
rect 27 42 33 72
rect 27 38 28 42
rect 32 38 33 42
rect 27 37 33 38
rect 37 43 43 72
rect 54 68 68 72
rect 53 62 59 63
rect 53 58 54 62
rect 58 58 59 62
rect 53 57 59 58
rect 37 42 50 43
rect 37 38 38 42
rect 42 38 50 42
rect 54 42 58 57
rect 64 53 68 68
rect 77 68 78 72
rect 82 68 83 72
rect 77 62 83 68
rect 77 58 78 62
rect 82 58 83 62
rect 63 52 69 53
rect 63 48 64 52
rect 68 48 69 52
rect 63 47 69 48
rect 67 42 73 43
rect 54 38 68 42
rect 72 38 73 42
rect 37 37 50 38
rect 67 37 73 38
rect 46 33 50 37
rect 29 32 35 33
rect 18 28 30 32
rect 34 28 35 32
rect 46 28 52 33
rect 29 27 35 28
rect 48 27 52 28
rect 17 22 23 23
rect 41 22 47 23
rect 17 18 18 22
rect 22 18 42 22
rect 46 18 47 22
rect 17 17 23 18
rect 41 17 47 18
rect 53 22 59 23
rect 68 22 72 37
rect 53 18 54 22
rect 58 18 72 22
rect 77 22 83 58
rect 89 82 95 87
rect 89 78 90 82
rect 94 78 95 82
rect 89 72 95 78
rect 89 68 90 72
rect 94 68 95 72
rect 89 62 95 68
rect 89 58 90 62
rect 94 58 95 62
rect 89 57 95 58
rect 77 18 78 22
rect 82 18 83 22
rect 53 17 59 18
rect 77 17 83 18
rect 89 22 95 23
rect 89 18 90 22
rect 94 18 95 22
rect 89 13 95 18
rect -2 12 102 13
rect -2 8 6 12
rect 10 8 66 12
rect 70 8 90 12
rect 94 8 102 12
rect -2 4 18 8
rect 22 4 30 8
rect 34 4 42 8
rect 46 4 54 8
rect 58 4 102 8
rect -2 -1 102 4
<< ntransistor >>
rect 13 15 15 25
rect 25 15 27 25
rect 37 15 39 25
rect 61 15 63 25
rect 73 5 75 25
rect 85 5 87 25
<< ptransistor >>
rect 13 65 15 85
rect 25 65 27 85
rect 37 65 39 85
rect 61 55 63 75
rect 73 55 75 95
rect 85 55 87 95
<< polycontact >>
rect 8 38 12 42
rect 64 48 68 52
rect 28 38 32 42
rect 38 38 42 42
rect 68 38 72 42
<< ndcontact >>
rect 30 28 34 32
rect 18 18 22 22
rect 42 18 46 22
rect 54 18 58 22
rect 6 8 10 12
rect 66 8 70 12
rect 78 18 82 22
rect 90 18 94 22
rect 90 8 94 12
<< pdcontact >>
rect 6 88 10 92
rect 42 88 46 92
rect 66 88 70 92
rect 18 78 22 82
rect 18 68 22 72
rect 66 78 70 82
rect 54 58 58 62
rect 78 78 82 82
rect 78 68 82 72
rect 78 58 82 62
rect 90 88 94 92
rect 90 78 94 82
rect 90 68 94 72
rect 90 58 94 62
<< psubstratepcontact >>
rect 18 4 22 8
rect 30 4 34 8
rect 42 4 46 8
rect 54 4 58 8
<< nsubstratencontact >>
rect 18 92 22 96
rect 30 92 34 96
rect 54 92 58 96
<< psubstratepdiff >>
rect 17 8 59 9
rect 17 4 18 8
rect 22 4 30 8
rect 34 4 42 8
rect 46 4 54 8
rect 58 4 59 8
rect 17 3 59 4
<< nsubstratendiff >>
rect 17 96 35 97
rect 17 92 18 96
rect 22 92 30 96
rect 34 92 35 96
rect 53 96 59 97
rect 17 91 35 92
rect 53 92 54 96
rect 58 92 59 96
rect 53 85 59 92
<< labels >>
rlabel metal1 10 50 10 50 6 i2
rlabel metal1 10 50 10 50 6 i2
rlabel metal1 30 55 30 55 6 i1
rlabel metal1 40 55 40 55 6 i0
rlabel metal1 40 55 40 55 6 i0
rlabel metal1 30 55 30 55 6 i1
rlabel metal1 50 6 50 6 6 vss
rlabel metal1 50 6 50 6 6 vss
rlabel metal1 50 30 50 30 6 i0
rlabel metal1 50 30 50 30 6 i0
rlabel metal1 50 94 50 94 6 vdd
rlabel metal1 50 94 50 94 6 vdd
rlabel metal1 80 50 80 50 6 nq
rlabel metal1 80 50 80 50 6 nq
<< end >>
