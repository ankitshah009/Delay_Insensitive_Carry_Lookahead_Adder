.subckt noa22_x1 i0 i1 i2 nq vdd vss
*   SPICE3 file   created from noa22_x1.ext -      technology: scmos
m00 nq     i0     w1     vdd p w=39u  l=2.3636u ad=195p     pd=49u      as=234p     ps=64u
m01 w1     i1     nq     vdd p w=39u  l=2.3636u ad=234p     pd=64u      as=195p     ps=49u
m02 vdd    i2     w1     vdd p w=39u  l=2.3636u ad=312p     pd=94u      as=234p     ps=64u
m03 w2     i0     vss    vss n w=19u  l=2.3636u ad=95p      pd=29u      as=152p     ps=54u
m04 nq     i1     w2     vss n w=19u  l=2.3636u ad=95p      pd=29u      as=95p      ps=29u
m05 vss    i2     nq     vss n w=19u  l=2.3636u ad=152p     pd=54u      as=95p      ps=29u
C0  vdd    i1     0.016f
C1  w1     i0     0.024f
C2  w2     vss    0.019f
C3  i2     i0     0.082f
C4  vss    nq     0.070f
C5  vss    vdd    0.012f
C6  nq     w1     0.171f
C7  w1     vdd    0.191f
C8  nq     i2     0.283f
C9  vss    i1     0.047f
C10 w1     i1     0.013f
C11 vdd    i2     0.164f
C12 nq     i0     0.087f
C13 i2     i1     0.150f
C14 vdd    i0     0.014f
C15 i1     i0     0.310f
C16 nq     vdd    0.076f
C17 vss    i2     0.101f
C18 w2     i1     0.018f
C19 vss    i0     0.054f
C20 w1     i2     0.036f
C21 nq     i1     0.280f
C23 nq     vss    0.015f
C25 i2     vss    0.035f
C26 i1     vss    0.035f
C27 i0     vss    0.030f
.ends
