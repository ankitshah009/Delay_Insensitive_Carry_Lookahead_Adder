magic
tech scmos
timestamp 1185039010
<< checkpaint >>
rect -22 -24 92 124
<< ab >>
rect 0 0 70 100
<< pwell >>
rect -2 -4 72 49
<< nwell >>
rect -2 49 72 104
<< polysilicon >>
rect 11 95 13 98
rect 23 95 25 98
rect 35 95 37 98
rect 47 95 49 98
rect 11 43 13 55
rect 23 43 25 55
rect 7 42 13 43
rect 7 38 8 42
rect 12 38 13 42
rect 7 37 13 38
rect 17 42 25 43
rect 17 38 18 42
rect 22 38 25 42
rect 17 37 25 38
rect 11 25 13 37
rect 23 25 25 37
rect 35 43 37 55
rect 47 43 49 55
rect 35 42 43 43
rect 35 38 38 42
rect 42 38 43 42
rect 35 37 43 38
rect 47 42 53 43
rect 47 38 48 42
rect 52 38 53 42
rect 47 37 53 38
rect 35 25 37 37
rect 47 25 49 37
rect 11 2 13 5
rect 23 2 25 5
rect 35 2 37 5
rect 47 2 49 5
<< ndiffusion >>
rect 15 32 21 33
rect 15 28 16 32
rect 20 28 21 32
rect 15 25 21 28
rect 3 22 11 25
rect 3 18 4 22
rect 8 18 11 22
rect 3 5 11 18
rect 13 5 23 25
rect 25 22 35 25
rect 25 18 28 22
rect 32 18 35 22
rect 25 5 35 18
rect 37 12 47 25
rect 37 8 40 12
rect 44 8 47 12
rect 37 5 47 8
rect 49 22 57 25
rect 49 18 52 22
rect 56 18 57 22
rect 49 5 57 18
<< pdiffusion >>
rect 3 92 11 95
rect 3 88 4 92
rect 8 88 11 92
rect 3 55 11 88
rect 13 55 23 95
rect 25 82 35 95
rect 25 78 28 82
rect 32 78 35 82
rect 25 72 35 78
rect 25 68 28 72
rect 32 68 35 72
rect 25 62 35 68
rect 25 58 28 62
rect 32 58 35 62
rect 25 55 35 58
rect 37 55 47 95
rect 49 92 57 95
rect 49 88 52 92
rect 56 88 57 92
rect 49 73 57 88
rect 49 55 55 73
<< metal1 >>
rect -2 92 72 101
rect -2 88 4 92
rect 8 88 52 92
rect 56 88 72 92
rect -2 87 72 88
rect 27 82 33 83
rect 7 42 13 82
rect 7 38 8 42
rect 12 38 13 42
rect 7 37 13 38
rect 17 42 23 82
rect 17 38 18 42
rect 22 38 23 42
rect 17 37 23 38
rect 27 78 28 82
rect 32 78 33 82
rect 27 72 33 78
rect 27 68 28 72
rect 32 68 33 72
rect 27 62 33 68
rect 27 58 28 62
rect 32 58 33 62
rect 27 33 33 58
rect 15 32 33 33
rect 15 28 16 32
rect 20 28 33 32
rect 37 42 43 82
rect 37 38 38 42
rect 42 38 43 42
rect 37 28 43 38
rect 47 42 53 82
rect 61 60 67 87
rect 61 56 62 60
rect 66 56 67 60
rect 61 55 67 56
rect 47 38 48 42
rect 52 38 53 42
rect 47 28 53 38
rect 15 27 33 28
rect 3 22 9 23
rect 27 22 33 23
rect 51 22 57 23
rect 3 18 4 22
rect 8 18 28 22
rect 32 18 52 22
rect 56 18 57 22
rect 3 17 9 18
rect 27 17 33 18
rect 51 17 57 18
rect -2 12 72 13
rect -2 8 40 12
rect 44 8 72 12
rect -2 -1 72 8
<< ntransistor >>
rect 11 5 13 25
rect 23 5 25 25
rect 35 5 37 25
rect 47 5 49 25
<< ptransistor >>
rect 11 55 13 95
rect 23 55 25 95
rect 35 55 37 95
rect 47 55 49 95
<< polycontact >>
rect 8 38 12 42
rect 18 38 22 42
rect 38 38 42 42
rect 48 38 52 42
<< ndcontact >>
rect 16 28 20 32
rect 4 18 8 22
rect 28 18 32 22
rect 40 8 44 12
rect 52 18 56 22
<< pdcontact >>
rect 4 88 8 92
rect 28 78 32 82
rect 28 68 32 72
rect 28 58 32 62
rect 52 88 56 92
<< nsubstratencontact >>
rect 62 56 66 60
<< nsubstratendiff >>
rect 61 60 67 67
rect 61 56 62 60
rect 66 56 67 60
rect 61 55 67 56
<< labels >>
rlabel metal1 10 60 10 60 6 i0
rlabel metal1 10 60 10 60 6 i0
rlabel metal1 30 55 30 55 6 nq
rlabel metal1 20 60 20 60 6 i1
rlabel metal1 30 55 30 55 6 nq
rlabel metal1 20 60 20 60 6 i1
rlabel metal1 35 6 35 6 6 vss
rlabel metal1 35 6 35 6 6 vss
rlabel metal1 50 55 50 55 6 i2
rlabel metal1 40 55 40 55 6 i3
rlabel metal1 50 55 50 55 6 i2
rlabel metal1 40 55 40 55 6 i3
rlabel metal1 35 94 35 94 6 vdd
rlabel metal1 35 94 35 94 6 vdd
<< end >>
