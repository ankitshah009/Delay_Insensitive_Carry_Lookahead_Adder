magic
tech scmos
timestamp 1179385441
<< checkpaint >>
rect -22 -25 86 105
<< ab >>
rect 0 0 64 80
<< pwell >>
rect -4 -7 68 36
<< nwell >>
rect -4 36 68 87
<< polysilicon >>
rect 31 64 33 69
rect 41 64 43 69
rect 53 64 55 69
rect 9 54 11 59
rect 9 39 11 42
rect 31 39 33 48
rect 41 39 43 48
rect 53 45 55 48
rect 53 44 62 45
rect 53 40 57 44
rect 61 40 62 44
rect 53 39 62 40
rect 9 38 19 39
rect 9 37 14 38
rect 13 34 14 37
rect 18 34 19 38
rect 13 33 19 34
rect 31 38 37 39
rect 31 34 32 38
rect 36 34 37 38
rect 31 33 37 34
rect 41 38 47 39
rect 41 34 42 38
rect 46 34 47 38
rect 41 33 47 34
rect 13 30 15 33
rect 13 19 15 24
rect 31 23 33 33
rect 41 23 43 33
rect 53 28 55 39
rect 48 26 55 28
rect 48 23 50 26
rect 31 12 33 17
rect 41 11 43 16
rect 48 11 50 16
<< ndiffusion >>
rect 6 29 13 30
rect 6 25 7 29
rect 11 25 13 29
rect 6 24 13 25
rect 15 29 23 30
rect 15 25 18 29
rect 22 25 23 29
rect 15 24 23 25
rect 17 23 23 24
rect 17 22 31 23
rect 17 18 18 22
rect 22 18 25 22
rect 29 18 31 22
rect 17 17 31 18
rect 33 22 41 23
rect 33 18 35 22
rect 39 18 41 22
rect 33 17 41 18
rect 36 16 41 17
rect 43 16 48 23
rect 50 21 57 23
rect 50 17 52 21
rect 56 17 57 21
rect 50 16 57 17
<< pdiffusion >>
rect 45 72 51 73
rect 45 68 46 72
rect 50 68 51 72
rect 45 64 51 68
rect 26 61 31 64
rect 24 60 31 61
rect 24 56 25 60
rect 29 56 31 60
rect 4 48 9 54
rect 2 47 9 48
rect 2 43 3 47
rect 7 43 9 47
rect 2 42 9 43
rect 11 53 18 54
rect 11 49 13 53
rect 17 49 18 53
rect 11 42 18 49
rect 24 53 31 56
rect 24 49 25 53
rect 29 49 31 53
rect 24 48 31 49
rect 33 63 41 64
rect 33 59 35 63
rect 39 59 41 63
rect 33 48 41 59
rect 43 48 53 64
rect 55 63 62 64
rect 55 59 57 63
rect 61 59 62 63
rect 55 58 62 59
rect 55 48 60 58
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect -2 72 66 78
rect -2 68 46 72
rect 50 68 66 72
rect 13 53 17 68
rect 13 48 17 49
rect 25 60 29 61
rect 34 59 35 63
rect 39 59 57 63
rect 61 59 62 63
rect 25 53 29 56
rect 2 47 7 48
rect 2 43 3 47
rect 2 42 7 43
rect 2 31 6 42
rect 25 38 29 49
rect 34 49 46 55
rect 50 49 62 55
rect 34 39 38 49
rect 57 44 62 49
rect 61 40 62 44
rect 57 39 62 40
rect 13 34 14 38
rect 18 34 29 38
rect 2 29 14 31
rect 25 30 29 34
rect 32 38 38 39
rect 36 34 38 38
rect 32 33 38 34
rect 42 38 46 39
rect 42 30 46 34
rect 2 25 7 29
rect 11 25 14 29
rect 18 29 22 30
rect 25 26 39 30
rect 42 26 55 30
rect 2 17 6 25
rect 18 22 22 25
rect 35 22 39 26
rect 22 18 25 22
rect 29 18 30 22
rect 18 12 22 18
rect 35 17 39 18
rect 52 21 56 22
rect 52 12 56 17
rect -2 2 66 12
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
<< ntransistor >>
rect 13 24 15 30
rect 31 17 33 23
rect 41 16 43 23
rect 48 16 50 23
<< ptransistor >>
rect 9 42 11 54
rect 31 48 33 64
rect 41 48 43 64
rect 53 48 55 64
<< polycontact >>
rect 57 40 61 44
rect 14 34 18 38
rect 32 34 36 38
rect 42 34 46 38
<< ndcontact >>
rect 7 25 11 29
rect 18 25 22 29
rect 18 18 22 22
rect 25 18 29 22
rect 35 18 39 22
rect 52 17 56 21
<< pdcontact >>
rect 46 68 50 72
rect 25 56 29 60
rect 3 43 7 47
rect 13 49 17 53
rect 25 49 29 53
rect 35 59 39 63
rect 57 59 61 63
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
<< psubstratepdiff >>
rect 0 2 64 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 64 2
rect 0 -3 64 -2
<< nsubstratendiff >>
rect 0 82 64 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 64 82
rect 0 77 64 78
<< labels >>
rlabel metal1 4 32 4 32 6 z
rlabel metal1 12 28 12 28 6 z
rlabel metal1 32 6 32 6 6 vss
rlabel polycontact 44 36 44 36 6 a2
rlabel metal1 36 44 36 44 6 b
rlabel metal1 44 52 44 52 6 b
rlabel metal1 32 74 32 74 6 vdd
rlabel metal1 52 28 52 28 6 a2
rlabel metal1 52 52 52 52 6 a1
rlabel metal1 60 48 60 48 6 a1
rlabel metal1 48 61 48 61 6 n1
<< end >>
