magic
tech scmos
timestamp 1185039156
<< checkpaint >>
rect -22 -24 302 124
<< ab >>
rect 0 0 280 100
<< pwell >>
rect -2 -4 282 49
<< nwell >>
rect -2 49 282 104
<< polysilicon >>
rect 27 95 29 98
rect 39 95 41 98
rect 51 95 53 98
rect 59 95 61 98
rect 71 95 73 98
rect 83 95 85 98
rect 91 95 93 98
rect 195 95 197 98
rect 207 95 209 98
rect 219 95 221 98
rect 231 95 233 98
rect 243 95 245 98
rect 255 95 257 98
rect 267 95 269 98
rect 121 85 123 88
rect 147 85 149 88
rect 159 85 161 88
rect 171 85 173 88
rect 183 85 185 88
rect 15 69 17 72
rect 15 53 17 55
rect 7 52 17 53
rect 7 48 8 52
rect 12 48 17 52
rect 7 47 17 48
rect 15 37 17 47
rect 27 53 29 75
rect 39 73 41 75
rect 33 72 41 73
rect 33 68 34 72
rect 38 68 41 72
rect 33 67 41 68
rect 27 52 33 53
rect 27 48 28 52
rect 32 48 33 52
rect 27 47 33 48
rect 15 26 17 29
rect 27 23 29 47
rect 39 41 41 67
rect 51 63 53 75
rect 47 62 53 63
rect 47 58 48 62
rect 52 58 53 62
rect 47 57 53 58
rect 47 52 53 53
rect 47 48 48 52
rect 52 51 53 52
rect 59 51 61 75
rect 71 73 73 75
rect 83 73 85 75
rect 52 49 61 51
rect 52 48 53 49
rect 47 47 53 48
rect 39 39 53 41
rect 33 32 41 33
rect 33 28 34 32
rect 38 28 41 32
rect 33 27 41 28
rect 39 23 41 27
rect 51 23 53 39
rect 59 23 61 49
rect 69 71 73 73
rect 79 71 85 73
rect 69 33 71 71
rect 79 53 81 71
rect 91 63 93 75
rect 103 69 105 72
rect 85 62 93 63
rect 85 58 86 62
rect 90 58 93 62
rect 85 57 93 58
rect 195 73 197 75
rect 195 72 203 73
rect 195 68 198 72
rect 202 68 203 72
rect 195 67 203 68
rect 75 52 81 53
rect 75 48 76 52
rect 80 51 81 52
rect 103 51 105 55
rect 121 53 123 65
rect 147 63 149 65
rect 159 63 161 65
rect 171 63 173 65
rect 141 61 149 63
rect 157 62 163 63
rect 80 49 105 51
rect 80 48 81 49
rect 75 47 81 48
rect 79 39 81 47
rect 65 32 71 33
rect 65 28 66 32
rect 70 28 71 32
rect 65 27 71 28
rect 75 37 81 39
rect 85 42 93 43
rect 85 38 86 42
rect 90 38 93 42
rect 85 37 93 38
rect 103 37 105 49
rect 117 52 123 53
rect 117 48 118 52
rect 122 48 123 52
rect 117 47 123 48
rect 129 52 135 53
rect 129 48 130 52
rect 134 51 135 52
rect 141 51 143 61
rect 157 58 158 62
rect 162 58 163 62
rect 157 57 163 58
rect 169 62 175 63
rect 169 58 170 62
rect 174 58 175 62
rect 169 57 175 58
rect 167 52 173 53
rect 167 51 168 52
rect 134 49 168 51
rect 134 48 135 49
rect 129 47 135 48
rect 75 23 77 37
rect 81 32 87 33
rect 81 28 82 32
rect 86 28 87 32
rect 81 27 87 28
rect 71 21 77 23
rect 71 19 73 21
rect 83 19 85 27
rect 91 19 93 37
rect 103 26 105 29
rect 121 25 123 47
rect 141 29 143 49
rect 167 48 168 49
rect 172 51 173 52
rect 183 51 185 65
rect 207 63 209 75
rect 201 62 209 63
rect 201 58 202 62
rect 206 58 209 62
rect 201 57 209 58
rect 219 51 221 75
rect 231 73 233 75
rect 225 72 233 73
rect 225 68 226 72
rect 230 68 233 72
rect 225 67 233 68
rect 243 53 245 75
rect 243 52 251 53
rect 172 49 233 51
rect 172 48 173 49
rect 167 47 173 48
rect 147 42 153 43
rect 147 38 148 42
rect 152 41 153 42
rect 177 42 185 43
rect 177 41 178 42
rect 152 39 178 41
rect 152 38 153 39
rect 147 37 153 38
rect 177 38 178 39
rect 182 41 185 42
rect 219 42 227 43
rect 219 41 222 42
rect 182 39 222 41
rect 182 38 185 39
rect 177 37 185 38
rect 157 32 163 33
rect 141 27 149 29
rect 157 28 158 32
rect 162 28 163 32
rect 157 27 163 28
rect 169 32 175 33
rect 169 28 170 32
rect 174 28 175 32
rect 169 27 175 28
rect 147 25 149 27
rect 159 25 161 27
rect 171 25 173 27
rect 183 25 185 37
rect 219 38 222 39
rect 226 38 227 42
rect 219 37 227 38
rect 201 32 209 33
rect 201 28 202 32
rect 206 28 209 32
rect 201 27 209 28
rect 27 8 29 11
rect 39 8 41 11
rect 51 8 53 11
rect 59 8 61 11
rect 195 22 203 23
rect 195 18 198 22
rect 202 18 203 22
rect 195 17 203 18
rect 195 15 197 17
rect 207 15 209 27
rect 219 25 221 37
rect 231 25 233 49
rect 243 48 246 52
rect 250 48 251 52
rect 243 47 251 48
rect 255 43 257 55
rect 267 43 269 55
rect 245 42 269 43
rect 245 38 246 42
rect 250 38 269 42
rect 245 37 269 38
rect 243 32 251 33
rect 243 28 246 32
rect 250 28 251 32
rect 243 27 251 28
rect 243 25 245 27
rect 255 25 257 37
rect 267 25 269 37
rect 121 12 123 15
rect 147 12 149 15
rect 159 12 161 15
rect 171 12 173 15
rect 183 12 185 15
rect 71 4 73 7
rect 83 4 85 7
rect 91 4 93 7
rect 219 12 221 15
rect 231 12 233 15
rect 243 12 245 15
rect 195 2 197 5
rect 207 2 209 5
rect 255 2 257 5
rect 267 2 269 5
<< ndiffusion >>
rect 7 29 15 37
rect 17 34 25 37
rect 17 30 20 34
rect 24 30 25 34
rect 17 29 25 30
rect 7 22 13 29
rect 43 32 49 33
rect 43 28 44 32
rect 48 28 49 32
rect 43 23 49 28
rect 7 18 8 22
rect 12 18 13 22
rect 7 17 13 18
rect 19 22 27 23
rect 19 18 20 22
rect 24 18 27 22
rect 19 11 27 18
rect 29 11 39 23
rect 41 11 51 23
rect 53 11 59 23
rect 61 22 69 23
rect 61 18 64 22
rect 68 19 69 22
rect 95 36 103 37
rect 95 32 96 36
rect 100 32 103 36
rect 95 29 103 32
rect 105 29 117 37
rect 107 25 117 29
rect 95 22 101 23
rect 95 19 96 22
rect 68 18 71 19
rect 61 11 71 18
rect 63 7 71 11
rect 73 12 83 19
rect 73 8 76 12
rect 80 8 83 12
rect 73 7 83 8
rect 85 7 91 19
rect 93 18 96 19
rect 100 18 101 22
rect 93 9 101 18
rect 107 15 121 25
rect 123 22 133 25
rect 123 18 128 22
rect 132 18 133 22
rect 123 15 133 18
rect 139 22 147 25
rect 139 18 140 22
rect 144 18 147 22
rect 139 15 147 18
rect 149 15 159 25
rect 161 15 171 25
rect 173 22 183 25
rect 173 18 176 22
rect 180 18 183 22
rect 173 15 183 18
rect 185 15 193 25
rect 211 22 219 25
rect 211 18 212 22
rect 216 18 219 22
rect 211 15 219 18
rect 221 22 231 25
rect 221 18 224 22
rect 228 18 231 22
rect 221 15 231 18
rect 233 15 243 25
rect 245 22 255 25
rect 245 18 248 22
rect 252 18 255 22
rect 245 15 255 18
rect 107 12 117 15
rect 151 12 157 15
rect 93 7 97 9
rect 107 8 108 12
rect 112 8 117 12
rect 107 7 117 8
rect 151 8 152 12
rect 156 8 157 12
rect 151 7 157 8
rect 187 5 195 15
rect 197 12 207 15
rect 197 8 200 12
rect 204 8 207 12
rect 197 5 207 8
rect 209 5 217 15
rect 247 12 255 15
rect 247 8 248 12
rect 252 8 255 12
rect 247 5 255 8
rect 257 22 267 25
rect 257 18 260 22
rect 264 18 267 22
rect 257 5 267 18
rect 269 22 277 25
rect 269 18 272 22
rect 276 18 277 22
rect 269 12 277 18
rect 269 8 272 12
rect 276 8 277 12
rect 269 5 277 8
<< pdiffusion >>
rect 7 82 13 83
rect 7 78 8 82
rect 12 78 13 82
rect 7 69 13 78
rect 19 82 27 95
rect 19 78 20 82
rect 24 78 27 82
rect 19 75 27 78
rect 29 75 39 95
rect 41 75 51 95
rect 53 75 59 95
rect 61 82 71 95
rect 61 78 64 82
rect 68 78 71 82
rect 61 75 71 78
rect 73 92 83 95
rect 73 88 76 92
rect 80 88 83 92
rect 73 75 83 88
rect 85 75 91 95
rect 93 82 101 95
rect 93 78 96 82
rect 100 78 101 82
rect 93 75 101 78
rect 107 92 117 93
rect 107 88 108 92
rect 112 88 117 92
rect 151 94 157 95
rect 151 90 152 94
rect 156 90 157 94
rect 107 85 117 88
rect 151 85 157 90
rect 187 85 195 95
rect 7 55 15 69
rect 17 62 25 69
rect 17 58 20 62
rect 24 58 25 62
rect 17 55 25 58
rect 43 72 49 75
rect 43 68 44 72
rect 48 68 49 72
rect 43 67 49 68
rect 107 69 121 85
rect 95 62 103 69
rect 95 58 96 62
rect 100 58 103 62
rect 95 55 103 58
rect 105 65 121 69
rect 123 72 133 85
rect 123 68 128 72
rect 132 68 133 72
rect 123 65 133 68
rect 139 72 147 85
rect 139 68 140 72
rect 144 68 147 72
rect 139 65 147 68
rect 149 65 159 85
rect 161 65 171 85
rect 173 72 183 85
rect 173 68 176 72
rect 180 68 183 72
rect 173 65 183 68
rect 185 75 195 85
rect 197 92 207 95
rect 197 88 200 92
rect 204 88 207 92
rect 197 75 207 88
rect 209 82 219 95
rect 209 78 212 82
rect 216 78 219 82
rect 209 75 219 78
rect 221 82 231 95
rect 221 78 224 82
rect 228 78 231 82
rect 221 75 231 78
rect 233 75 243 95
rect 245 92 255 95
rect 245 88 248 92
rect 252 88 255 92
rect 245 82 255 88
rect 245 78 248 82
rect 252 78 255 82
rect 245 75 255 78
rect 185 65 193 75
rect 105 55 117 65
rect 247 72 255 75
rect 247 68 248 72
rect 252 68 255 72
rect 247 62 255 68
rect 247 58 248 62
rect 252 58 255 62
rect 247 55 255 58
rect 257 82 267 95
rect 257 78 260 82
rect 264 78 267 82
rect 257 72 267 78
rect 257 68 260 72
rect 264 68 267 72
rect 257 62 267 68
rect 257 58 260 62
rect 264 58 267 62
rect 257 55 267 58
rect 269 92 277 95
rect 269 88 272 92
rect 276 88 277 92
rect 269 82 277 88
rect 269 78 272 82
rect 276 78 277 82
rect 269 72 277 78
rect 269 68 272 72
rect 276 68 277 72
rect 269 62 277 68
rect 269 58 272 62
rect 276 58 277 62
rect 269 55 277 58
<< metal1 >>
rect -2 96 282 101
rect -2 92 126 96
rect 130 92 140 96
rect 144 94 164 96
rect 144 92 152 94
rect -2 88 76 92
rect 80 88 108 92
rect 112 90 152 92
rect 156 92 164 94
rect 168 92 176 96
rect 180 92 282 96
rect 156 90 200 92
rect 112 88 200 90
rect 204 88 248 92
rect 252 88 272 92
rect 276 88 282 92
rect -2 87 282 88
rect 7 82 13 87
rect 7 78 8 82
rect 12 78 13 82
rect 7 77 13 78
rect 19 82 69 83
rect 19 78 20 82
rect 24 78 64 82
rect 68 78 69 82
rect 19 77 69 78
rect 95 82 162 83
rect 211 82 217 83
rect 95 78 96 82
rect 100 78 163 82
rect 95 77 163 78
rect 95 73 101 77
rect 8 72 39 73
rect 7 68 34 72
rect 38 68 39 72
rect 7 67 39 68
rect 43 72 112 73
rect 127 72 133 73
rect 43 68 44 72
rect 48 68 113 72
rect 43 67 113 68
rect 7 52 13 67
rect 19 62 53 63
rect 7 48 8 52
rect 12 48 13 52
rect 7 28 13 48
rect 17 58 20 62
rect 24 58 48 62
rect 52 58 53 62
rect 17 57 53 58
rect 17 35 23 57
rect 27 52 33 53
rect 27 48 28 52
rect 32 48 33 52
rect 27 40 33 48
rect 38 52 53 53
rect 38 48 48 52
rect 52 48 53 52
rect 38 47 53 48
rect 57 43 63 67
rect 78 62 91 63
rect 54 42 63 43
rect 53 38 63 42
rect 67 53 73 62
rect 78 58 86 62
rect 90 58 91 62
rect 78 57 91 58
rect 95 62 101 63
rect 95 58 96 62
rect 100 58 103 62
rect 95 57 103 58
rect 86 53 90 57
rect 67 52 81 53
rect 67 48 76 52
rect 80 48 81 52
rect 67 47 81 48
rect 86 47 92 53
rect 67 38 73 47
rect 86 43 90 47
rect 78 42 91 43
rect 78 38 86 42
rect 90 38 91 42
rect 53 37 62 38
rect 78 37 91 38
rect 97 37 103 57
rect 17 34 25 35
rect 17 30 20 34
rect 24 33 25 34
rect 53 33 59 37
rect 95 36 103 37
rect 95 33 96 36
rect 24 32 39 33
rect 24 30 34 32
rect 19 29 34 30
rect 20 28 34 29
rect 38 28 39 32
rect 20 27 39 28
rect 43 32 59 33
rect 43 28 44 32
rect 48 28 59 32
rect 65 32 96 33
rect 100 32 103 36
rect 65 28 66 32
rect 70 28 82 32
rect 86 28 101 32
rect 43 27 58 28
rect 65 27 100 28
rect 107 23 113 67
rect 7 22 13 23
rect 7 18 8 22
rect 12 18 13 22
rect 7 13 13 18
rect 19 22 25 23
rect 63 22 69 23
rect 19 18 20 22
rect 24 18 64 22
rect 68 18 69 22
rect 19 17 25 18
rect 63 17 69 18
rect 95 22 113 23
rect 95 18 96 22
rect 100 18 113 22
rect 117 52 123 72
rect 117 48 118 52
rect 122 48 123 52
rect 117 18 123 48
rect 127 68 128 72
rect 132 68 133 72
rect 127 53 133 68
rect 139 72 145 73
rect 139 68 140 72
rect 144 71 152 72
rect 144 68 153 71
rect 139 67 153 68
rect 140 66 153 67
rect 127 52 135 53
rect 127 48 130 52
rect 134 48 135 52
rect 127 47 135 48
rect 127 22 133 47
rect 147 42 153 66
rect 147 38 148 42
rect 152 38 153 42
rect 147 24 153 38
rect 157 62 163 77
rect 211 78 212 82
rect 216 78 217 82
rect 211 73 217 78
rect 223 82 240 83
rect 247 82 253 87
rect 259 82 265 83
rect 223 78 224 82
rect 228 78 241 82
rect 223 77 241 78
rect 175 72 192 73
rect 197 72 217 73
rect 225 72 231 73
rect 175 68 176 72
rect 180 68 193 72
rect 175 67 193 68
rect 197 68 198 72
rect 202 68 217 72
rect 197 67 217 68
rect 187 63 193 67
rect 157 58 158 62
rect 162 58 163 62
rect 157 32 163 58
rect 169 62 182 63
rect 187 62 207 63
rect 169 58 170 62
rect 174 58 183 62
rect 169 57 183 58
rect 157 28 158 32
rect 162 28 163 32
rect 167 52 173 53
rect 167 48 168 52
rect 172 48 173 52
rect 167 33 173 48
rect 177 42 183 57
rect 177 38 178 42
rect 182 38 183 42
rect 177 37 183 38
rect 187 58 202 62
rect 206 58 207 62
rect 187 57 207 58
rect 187 33 193 57
rect 167 32 175 33
rect 167 28 170 32
rect 174 28 175 32
rect 157 27 163 28
rect 169 27 175 28
rect 187 32 207 33
rect 187 28 202 32
rect 206 28 207 32
rect 187 27 207 28
rect 140 23 153 24
rect 187 23 193 27
rect 211 23 217 67
rect 223 68 226 72
rect 230 68 231 72
rect 223 67 231 68
rect 223 43 229 67
rect 221 42 229 43
rect 221 38 222 42
rect 226 38 229 42
rect 235 43 241 77
rect 247 78 248 82
rect 252 78 253 82
rect 247 72 253 78
rect 247 68 248 72
rect 252 68 253 72
rect 247 62 253 68
rect 247 58 248 62
rect 252 58 253 62
rect 247 57 253 58
rect 257 78 260 82
rect 264 78 265 82
rect 257 77 265 78
rect 271 82 277 87
rect 271 78 272 82
rect 276 78 277 82
rect 257 73 263 77
rect 257 72 265 73
rect 257 68 260 72
rect 264 68 265 72
rect 257 67 265 68
rect 271 72 277 78
rect 271 68 272 72
rect 276 68 277 72
rect 257 63 263 67
rect 257 62 265 63
rect 257 58 260 62
rect 264 58 265 62
rect 257 57 265 58
rect 271 62 277 68
rect 271 58 272 62
rect 276 58 277 62
rect 271 57 277 58
rect 257 53 263 57
rect 245 52 264 53
rect 245 48 246 52
rect 250 48 264 52
rect 245 47 264 48
rect 235 42 251 43
rect 235 38 246 42
rect 250 38 251 42
rect 221 37 227 38
rect 235 37 251 38
rect 235 23 241 37
rect 257 33 263 47
rect 245 32 264 33
rect 245 28 246 32
rect 250 28 264 32
rect 245 27 264 28
rect 257 23 263 27
rect 127 18 128 22
rect 132 18 133 22
rect 95 17 112 18
rect 127 17 133 18
rect 139 22 153 23
rect 139 18 140 22
rect 144 19 153 22
rect 175 22 193 23
rect 144 18 152 19
rect 175 18 176 22
rect 180 18 193 22
rect 197 22 217 23
rect 197 18 198 22
rect 202 18 212 22
rect 216 18 217 22
rect 139 17 145 18
rect 175 17 192 18
rect 197 17 217 18
rect 223 22 241 23
rect 223 18 224 22
rect 228 18 241 22
rect 247 22 253 23
rect 247 18 248 22
rect 252 18 253 22
rect 257 22 265 23
rect 257 18 260 22
rect 264 18 265 22
rect 223 17 240 18
rect 247 13 253 18
rect 259 17 265 18
rect 271 22 277 23
rect 271 18 272 22
rect 276 18 277 22
rect 271 13 277 18
rect -2 12 282 13
rect -2 8 76 12
rect 80 8 108 12
rect 112 8 152 12
rect 156 8 200 12
rect 204 8 248 12
rect 252 8 272 12
rect 276 8 282 12
rect -2 4 126 8
rect 130 4 140 8
rect 144 4 164 8
rect 168 4 176 8
rect 180 4 224 8
rect 228 4 236 8
rect 240 4 282 8
rect -2 -1 282 4
<< ntransistor >>
rect 15 29 17 37
rect 27 11 29 23
rect 39 11 41 23
rect 51 11 53 23
rect 59 11 61 23
rect 103 29 105 37
rect 71 7 73 19
rect 83 7 85 19
rect 91 7 93 19
rect 121 15 123 25
rect 147 15 149 25
rect 159 15 161 25
rect 171 15 173 25
rect 183 15 185 25
rect 219 15 221 25
rect 231 15 233 25
rect 243 15 245 25
rect 195 5 197 15
rect 207 5 209 15
rect 255 5 257 25
rect 267 5 269 25
<< ptransistor >>
rect 27 75 29 95
rect 39 75 41 95
rect 51 75 53 95
rect 59 75 61 95
rect 71 75 73 95
rect 83 75 85 95
rect 91 75 93 95
rect 15 55 17 69
rect 103 55 105 69
rect 121 65 123 85
rect 147 65 149 85
rect 159 65 161 85
rect 171 65 173 85
rect 183 65 185 85
rect 195 75 197 95
rect 207 75 209 95
rect 219 75 221 95
rect 231 75 233 95
rect 243 75 245 95
rect 255 55 257 95
rect 267 55 269 95
<< polycontact >>
rect 8 48 12 52
rect 34 68 38 72
rect 28 48 32 52
rect 48 58 52 62
rect 48 48 52 52
rect 34 28 38 32
rect 86 58 90 62
rect 198 68 202 72
rect 76 48 80 52
rect 66 28 70 32
rect 86 38 90 42
rect 118 48 122 52
rect 130 48 134 52
rect 158 58 162 62
rect 170 58 174 62
rect 82 28 86 32
rect 168 48 172 52
rect 202 58 206 62
rect 226 68 230 72
rect 148 38 152 42
rect 178 38 182 42
rect 158 28 162 32
rect 170 28 174 32
rect 222 38 226 42
rect 202 28 206 32
rect 198 18 202 22
rect 246 48 250 52
rect 246 38 250 42
rect 246 28 250 32
<< ndcontact >>
rect 20 30 24 34
rect 44 28 48 32
rect 8 18 12 22
rect 20 18 24 22
rect 64 18 68 22
rect 96 32 100 36
rect 76 8 80 12
rect 96 18 100 22
rect 128 18 132 22
rect 140 18 144 22
rect 176 18 180 22
rect 212 18 216 22
rect 224 18 228 22
rect 248 18 252 22
rect 108 8 112 12
rect 152 8 156 12
rect 200 8 204 12
rect 248 8 252 12
rect 260 18 264 22
rect 272 18 276 22
rect 272 8 276 12
<< pdcontact >>
rect 8 78 12 82
rect 20 78 24 82
rect 64 78 68 82
rect 76 88 80 92
rect 96 78 100 82
rect 108 88 112 92
rect 152 90 156 94
rect 20 58 24 62
rect 44 68 48 72
rect 96 58 100 62
rect 128 68 132 72
rect 140 68 144 72
rect 176 68 180 72
rect 200 88 204 92
rect 212 78 216 82
rect 224 78 228 82
rect 248 88 252 92
rect 248 78 252 82
rect 248 68 252 72
rect 248 58 252 62
rect 260 78 264 82
rect 260 68 264 72
rect 260 58 264 62
rect 272 88 276 92
rect 272 78 276 82
rect 272 68 276 72
rect 272 58 276 62
<< psubstratepcontact >>
rect 126 4 130 8
rect 140 4 144 8
rect 164 4 168 8
rect 176 4 180 8
rect 224 4 228 8
rect 236 4 240 8
<< nsubstratencontact >>
rect 126 92 130 96
rect 140 92 144 96
rect 164 92 168 96
rect 176 92 180 96
<< psubstratepdiff >>
rect 125 8 145 9
rect 125 4 126 8
rect 130 4 140 8
rect 144 4 145 8
rect 163 8 181 9
rect 125 3 145 4
rect 163 4 164 8
rect 168 4 176 8
rect 180 4 181 8
rect 223 8 241 9
rect 163 3 181 4
rect 223 4 224 8
rect 228 4 236 8
rect 240 4 241 8
rect 223 3 241 4
<< nsubstratendiff >>
rect 125 96 145 97
rect 125 92 126 96
rect 130 92 140 96
rect 144 92 145 96
rect 163 96 181 97
rect 125 91 145 92
rect 163 92 164 96
rect 168 92 176 96
rect 180 92 181 96
rect 163 91 181 92
<< labels >>
rlabel polycontact 30 50 30 50 6 i2
rlabel polycontact 10 50 10 50 6 cmd1
rlabel polycontact 30 50 30 50 6 i2
rlabel polycontact 10 50 10 50 6 cmd1
rlabel metal1 80 40 80 40 6 i0
rlabel metal1 80 40 80 40 6 i0
rlabel polycontact 50 50 50 50 6 i1
rlabel metal1 70 50 70 50 6 cmd0
rlabel metal1 90 50 90 50 6 i0
rlabel metal1 90 50 90 50 6 i0
rlabel metal1 70 50 70 50 6 cmd0
rlabel polycontact 50 50 50 50 6 i1
rlabel metal1 80 60 80 60 6 i0
rlabel metal1 80 60 80 60 6 i0
rlabel metal1 120 45 120 45 6 ck
rlabel metal1 120 45 120 45 6 ck
rlabel metal1 140 6 140 6 6 vss
rlabel metal1 140 6 140 6 6 vss
rlabel metal1 140 94 140 94 6 vdd
rlabel metal1 140 94 140 94 6 vdd
rlabel metal1 260 50 260 50 6 q
rlabel metal1 260 50 260 50 6 q
<< end >>
