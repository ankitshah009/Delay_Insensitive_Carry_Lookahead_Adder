magic
tech scmos
timestamp 1179386417
<< checkpaint >>
rect -22 -25 94 105
<< ab >>
rect 0 0 72 80
<< pwell >>
rect -4 -7 76 36
<< nwell >>
rect -4 36 76 87
<< polysilicon >>
rect 9 66 11 71
rect 19 66 21 71
rect 29 66 31 71
rect 39 66 41 71
rect 50 56 52 61
rect 60 56 62 61
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 39 39 41 42
rect 50 39 52 42
rect 60 39 62 42
rect 9 38 15 39
rect 9 34 10 38
rect 14 34 15 38
rect 9 33 15 34
rect 19 38 31 39
rect 19 34 26 38
rect 30 34 31 38
rect 19 33 31 34
rect 12 30 14 33
rect 19 30 21 33
rect 29 30 31 33
rect 36 38 52 39
rect 36 34 42 38
rect 46 37 52 38
rect 56 38 62 39
rect 46 34 47 37
rect 36 33 47 34
rect 56 34 57 38
rect 61 34 62 38
rect 56 33 62 34
rect 36 30 38 33
rect 12 12 14 17
rect 19 12 21 17
rect 29 12 31 17
rect 36 12 38 17
<< ndiffusion >>
rect 3 17 12 30
rect 14 17 19 30
rect 21 22 29 30
rect 21 18 23 22
rect 27 18 29 22
rect 21 17 29 18
rect 31 17 36 30
rect 38 17 47 30
rect 3 12 10 17
rect 40 12 47 17
rect 3 8 5 12
rect 9 8 10 12
rect 3 7 10 8
rect 40 8 41 12
rect 45 8 47 12
rect 40 7 47 8
<< pdiffusion >>
rect 2 65 9 66
rect 2 61 3 65
rect 7 61 9 65
rect 2 42 9 61
rect 11 62 19 66
rect 11 58 13 62
rect 17 58 19 62
rect 11 54 19 58
rect 11 50 13 54
rect 17 50 19 54
rect 11 42 19 50
rect 21 65 29 66
rect 21 61 23 65
rect 27 61 29 65
rect 21 42 29 61
rect 31 62 39 66
rect 31 58 33 62
rect 37 58 39 62
rect 31 54 39 58
rect 31 50 33 54
rect 37 50 39 54
rect 31 42 39 50
rect 41 65 48 66
rect 41 61 43 65
rect 47 61 48 65
rect 41 56 48 61
rect 41 42 50 56
rect 52 54 60 56
rect 52 50 54 54
rect 58 50 60 54
rect 52 42 60 50
rect 62 55 70 56
rect 62 51 64 55
rect 68 51 70 55
rect 62 47 70 51
rect 62 43 64 47
rect 68 43 70 47
rect 62 42 70 43
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect -2 68 74 78
rect 3 65 7 68
rect 23 65 27 68
rect 3 60 7 61
rect 13 62 17 63
rect 43 65 47 68
rect 23 60 27 61
rect 33 62 38 63
rect 13 54 17 58
rect 37 58 38 62
rect 43 60 47 61
rect 33 54 38 58
rect 64 55 68 68
rect 2 50 13 54
rect 17 50 33 54
rect 37 50 54 54
rect 58 50 59 54
rect 2 22 6 50
rect 64 47 68 51
rect 25 42 57 46
rect 64 42 68 43
rect 10 38 21 39
rect 14 34 21 38
rect 25 38 31 42
rect 25 34 26 38
rect 30 34 31 38
rect 41 34 42 38
rect 46 34 47 38
rect 53 34 57 42
rect 61 34 63 38
rect 10 33 21 34
rect 17 30 21 33
rect 41 30 47 34
rect 17 26 47 30
rect 2 18 23 22
rect 27 18 31 22
rect -2 8 5 12
rect 9 8 41 12
rect 45 8 74 12
rect -2 2 74 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
<< ntransistor >>
rect 12 17 14 30
rect 19 17 21 30
rect 29 17 31 30
rect 36 17 38 30
<< ptransistor >>
rect 9 42 11 66
rect 19 42 21 66
rect 29 42 31 66
rect 39 42 41 66
rect 50 42 52 56
rect 60 42 62 56
<< polycontact >>
rect 10 34 14 38
rect 26 34 30 38
rect 42 34 46 38
rect 57 34 61 38
<< ndcontact >>
rect 23 18 27 22
rect 5 8 9 12
rect 41 8 45 12
<< pdcontact >>
rect 3 61 7 65
rect 13 58 17 62
rect 13 50 17 54
rect 23 61 27 65
rect 33 58 37 62
rect 33 50 37 54
rect 43 61 47 65
rect 54 50 58 54
rect 64 51 68 55
rect 64 43 68 47
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
<< psubstratepdiff >>
rect 0 2 72 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 72 2
rect 0 -3 72 -2
<< nsubstratendiff >>
rect 0 82 72 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 72 82
rect 0 77 72 78
<< labels >>
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 20 12 20 6 z
rlabel metal1 20 20 20 20 6 z
rlabel metal1 20 28 20 28 6 a
rlabel polycontact 12 36 12 36 6 a
rlabel metal1 20 52 20 52 6 z
rlabel metal1 12 52 12 52 6 z
rlabel metal1 36 6 36 6 6 vss
rlabel metal1 28 20 28 20 6 z
rlabel metal1 28 28 28 28 6 a
rlabel metal1 36 28 36 28 6 a
rlabel metal1 28 40 28 40 6 b
rlabel metal1 36 44 36 44 6 b
rlabel metal1 28 52 28 52 6 z
rlabel metal1 36 56 36 56 6 z
rlabel metal1 36 74 36 74 6 vdd
rlabel metal1 44 32 44 32 6 a
rlabel metal1 44 44 44 44 6 b
rlabel metal1 52 44 52 44 6 b
rlabel metal1 52 52 52 52 6 z
rlabel metal1 44 52 44 52 6 z
rlabel polycontact 60 36 60 36 6 b
<< end >>
