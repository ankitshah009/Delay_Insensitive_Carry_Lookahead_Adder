magic
tech scmos
timestamp 1179387554
<< checkpaint >>
rect -22 -25 150 105
<< ab >>
rect 0 0 128 80
<< pwell >>
rect -4 -7 132 36
<< nwell >>
rect -4 36 132 87
<< polysilicon >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 39 70 41 74
rect 72 70 74 74
rect 79 70 81 74
rect 89 70 91 74
rect 107 70 109 74
rect 117 70 119 74
rect 49 62 51 67
rect 39 49 41 52
rect 49 49 51 52
rect 39 48 51 49
rect 39 47 43 48
rect 42 44 43 47
rect 47 47 51 48
rect 47 44 48 47
rect 42 43 48 44
rect 57 42 63 43
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 57 39 58 42
rect 9 38 15 39
rect 9 34 10 38
rect 14 34 15 38
rect 9 33 15 34
rect 19 38 25 39
rect 19 34 20 38
rect 24 34 25 38
rect 29 38 58 39
rect 62 38 63 42
rect 72 39 74 42
rect 29 37 63 38
rect 69 38 75 39
rect 19 33 25 34
rect 10 24 12 33
rect 19 29 21 33
rect 37 29 39 37
rect 69 34 70 38
rect 74 34 75 38
rect 69 33 75 34
rect 49 32 55 33
rect 17 27 21 29
rect 17 24 19 27
rect 27 24 29 29
rect 49 28 50 32
rect 54 28 55 32
rect 69 30 71 33
rect 79 30 81 42
rect 89 39 91 42
rect 89 38 95 39
rect 89 34 90 38
rect 94 35 95 38
rect 107 35 109 42
rect 117 39 119 42
rect 94 34 109 35
rect 89 33 109 34
rect 113 38 119 39
rect 113 34 114 38
rect 118 34 119 38
rect 113 33 119 34
rect 101 30 103 33
rect 49 27 55 28
rect 49 23 51 27
rect 37 12 39 16
rect 88 21 94 22
rect 88 17 89 21
rect 93 17 94 21
rect 117 27 119 33
rect 88 16 94 17
rect 10 6 12 11
rect 17 6 19 11
rect 27 8 29 11
rect 49 8 51 12
rect 69 11 71 16
rect 79 13 81 16
rect 88 13 90 16
rect 101 14 103 19
rect 79 11 90 13
rect 27 6 51 8
rect 117 11 119 16
<< ndiffusion >>
rect 32 24 37 29
rect 2 12 10 24
rect 2 8 3 12
rect 7 11 10 12
rect 12 11 17 24
rect 19 22 27 24
rect 19 18 21 22
rect 25 18 27 22
rect 19 11 27 18
rect 29 23 37 24
rect 29 19 31 23
rect 35 19 37 23
rect 29 16 37 19
rect 39 23 47 29
rect 39 17 49 23
rect 39 16 42 17
rect 29 11 34 16
rect 41 13 42 16
rect 46 13 49 17
rect 41 12 49 13
rect 51 22 58 23
rect 64 22 69 30
rect 51 18 53 22
rect 57 18 58 22
rect 51 17 58 18
rect 62 21 69 22
rect 62 17 63 21
rect 67 17 69 21
rect 51 12 56 17
rect 62 16 69 17
rect 71 29 79 30
rect 71 25 73 29
rect 77 25 79 29
rect 71 16 79 25
rect 81 29 88 30
rect 81 25 83 29
rect 87 25 88 29
rect 81 24 88 25
rect 94 29 101 30
rect 94 25 95 29
rect 99 25 101 29
rect 94 24 101 25
rect 81 16 86 24
rect 96 19 101 24
rect 103 27 115 30
rect 103 19 117 27
rect 7 8 8 11
rect 2 7 8 8
rect 105 16 117 19
rect 119 22 124 27
rect 119 21 126 22
rect 119 17 121 21
rect 125 17 126 21
rect 119 16 126 17
rect 105 12 115 16
rect 105 8 108 12
rect 112 8 115 12
rect 105 7 115 8
<< pdiffusion >>
rect 4 64 9 70
rect 2 63 9 64
rect 2 59 3 63
rect 7 59 9 63
rect 2 58 9 59
rect 4 42 9 58
rect 11 55 19 70
rect 11 51 13 55
rect 17 51 19 55
rect 11 42 19 51
rect 21 47 29 70
rect 21 43 23 47
rect 27 43 29 47
rect 21 42 29 43
rect 31 69 39 70
rect 31 65 33 69
rect 37 65 39 69
rect 31 62 39 65
rect 31 58 33 62
rect 37 58 39 62
rect 31 52 39 58
rect 41 62 46 70
rect 67 63 72 70
rect 65 62 72 63
rect 41 58 49 62
rect 41 54 43 58
rect 47 54 49 58
rect 41 52 49 54
rect 51 61 58 62
rect 51 57 53 61
rect 57 57 58 61
rect 51 52 58 57
rect 65 58 66 62
rect 70 58 72 62
rect 65 55 72 58
rect 31 42 37 52
rect 65 51 66 55
rect 70 51 72 55
rect 65 42 72 51
rect 74 42 79 70
rect 81 63 89 70
rect 81 59 83 63
rect 87 59 89 63
rect 81 56 89 59
rect 81 52 83 56
rect 87 52 89 56
rect 81 42 89 52
rect 91 65 96 70
rect 91 64 98 65
rect 91 60 93 64
rect 97 60 98 64
rect 91 57 98 60
rect 91 53 93 57
rect 97 53 98 57
rect 91 52 98 53
rect 91 42 96 52
rect 102 48 107 70
rect 100 47 107 48
rect 100 43 101 47
rect 105 43 107 47
rect 100 42 107 43
rect 109 69 117 70
rect 109 65 111 69
rect 115 65 117 69
rect 109 62 117 65
rect 109 58 111 62
rect 115 58 117 62
rect 109 42 117 58
rect 119 55 124 70
rect 119 54 126 55
rect 119 50 121 54
rect 125 50 126 54
rect 119 47 126 50
rect 119 43 121 47
rect 125 43 126 47
rect 119 42 126 43
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect 118 78 122 82
rect 126 78 130 82
rect -2 69 130 78
rect -2 68 33 69
rect 32 65 33 68
rect 37 68 111 69
rect 37 65 38 68
rect 2 59 3 63
rect 7 59 27 63
rect 23 55 27 59
rect 32 62 38 65
rect 32 58 33 62
rect 37 58 38 62
rect 53 61 57 68
rect 43 58 47 59
rect 2 51 13 55
rect 17 51 18 55
rect 23 54 43 55
rect 53 56 57 57
rect 66 62 70 68
rect 110 65 111 68
rect 115 68 130 69
rect 115 65 116 68
rect 23 51 47 54
rect 66 55 70 58
rect 83 63 87 64
rect 83 56 87 59
rect 2 50 18 51
rect 2 22 6 50
rect 10 43 23 47
rect 27 43 28 47
rect 10 38 14 43
rect 32 38 36 51
rect 66 50 70 51
rect 74 52 83 55
rect 74 51 87 52
rect 92 60 93 64
rect 97 60 98 64
rect 92 57 98 60
rect 110 62 116 65
rect 110 58 111 62
rect 115 58 116 62
rect 92 53 93 57
rect 97 55 98 57
rect 97 54 126 55
rect 97 53 121 54
rect 92 51 121 53
rect 41 44 43 48
rect 47 44 54 48
rect 74 46 78 51
rect 125 50 126 54
rect 121 47 126 50
rect 41 42 54 44
rect 61 43 78 46
rect 19 34 20 38
rect 24 34 44 38
rect 10 30 14 34
rect 10 26 35 30
rect 31 23 35 26
rect 2 18 21 22
rect 25 18 26 22
rect 40 24 44 34
rect 50 32 54 42
rect 58 42 78 43
rect 62 38 65 42
rect 82 41 94 47
rect 90 38 94 41
rect 58 37 65 38
rect 50 27 54 28
rect 61 29 65 37
rect 69 34 70 38
rect 74 34 86 38
rect 82 29 86 34
rect 90 33 94 34
rect 98 43 101 47
rect 105 43 106 47
rect 98 29 102 43
rect 114 38 118 47
rect 125 43 126 47
rect 121 42 126 43
rect 114 31 118 34
rect 61 25 73 29
rect 77 25 78 29
rect 82 25 83 29
rect 87 25 95 29
rect 99 25 102 29
rect 106 25 118 31
rect 40 22 57 24
rect 40 20 53 22
rect 31 18 35 19
rect 122 21 126 42
rect 53 17 57 18
rect 62 17 63 21
rect 67 17 89 21
rect 93 17 121 21
rect 125 17 126 21
rect 41 13 42 17
rect 46 13 47 17
rect 41 12 47 13
rect -2 8 3 12
rect 7 8 108 12
rect 112 8 130 12
rect -2 2 130 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 122 2
rect 126 -2 130 2
<< ntransistor >>
rect 10 11 12 24
rect 17 11 19 24
rect 27 11 29 24
rect 37 16 39 29
rect 49 12 51 23
rect 69 16 71 30
rect 79 16 81 30
rect 101 19 103 30
rect 117 16 119 27
<< ptransistor >>
rect 9 42 11 70
rect 19 42 21 70
rect 29 42 31 70
rect 39 52 41 70
rect 49 52 51 62
rect 72 42 74 70
rect 79 42 81 70
rect 89 42 91 70
rect 107 42 109 70
rect 117 42 119 70
<< polycontact >>
rect 43 44 47 48
rect 10 34 14 38
rect 20 34 24 38
rect 58 38 62 42
rect 70 34 74 38
rect 50 28 54 32
rect 90 34 94 38
rect 114 34 118 38
rect 89 17 93 21
<< ndcontact >>
rect 3 8 7 12
rect 21 18 25 22
rect 31 19 35 23
rect 42 13 46 17
rect 53 18 57 22
rect 63 17 67 21
rect 73 25 77 29
rect 83 25 87 29
rect 95 25 99 29
rect 121 17 125 21
rect 108 8 112 12
<< pdcontact >>
rect 3 59 7 63
rect 13 51 17 55
rect 23 43 27 47
rect 33 65 37 69
rect 33 58 37 62
rect 43 54 47 58
rect 53 57 57 61
rect 66 58 70 62
rect 66 51 70 55
rect 83 59 87 63
rect 83 52 87 56
rect 93 60 97 64
rect 93 53 97 57
rect 101 43 105 47
rect 111 65 115 69
rect 111 58 115 62
rect 121 50 125 54
rect 121 43 125 47
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
rect 90 -2 94 2
rect 98 -2 102 2
rect 106 -2 110 2
rect 114 -2 118 2
rect 122 -2 126 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
rect 90 78 94 82
rect 98 78 102 82
rect 106 78 110 82
rect 114 78 118 82
rect 122 78 126 82
<< psubstratepdiff >>
rect 0 2 128 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 122 2
rect 126 -2 128 2
rect 0 -3 128 -2
<< nsubstratendiff >>
rect 0 82 128 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect 118 78 122 82
rect 126 78 128 82
rect 0 77 128 78
<< labels >>
rlabel ntransistor 11 22 11 22 6 zn
rlabel polycontact 22 36 22 36 6 cn
rlabel polycontact 60 40 60 40 6 iz
rlabel ptransistor 73 53 73 53 6 bn
rlabel polycontact 91 19 91 19 6 an
rlabel metal1 20 20 20 20 6 z
rlabel metal1 12 20 12 20 6 z
rlabel polycontact 12 36 12 36 6 zn
rlabel metal1 4 40 4 40 6 z
rlabel metal1 12 52 12 52 6 z
rlabel metal1 33 24 33 24 6 zn
rlabel metal1 19 45 19 45 6 zn
rlabel metal1 31 36 31 36 6 cn
rlabel metal1 44 44 44 44 6 c
rlabel metal1 14 61 14 61 6 cn
rlabel pdcontact 45 55 45 55 6 cn
rlabel metal1 64 6 64 6 6 vss
rlabel metal1 48 22 48 22 6 cn
rlabel metal1 52 40 52 40 6 c
rlabel polycontact 61 40 61 40 6 iz
rlabel metal1 64 74 64 74 6 vdd
rlabel metal1 69 27 69 27 6 iz
rlabel metal1 92 27 92 27 6 bn
rlabel metal1 77 36 77 36 6 bn
rlabel metal1 92 40 92 40 6 b
rlabel metal1 84 44 84 44 6 b
rlabel metal1 85 57 85 57 6 iz
rlabel metal1 95 57 95 57 6 an
rlabel metal1 94 19 94 19 6 an
rlabel metal1 108 28 108 28 6 a
rlabel pdcontact 102 45 102 45 6 bn
rlabel polycontact 116 36 116 36 6 a
rlabel metal1 124 36 124 36 6 an
<< end >>
