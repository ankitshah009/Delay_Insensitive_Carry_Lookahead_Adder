magic
tech scmos
timestamp 1179384981
<< checkpaint >>
rect -22 -25 78 105
<< ab >>
rect 0 0 56 80
<< pwell >>
rect -4 -7 60 36
<< nwell >>
rect -4 36 60 87
<< polysilicon >>
rect 9 65 11 70
rect 19 65 21 70
rect 29 65 31 70
rect 39 62 41 66
rect 9 42 11 45
rect 19 42 21 45
rect 9 41 21 42
rect 9 37 16 41
rect 20 37 21 41
rect 29 39 31 45
rect 9 36 21 37
rect 25 38 31 39
rect 9 30 11 36
rect 25 34 26 38
rect 30 34 31 38
rect 39 39 41 42
rect 39 38 47 39
rect 39 35 42 38
rect 25 33 31 34
rect 35 34 42 35
rect 46 34 47 38
rect 35 33 47 34
rect 28 30 30 33
rect 35 30 37 33
rect 9 6 11 10
rect 28 8 30 13
rect 35 8 37 13
<< ndiffusion >>
rect 2 29 9 30
rect 2 25 3 29
rect 7 25 9 29
rect 2 22 9 25
rect 2 18 3 22
rect 7 18 9 22
rect 2 17 9 18
rect 4 10 9 17
rect 11 22 28 30
rect 11 18 14 22
rect 18 18 28 22
rect 11 15 28 18
rect 11 11 14 15
rect 18 13 28 15
rect 30 13 35 30
rect 37 23 42 30
rect 37 22 44 23
rect 37 18 39 22
rect 43 18 44 22
rect 37 17 44 18
rect 37 13 42 17
rect 18 11 26 13
rect 11 10 26 11
<< pdiffusion >>
rect 2 64 9 65
rect 2 60 3 64
rect 7 60 9 64
rect 2 45 9 60
rect 11 62 19 65
rect 11 58 13 62
rect 17 58 19 62
rect 11 55 19 58
rect 11 51 13 55
rect 17 51 19 55
rect 11 45 19 51
rect 21 64 29 65
rect 21 60 23 64
rect 27 60 29 64
rect 21 45 29 60
rect 31 62 36 65
rect 31 61 39 62
rect 31 57 33 61
rect 37 57 39 61
rect 31 54 39 57
rect 31 50 33 54
rect 37 50 39 54
rect 31 45 39 50
rect 34 42 39 45
rect 41 61 48 62
rect 41 57 43 61
rect 47 57 48 61
rect 41 54 48 57
rect 41 50 43 54
rect 47 50 48 54
rect 41 42 48 50
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect -2 68 58 78
rect 3 64 7 68
rect 23 64 27 68
rect 3 59 7 60
rect 13 62 17 63
rect 23 59 27 60
rect 33 61 38 62
rect 13 55 17 58
rect 2 51 13 55
rect 37 57 38 61
rect 33 54 38 57
rect 2 50 17 51
rect 23 50 33 54
rect 37 50 38 54
rect 42 61 48 68
rect 42 57 43 61
rect 47 57 48 61
rect 42 54 48 57
rect 42 50 43 54
rect 47 50 48 54
rect 2 30 6 50
rect 23 46 27 50
rect 16 42 27 46
rect 33 42 47 46
rect 16 41 20 42
rect 41 38 47 42
rect 16 30 20 37
rect 25 34 26 38
rect 30 34 37 38
rect 41 34 42 38
rect 46 34 47 38
rect 33 30 37 34
rect 2 29 7 30
rect 2 25 3 29
rect 16 26 28 30
rect 33 26 47 30
rect 2 22 7 25
rect 24 22 28 26
rect 2 18 3 22
rect 2 17 7 18
rect 13 18 14 22
rect 18 18 19 22
rect 24 18 39 22
rect 43 18 44 22
rect 13 15 19 18
rect 13 12 14 15
rect -2 11 14 12
rect 18 12 19 15
rect 18 11 58 12
rect -2 2 58 11
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
<< ntransistor >>
rect 9 10 11 30
rect 28 13 30 30
rect 35 13 37 30
<< ptransistor >>
rect 9 45 11 65
rect 19 45 21 65
rect 29 45 31 65
rect 39 42 41 62
<< polycontact >>
rect 16 37 20 41
rect 26 34 30 38
rect 42 34 46 38
<< ndcontact >>
rect 3 25 7 29
rect 3 18 7 22
rect 14 18 18 22
rect 14 11 18 15
rect 39 18 43 22
<< pdcontact >>
rect 3 60 7 64
rect 13 58 17 62
rect 13 51 17 55
rect 23 60 27 64
rect 33 57 37 61
rect 33 50 37 54
rect 43 57 47 61
rect 43 50 47 54
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
<< psubstratepdiff >>
rect 0 2 56 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 56 2
rect 0 -3 56 -2
<< nsubstratendiff >>
rect 0 82 56 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 56 82
rect 0 77 56 78
<< labels >>
rlabel metal1 4 36 4 36 6 z
rlabel metal1 18 36 18 36 6 zn
rlabel metal1 12 52 12 52 6 z
rlabel metal1 28 6 28 6 6 vss
rlabel polycontact 28 36 28 36 6 a
rlabel metal1 36 28 36 28 6 a
rlabel metal1 36 44 36 44 6 b
rlabel metal1 30 52 30 52 6 zn
rlabel metal1 35 56 35 56 6 zn
rlabel metal1 28 74 28 74 6 vdd
rlabel metal1 34 20 34 20 6 zn
rlabel metal1 44 28 44 28 6 a
rlabel metal1 44 40 44 40 6 b
<< end >>
