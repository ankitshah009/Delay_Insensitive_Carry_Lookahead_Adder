magic
tech scmos
timestamp 1179386476
<< checkpaint >>
rect -22 -22 78 94
<< ab >>
rect 0 0 56 72
<< pwell >>
rect -4 -4 60 32
<< nwell >>
rect -4 32 60 76
<< polysilicon >>
rect 9 66 11 70
rect 19 66 21 70
rect 30 66 32 70
rect 40 66 42 70
rect 9 35 11 38
rect 19 35 21 38
rect 30 35 32 38
rect 9 34 15 35
rect 9 30 10 34
rect 14 30 15 34
rect 9 29 15 30
rect 19 34 32 35
rect 19 30 26 34
rect 30 30 32 34
rect 40 35 42 38
rect 40 34 47 35
rect 40 31 42 34
rect 19 29 32 30
rect 13 25 15 29
rect 20 25 22 29
rect 30 25 32 29
rect 37 30 42 31
rect 46 30 47 34
rect 37 29 47 30
rect 37 25 39 29
rect 13 2 15 7
rect 20 2 22 7
rect 30 2 32 7
rect 37 2 39 7
<< ndiffusion >>
rect 4 11 13 25
rect 4 7 6 11
rect 10 7 13 11
rect 15 7 20 25
rect 22 18 30 25
rect 22 14 24 18
rect 28 14 30 18
rect 22 7 30 14
rect 32 7 37 25
rect 39 19 47 25
rect 39 15 41 19
rect 45 15 47 19
rect 39 12 47 15
rect 39 8 41 12
rect 45 8 47 12
rect 39 7 47 8
rect 4 5 11 7
<< pdiffusion >>
rect 2 65 9 66
rect 2 61 3 65
rect 7 61 9 65
rect 2 57 9 61
rect 2 53 3 57
rect 7 53 9 57
rect 2 38 9 53
rect 11 50 19 66
rect 11 46 13 50
rect 17 46 19 50
rect 11 43 19 46
rect 11 39 13 43
rect 17 39 19 43
rect 11 38 19 39
rect 21 65 30 66
rect 21 61 23 65
rect 27 61 30 65
rect 21 58 30 61
rect 21 54 23 58
rect 27 54 30 58
rect 21 38 30 54
rect 32 57 40 66
rect 32 53 34 57
rect 38 53 40 57
rect 32 50 40 53
rect 32 46 34 50
rect 38 46 40 50
rect 32 38 40 46
rect 42 65 50 66
rect 42 61 44 65
rect 48 61 50 65
rect 42 58 50 61
rect 42 54 44 58
rect 48 54 50 58
rect 42 38 50 54
<< metal1 >>
rect -2 65 58 72
rect -2 64 3 65
rect 7 64 23 65
rect 3 57 7 61
rect 22 61 23 64
rect 27 64 44 65
rect 27 61 28 64
rect 22 58 28 61
rect 43 61 44 64
rect 48 64 58 65
rect 48 61 49 64
rect 22 54 23 58
rect 27 54 28 58
rect 34 57 39 59
rect 3 52 7 53
rect 38 53 39 57
rect 43 58 49 61
rect 43 54 44 58
rect 48 54 49 58
rect 34 50 39 53
rect 12 46 13 50
rect 17 46 34 50
rect 38 46 39 50
rect 12 43 18 46
rect 2 39 13 43
rect 17 39 18 43
rect 2 18 6 39
rect 25 38 39 42
rect 10 34 14 35
rect 25 34 31 38
rect 25 30 26 34
rect 30 30 31 34
rect 41 30 42 34
rect 46 30 47 34
rect 10 26 14 30
rect 41 26 47 30
rect 10 22 47 26
rect 2 14 24 18
rect 28 14 31 18
rect 40 15 41 19
rect 45 15 46 19
rect 40 12 46 15
rect 5 8 6 11
rect -2 7 6 8
rect 10 8 11 11
rect 40 8 41 12
rect 45 8 46 12
rect 10 7 58 8
rect -2 0 58 7
<< ntransistor >>
rect 13 7 15 25
rect 20 7 22 25
rect 30 7 32 25
rect 37 7 39 25
<< ptransistor >>
rect 9 38 11 66
rect 19 38 21 66
rect 30 38 32 66
rect 40 38 42 66
<< polycontact >>
rect 10 30 14 34
rect 26 30 30 34
rect 42 30 46 34
<< ndcontact >>
rect 6 7 10 11
rect 24 14 28 18
rect 41 15 45 19
rect 41 8 45 12
<< pdcontact >>
rect 3 61 7 65
rect 3 53 7 57
rect 13 46 17 50
rect 13 39 17 43
rect 23 61 27 65
rect 23 54 27 58
rect 34 53 38 57
rect 34 46 38 50
rect 44 61 48 65
rect 44 54 48 58
<< labels >>
rlabel metal1 4 32 4 32 6 z
rlabel metal1 20 16 20 16 6 z
rlabel metal1 12 16 12 16 6 z
rlabel polycontact 12 32 12 32 6 a
rlabel metal1 20 24 20 24 6 a
rlabel metal1 20 48 20 48 6 z
rlabel metal1 28 4 28 4 6 vss
rlabel metal1 28 16 28 16 6 z
rlabel metal1 28 24 28 24 6 a
rlabel metal1 36 24 36 24 6 a
rlabel metal1 36 40 36 40 6 b
rlabel metal1 28 36 28 36 6 b
rlabel metal1 28 48 28 48 6 z
rlabel metal1 36 52 36 52 6 z
rlabel metal1 28 68 28 68 6 vdd
rlabel metal1 44 28 44 28 6 a
<< end >>
