magic
tech scmos
timestamp 1179386223
<< checkpaint >>
rect -22 -22 62 94
<< ab >>
rect 0 0 40 72
<< pwell >>
rect -4 -4 44 32
<< nwell >>
rect -4 32 44 76
<< polysilicon >>
rect 10 59 16 60
rect 10 55 11 59
rect 15 55 16 59
rect 10 54 16 55
rect 10 52 12 54
rect 9 49 12 52
rect 29 51 31 56
rect 9 46 11 49
rect 19 46 21 50
rect 9 26 11 38
rect 19 35 21 38
rect 16 34 23 35
rect 16 30 18 34
rect 22 30 23 34
rect 16 29 23 30
rect 16 26 18 29
rect 29 27 31 41
rect 28 26 34 27
rect 9 14 11 19
rect 16 14 18 19
rect 28 22 29 26
rect 33 22 34 26
rect 28 21 34 22
rect 28 18 30 21
rect 28 7 30 12
<< ndiffusion >>
rect 2 25 9 26
rect 2 21 3 25
rect 7 21 9 25
rect 2 19 9 21
rect 11 19 16 26
rect 18 19 26 26
rect 20 18 26 19
rect 20 12 28 18
rect 30 17 37 18
rect 30 13 32 17
rect 36 13 37 17
rect 30 12 37 13
rect 20 8 26 12
rect 20 4 21 8
rect 25 4 26 8
rect 20 3 26 4
<< pdiffusion >>
rect 2 68 8 69
rect 2 64 3 68
rect 7 64 8 68
rect 2 54 8 64
rect 21 57 27 58
rect 2 46 7 54
rect 21 53 22 57
rect 26 53 27 57
rect 21 52 27 53
rect 23 51 27 52
rect 23 46 29 51
rect 2 38 9 46
rect 11 43 19 46
rect 11 39 13 43
rect 17 39 19 43
rect 11 38 19 39
rect 21 41 29 46
rect 31 50 38 51
rect 31 46 33 50
rect 37 46 38 50
rect 31 45 38 46
rect 31 41 36 45
rect 21 38 27 41
<< metal1 >>
rect -2 68 42 72
rect -2 64 3 68
rect 7 64 13 68
rect 17 64 32 68
rect 36 64 42 68
rect 2 55 11 59
rect 15 55 16 59
rect 2 53 16 55
rect 21 57 27 64
rect 21 53 22 57
rect 26 53 27 57
rect 2 37 6 53
rect 26 46 33 50
rect 37 46 38 50
rect 10 39 13 43
rect 17 39 23 43
rect 10 38 23 39
rect 10 27 14 38
rect 26 35 30 46
rect 2 25 14 27
rect 2 21 3 25
rect 7 21 14 25
rect 18 34 30 35
rect 22 31 30 34
rect 18 17 22 30
rect 34 27 38 43
rect 26 26 38 27
rect 26 22 29 26
rect 33 22 38 26
rect 26 21 38 22
rect 18 13 32 17
rect 36 13 37 17
rect -2 4 4 8
rect 8 4 11 8
rect 15 4 21 8
rect 25 4 42 8
rect -2 0 42 4
<< ntransistor >>
rect 9 19 11 26
rect 16 19 18 26
rect 28 12 30 18
<< ptransistor >>
rect 9 38 11 46
rect 19 38 21 46
rect 29 41 31 51
<< polycontact >>
rect 11 55 15 59
rect 18 30 22 34
rect 29 22 33 26
<< ndcontact >>
rect 3 21 7 25
rect 32 13 36 17
rect 21 4 25 8
<< pdcontact >>
rect 3 64 7 68
rect 22 53 26 57
rect 13 39 17 43
rect 33 46 37 50
<< psubstratepcontact >>
rect 4 4 8 8
rect 11 4 15 8
<< nsubstratencontact >>
rect 13 64 17 68
rect 32 64 36 68
<< psubstratepdiff >>
rect 3 8 16 11
rect 3 4 4 8
rect 8 4 11 8
rect 15 4 16 8
rect 3 3 16 4
<< nsubstratendiff >>
rect 12 68 37 69
rect 12 64 13 68
rect 17 64 32 68
rect 36 64 37 68
rect 12 63 37 64
<< labels >>
rlabel ptransistor 20 39 20 39 6 an
rlabel ndcontact 4 24 4 24 6 z
rlabel metal1 4 48 4 48 6 b
rlabel metal1 12 32 12 32 6 z
rlabel polycontact 12 56 12 56 6 b
rlabel metal1 20 4 20 4 6 vss
rlabel metal1 20 24 20 24 6 an
rlabel metal1 28 24 28 24 6 a
rlabel metal1 20 40 20 40 6 z
rlabel metal1 20 68 20 68 6 vdd
rlabel metal1 27 15 27 15 6 an
rlabel metal1 36 32 36 32 6 a
rlabel metal1 32 48 32 48 6 an
<< end >>
