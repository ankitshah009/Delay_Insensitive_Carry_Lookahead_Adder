magic
tech scmos
timestamp 1185039019
<< checkpaint >>
rect -22 -24 142 124
<< ab >>
rect 0 0 120 100
<< pwell >>
rect -2 -4 122 49
<< nwell >>
rect -2 49 122 104
<< polysilicon >>
rect 93 95 95 98
rect 105 95 107 98
rect 11 85 13 88
rect 23 85 25 88
rect 31 85 33 88
rect 47 85 49 88
rect 55 85 57 88
rect 67 85 69 88
rect 11 41 13 65
rect 23 63 25 65
rect 17 62 25 63
rect 17 58 18 62
rect 22 61 25 62
rect 22 58 23 61
rect 17 57 23 58
rect 31 43 33 65
rect 47 57 49 65
rect 55 63 57 65
rect 55 62 63 63
rect 55 61 58 62
rect 57 58 58 61
rect 62 58 63 62
rect 57 57 63 58
rect 47 56 53 57
rect 47 52 48 56
rect 52 52 53 56
rect 47 51 53 52
rect 37 50 43 51
rect 37 46 38 50
rect 42 47 43 50
rect 67 47 69 65
rect 73 52 79 53
rect 73 48 74 52
rect 78 51 79 52
rect 93 51 95 55
rect 105 51 107 55
rect 78 49 107 51
rect 78 48 79 49
rect 73 47 79 48
rect 42 46 69 47
rect 37 45 69 46
rect 27 42 33 43
rect 27 41 28 42
rect 11 39 28 41
rect 11 15 13 39
rect 27 38 28 39
rect 32 41 33 42
rect 32 39 49 41
rect 32 38 33 39
rect 27 37 33 38
rect 17 32 23 33
rect 17 28 18 32
rect 22 29 23 32
rect 22 28 25 29
rect 17 27 25 28
rect 23 15 25 27
rect 29 22 35 23
rect 29 18 30 22
rect 34 18 35 22
rect 29 17 35 18
rect 31 15 33 17
rect 47 15 49 39
rect 57 32 63 33
rect 57 29 58 32
rect 55 28 58 29
rect 62 28 63 32
rect 55 27 63 28
rect 55 15 57 27
rect 67 15 69 45
rect 93 25 95 49
rect 105 25 107 49
rect 11 2 13 5
rect 23 2 25 5
rect 31 2 33 5
rect 47 2 49 5
rect 55 2 57 5
rect 67 2 69 5
rect 93 2 95 5
rect 105 2 107 5
<< ndiffusion >>
rect 3 22 9 23
rect 3 18 4 22
rect 8 18 9 22
rect 3 15 9 18
rect 37 32 45 33
rect 37 28 38 32
rect 42 28 45 32
rect 37 15 45 28
rect 71 22 77 23
rect 71 18 72 22
rect 76 18 77 22
rect 71 15 77 18
rect 3 5 11 15
rect 13 12 23 15
rect 13 8 16 12
rect 20 8 23 12
rect 13 5 23 8
rect 25 5 31 15
rect 33 5 47 15
rect 49 5 55 15
rect 57 12 67 15
rect 57 8 60 12
rect 64 8 67 12
rect 57 5 67 8
rect 69 5 77 15
rect 85 22 93 25
rect 85 18 86 22
rect 90 18 93 22
rect 85 12 93 18
rect 85 8 86 12
rect 90 8 93 12
rect 85 5 93 8
rect 95 22 105 25
rect 95 18 98 22
rect 102 18 105 22
rect 95 5 105 18
rect 107 22 115 25
rect 107 18 110 22
rect 114 18 115 22
rect 107 12 115 18
rect 107 8 110 12
rect 114 8 115 12
rect 107 5 115 8
<< pdiffusion >>
rect 15 92 21 93
rect 15 88 16 92
rect 20 88 21 92
rect 59 92 65 93
rect 59 88 60 92
rect 64 88 65 92
rect 85 92 93 95
rect 85 88 86 92
rect 90 88 93 92
rect 15 85 21 88
rect 59 85 65 88
rect 3 82 11 85
rect 3 78 4 82
rect 8 78 11 82
rect 3 72 11 78
rect 3 68 4 72
rect 8 68 11 72
rect 3 65 11 68
rect 13 65 23 85
rect 25 65 31 85
rect 33 82 47 85
rect 33 78 38 82
rect 42 78 47 82
rect 33 72 47 78
rect 33 68 38 72
rect 42 68 47 72
rect 33 65 47 68
rect 49 65 55 85
rect 57 65 67 85
rect 69 82 77 85
rect 69 78 72 82
rect 76 78 77 82
rect 69 70 77 78
rect 69 66 72 70
rect 76 66 77 70
rect 69 65 77 66
rect 85 82 93 88
rect 85 78 86 82
rect 90 78 93 82
rect 85 72 93 78
rect 85 68 86 72
rect 90 68 93 72
rect 85 62 93 68
rect 85 58 86 62
rect 90 58 93 62
rect 85 55 93 58
rect 95 82 105 95
rect 95 78 98 82
rect 102 78 105 82
rect 95 72 105 78
rect 95 68 98 72
rect 102 68 105 72
rect 95 62 105 68
rect 95 58 98 62
rect 102 58 105 62
rect 95 55 105 58
rect 107 92 115 95
rect 107 88 110 92
rect 114 88 115 92
rect 107 82 115 88
rect 107 78 110 82
rect 114 78 115 82
rect 107 72 115 78
rect 107 68 110 72
rect 114 68 115 72
rect 107 62 115 68
rect 107 58 110 62
rect 114 58 115 62
rect 107 55 115 58
<< metal1 >>
rect -2 96 122 101
rect -2 92 28 96
rect 32 92 38 96
rect 42 92 48 96
rect 52 92 122 96
rect -2 88 16 92
rect 20 88 60 92
rect 64 88 86 92
rect 90 88 110 92
rect 114 88 122 92
rect -2 87 122 88
rect 3 82 9 83
rect 37 82 43 83
rect 71 82 77 83
rect 3 78 4 82
rect 8 78 9 82
rect 3 77 9 78
rect 4 73 8 77
rect 3 72 9 73
rect 3 68 4 72
rect 8 68 9 72
rect 3 67 9 68
rect 4 23 8 67
rect 17 62 23 82
rect 17 58 18 62
rect 22 58 23 62
rect 17 32 23 58
rect 17 28 18 32
rect 22 28 23 32
rect 27 42 33 82
rect 37 78 38 82
rect 42 78 43 82
rect 37 77 43 78
rect 38 73 42 77
rect 37 72 43 73
rect 37 68 38 72
rect 42 68 43 72
rect 37 67 43 68
rect 38 51 42 67
rect 57 62 63 82
rect 71 78 72 82
rect 76 78 77 82
rect 71 77 77 78
rect 85 82 91 87
rect 85 78 86 82
rect 90 78 91 82
rect 72 71 76 77
rect 85 72 91 78
rect 71 70 77 71
rect 71 66 72 70
rect 76 66 77 70
rect 71 65 77 66
rect 85 68 86 72
rect 90 68 91 72
rect 57 58 58 62
rect 62 58 63 62
rect 47 56 53 57
rect 47 52 48 56
rect 52 52 53 56
rect 47 51 53 52
rect 37 50 43 51
rect 37 46 38 50
rect 42 46 43 50
rect 37 45 43 46
rect 27 38 28 42
rect 32 38 33 42
rect 27 28 33 38
rect 38 33 42 45
rect 37 32 43 33
rect 37 28 38 32
rect 42 28 43 32
rect 17 27 23 28
rect 37 27 43 28
rect 3 22 9 23
rect 29 22 35 23
rect 48 22 52 51
rect 3 18 4 22
rect 8 18 30 22
rect 34 18 52 22
rect 57 32 63 58
rect 57 28 58 32
rect 62 28 63 32
rect 57 18 63 28
rect 72 53 76 65
rect 85 62 91 68
rect 85 58 86 62
rect 90 58 91 62
rect 85 57 91 58
rect 97 82 103 83
rect 97 78 98 82
rect 102 78 103 82
rect 97 72 103 78
rect 97 68 98 72
rect 102 68 103 72
rect 97 62 103 68
rect 97 58 98 62
rect 102 58 103 62
rect 72 52 79 53
rect 72 48 74 52
rect 78 48 79 52
rect 72 47 79 48
rect 72 23 76 47
rect 71 22 77 23
rect 71 18 72 22
rect 76 18 77 22
rect 3 17 9 18
rect 29 17 35 18
rect 71 17 77 18
rect 85 22 91 23
rect 85 18 86 22
rect 90 18 91 22
rect 85 13 91 18
rect 97 22 103 58
rect 109 82 115 87
rect 109 78 110 82
rect 114 78 115 82
rect 109 72 115 78
rect 109 68 110 72
rect 114 68 115 72
rect 109 62 115 68
rect 109 58 110 62
rect 114 58 115 62
rect 109 57 115 58
rect 97 18 98 22
rect 102 18 103 22
rect 97 17 103 18
rect 109 22 115 23
rect 109 18 110 22
rect 114 18 115 22
rect 109 13 115 18
rect -2 12 122 13
rect -2 8 16 12
rect 20 8 60 12
rect 64 8 86 12
rect 90 8 110 12
rect 114 8 122 12
rect -2 -1 122 8
<< ntransistor >>
rect 11 5 13 15
rect 23 5 25 15
rect 31 5 33 15
rect 47 5 49 15
rect 55 5 57 15
rect 67 5 69 15
rect 93 5 95 25
rect 105 5 107 25
<< ptransistor >>
rect 11 65 13 85
rect 23 65 25 85
rect 31 65 33 85
rect 47 65 49 85
rect 55 65 57 85
rect 67 65 69 85
rect 93 55 95 95
rect 105 55 107 95
<< polycontact >>
rect 18 58 22 62
rect 58 58 62 62
rect 48 52 52 56
rect 38 46 42 50
rect 74 48 78 52
rect 28 38 32 42
rect 18 28 22 32
rect 30 18 34 22
rect 58 28 62 32
<< ndcontact >>
rect 4 18 8 22
rect 38 28 42 32
rect 72 18 76 22
rect 16 8 20 12
rect 60 8 64 12
rect 86 18 90 22
rect 86 8 90 12
rect 98 18 102 22
rect 110 18 114 22
rect 110 8 114 12
<< pdcontact >>
rect 16 88 20 92
rect 60 88 64 92
rect 86 88 90 92
rect 4 78 8 82
rect 4 68 8 72
rect 38 78 42 82
rect 38 68 42 72
rect 72 78 76 82
rect 72 66 76 70
rect 86 78 90 82
rect 86 68 90 72
rect 86 58 90 62
rect 98 78 102 82
rect 98 68 102 72
rect 98 58 102 62
rect 110 88 114 92
rect 110 78 114 82
rect 110 68 114 72
rect 110 58 114 62
<< nsubstratencontact >>
rect 28 92 32 96
rect 38 92 42 96
rect 48 92 52 96
<< nsubstratendiff >>
rect 27 96 53 97
rect 27 92 28 96
rect 32 92 38 96
rect 42 92 48 96
rect 52 92 53 96
rect 27 91 53 92
<< labels >>
rlabel metal1 20 55 20 55 6 i0
rlabel metal1 20 55 20 55 6 i0
rlabel metal1 30 55 30 55 6 cmd
rlabel metal1 30 55 30 55 6 cmd
rlabel metal1 60 6 60 6 6 vss
rlabel metal1 60 6 60 6 6 vss
rlabel metal1 60 50 60 50 6 i1
rlabel metal1 60 50 60 50 6 i1
rlabel metal1 60 94 60 94 6 vdd
rlabel metal1 60 94 60 94 6 vdd
rlabel metal1 100 50 100 50 6 nq
rlabel metal1 100 50 100 50 6 nq
<< end >>
