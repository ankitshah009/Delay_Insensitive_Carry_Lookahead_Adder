magic
tech scmos
timestamp 1179387602
<< checkpaint >>
rect -22 -22 118 94
<< ab >>
rect 0 0 96 72
<< pwell >>
rect -4 -4 100 32
<< nwell >>
rect -4 32 100 76
<< polysilicon >>
rect 9 66 11 70
rect 19 66 21 70
rect 29 65 31 70
rect 36 68 64 70
rect 36 65 38 68
rect 55 60 57 64
rect 62 60 64 68
rect 74 66 76 70
rect 9 35 11 38
rect 19 35 21 38
rect 9 34 15 35
rect 9 30 10 34
rect 14 30 15 34
rect 9 29 15 30
rect 19 34 25 35
rect 19 30 20 34
rect 24 30 25 34
rect 19 29 25 30
rect 29 30 31 38
rect 36 34 38 38
rect 55 35 57 38
rect 51 34 57 35
rect 51 30 52 34
rect 56 30 57 34
rect 10 20 12 29
rect 19 25 21 29
rect 29 28 57 30
rect 62 34 64 38
rect 74 35 76 38
rect 74 34 81 35
rect 62 33 70 34
rect 62 29 65 33
rect 69 29 70 33
rect 62 28 70 29
rect 74 30 76 34
rect 80 30 81 34
rect 74 29 81 30
rect 17 23 21 25
rect 37 24 39 28
rect 62 25 64 28
rect 74 25 76 29
rect 17 20 19 23
rect 27 20 29 24
rect 37 8 39 12
rect 62 8 64 12
rect 10 2 12 7
rect 17 2 19 7
rect 27 4 29 7
rect 74 4 76 12
rect 27 2 76 4
<< ndiffusion >>
rect 55 24 62 25
rect 32 20 37 24
rect 2 8 10 20
rect 2 4 3 8
rect 7 7 10 8
rect 12 7 17 20
rect 19 18 27 20
rect 19 14 21 18
rect 25 14 27 18
rect 19 7 27 14
rect 29 19 37 20
rect 29 15 31 19
rect 35 15 37 19
rect 29 12 37 15
rect 39 17 46 24
rect 39 13 41 17
rect 45 13 46 17
rect 39 12 46 13
rect 55 20 56 24
rect 60 20 62 24
rect 55 17 62 20
rect 55 13 56 17
rect 60 13 62 17
rect 55 12 62 13
rect 64 17 74 25
rect 64 13 68 17
rect 72 13 74 17
rect 64 12 74 13
rect 76 18 81 25
rect 76 17 83 18
rect 76 13 78 17
rect 82 13 83 17
rect 76 12 83 13
rect 29 7 34 12
rect 7 4 8 7
rect 2 3 8 4
<< pdiffusion >>
rect 4 60 9 66
rect 2 59 9 60
rect 2 55 3 59
rect 7 55 9 59
rect 2 54 9 55
rect 4 38 9 54
rect 11 50 19 66
rect 11 46 13 50
rect 17 46 19 50
rect 11 38 19 46
rect 21 65 26 66
rect 21 50 29 65
rect 21 46 23 50
rect 27 46 29 50
rect 21 43 29 46
rect 21 39 23 43
rect 27 39 29 43
rect 21 38 29 39
rect 31 38 36 65
rect 38 64 46 65
rect 38 60 40 64
rect 44 60 46 64
rect 66 65 74 66
rect 66 61 68 65
rect 72 61 74 65
rect 66 60 74 61
rect 38 50 46 60
rect 38 38 44 50
rect 50 44 55 60
rect 48 43 55 44
rect 48 39 49 43
rect 53 39 55 43
rect 48 38 55 39
rect 57 38 62 60
rect 64 38 74 60
rect 76 59 81 66
rect 76 58 83 59
rect 76 54 78 58
rect 82 54 83 58
rect 76 53 83 54
rect 76 38 81 53
<< metal1 >>
rect -2 68 98 72
rect -2 65 88 68
rect -2 64 68 65
rect 67 61 68 64
rect 72 64 88 65
rect 92 64 98 68
rect 72 61 73 64
rect 40 59 44 60
rect 2 55 3 59
rect 7 55 36 59
rect 50 55 78 58
rect 32 54 78 55
rect 82 54 89 58
rect 32 51 54 54
rect 23 50 27 51
rect 2 46 13 50
rect 17 46 18 50
rect 2 18 6 46
rect 23 43 27 46
rect 10 39 23 42
rect 10 38 27 39
rect 10 34 14 38
rect 32 34 36 51
rect 19 30 20 34
rect 24 30 36 34
rect 42 39 49 43
rect 53 39 54 43
rect 10 26 14 30
rect 10 25 35 26
rect 42 25 46 39
rect 58 35 62 51
rect 66 45 78 51
rect 50 34 62 35
rect 66 34 70 35
rect 50 30 52 34
rect 56 30 62 34
rect 50 29 62 30
rect 65 33 70 34
rect 69 29 70 33
rect 74 34 78 45
rect 74 30 76 34
rect 80 30 81 34
rect 65 28 70 29
rect 66 26 70 28
rect 10 24 61 25
rect 10 22 56 24
rect 31 21 56 22
rect 31 19 35 21
rect 2 14 21 18
rect 25 14 26 18
rect 55 20 56 21
rect 60 20 61 24
rect 66 21 79 26
rect 55 17 61 20
rect 85 17 89 54
rect 31 14 35 15
rect 40 13 41 17
rect 45 13 46 17
rect 55 13 56 17
rect 60 13 61 17
rect 67 13 68 17
rect 72 13 73 17
rect 77 13 78 17
rect 82 13 89 17
rect 40 8 46 13
rect 67 8 73 13
rect -2 4 3 8
rect 7 4 88 8
rect 92 4 98 8
rect -2 0 98 4
<< ntransistor >>
rect 10 7 12 20
rect 17 7 19 20
rect 27 7 29 20
rect 37 12 39 24
rect 62 12 64 25
rect 74 12 76 25
<< ptransistor >>
rect 9 38 11 66
rect 19 38 21 66
rect 29 38 31 65
rect 36 38 38 65
rect 55 38 57 60
rect 62 38 64 60
rect 74 38 76 66
<< polycontact >>
rect 10 30 14 34
rect 20 30 24 34
rect 52 30 56 34
rect 65 29 69 33
rect 76 30 80 34
<< ndcontact >>
rect 3 4 7 8
rect 21 14 25 18
rect 31 15 35 19
rect 41 13 45 17
rect 56 20 60 24
rect 56 13 60 17
rect 68 13 72 17
rect 78 13 82 17
<< pdcontact >>
rect 3 55 7 59
rect 13 46 17 50
rect 23 46 27 50
rect 23 39 27 43
rect 40 60 44 64
rect 68 61 72 65
rect 49 39 53 43
rect 78 54 82 58
<< psubstratepcontact >>
rect 88 4 92 8
<< nsubstratencontact >>
rect 88 64 92 68
<< psubstratepdiff >>
rect 87 8 93 24
rect 87 4 88 8
rect 92 4 93 8
rect 87 3 93 4
<< nsubstratendiff >>
rect 87 68 93 69
rect 87 64 88 68
rect 92 64 93 68
rect 87 40 93 64
<< labels >>
rlabel polycontact 22 32 22 32 6 bn
rlabel polycontact 12 32 12 32 6 an
rlabel metal1 12 16 12 16 6 z
rlabel metal1 4 32 4 32 6 z
rlabel polycontact 12 32 12 32 6 an
rlabel metal1 12 48 12 48 6 z
rlabel metal1 33 20 33 20 6 an
rlabel metal1 20 16 20 16 6 z
rlabel metal1 27 32 27 32 6 bn
rlabel metal1 25 44 25 44 6 an
rlabel metal1 19 57 19 57 6 bn
rlabel metal1 48 4 48 4 6 vss
rlabel metal1 52 32 52 32 6 a2
rlabel metal1 48 41 48 41 6 an
rlabel metal1 48 68 48 68 6 vdd
rlabel metal1 58 19 58 19 6 an
rlabel metal1 76 24 76 24 6 a1
rlabel metal1 68 28 68 28 6 a1
rlabel metal1 60 40 60 40 6 a2
rlabel metal1 76 44 76 44 6 b
rlabel metal1 68 48 68 48 6 b
rlabel metal1 83 15 83 15 6 bn
rlabel metal1 69 56 69 56 6 bn
<< end >>
