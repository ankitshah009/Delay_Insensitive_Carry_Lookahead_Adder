magic
tech scmos
timestamp 1179386892
<< checkpaint >>
rect -22 -25 110 105
<< ab >>
rect 0 0 88 80
<< pwell >>
rect -4 -7 92 36
<< nwell >>
rect -4 36 92 87
<< polysilicon >>
rect 11 70 13 74
rect 18 70 20 74
rect 25 70 27 74
rect 35 70 37 74
rect 42 70 44 74
rect 49 70 51 74
rect 59 70 61 74
rect 66 70 68 74
rect 73 70 75 74
rect 11 34 13 43
rect 18 40 20 43
rect 25 40 27 43
rect 35 40 37 43
rect 18 38 21 40
rect 25 38 37 40
rect 19 34 21 38
rect 29 34 30 38
rect 34 34 35 38
rect 9 33 15 34
rect 9 29 10 33
rect 14 29 15 33
rect 9 28 15 29
rect 19 33 25 34
rect 19 29 20 33
rect 24 29 25 33
rect 19 28 25 29
rect 29 33 35 34
rect 9 25 11 28
rect 19 25 21 28
rect 29 25 31 33
rect 42 30 44 43
rect 49 40 51 43
rect 59 40 61 43
rect 49 39 62 40
rect 49 38 57 39
rect 56 35 57 38
rect 61 35 62 39
rect 56 34 62 35
rect 66 30 68 43
rect 42 28 68 30
rect 73 31 75 43
rect 73 30 79 31
rect 42 22 48 28
rect 73 26 74 30
rect 78 26 79 30
rect 73 25 79 26
rect 42 18 43 22
rect 47 18 48 22
rect 42 17 48 18
rect 9 6 11 10
rect 19 6 21 10
rect 29 6 31 10
<< ndiffusion >>
rect 4 23 9 25
rect 2 22 9 23
rect 2 18 3 22
rect 7 18 9 22
rect 2 17 9 18
rect 4 10 9 17
rect 11 15 19 25
rect 11 11 13 15
rect 17 11 19 15
rect 11 10 19 11
rect 21 22 29 25
rect 21 18 23 22
rect 27 18 29 22
rect 21 10 29 18
rect 31 22 39 25
rect 31 18 33 22
rect 37 18 39 22
rect 31 15 39 18
rect 31 11 33 15
rect 37 11 39 15
rect 31 10 39 11
<< pdiffusion >>
rect 6 62 11 70
rect 4 61 11 62
rect 4 57 5 61
rect 9 57 11 61
rect 4 54 11 57
rect 4 50 5 54
rect 9 50 11 54
rect 4 49 11 50
rect 6 43 11 49
rect 13 43 18 70
rect 20 43 25 70
rect 27 69 35 70
rect 27 65 29 69
rect 33 65 35 69
rect 27 62 35 65
rect 27 58 29 62
rect 33 58 35 62
rect 27 43 35 58
rect 37 43 42 70
rect 44 43 49 70
rect 51 62 59 70
rect 51 58 53 62
rect 57 58 59 62
rect 51 55 59 58
rect 51 51 53 55
rect 57 51 59 55
rect 51 43 59 51
rect 61 43 66 70
rect 68 43 73 70
rect 75 69 82 70
rect 75 65 77 69
rect 81 65 82 69
rect 75 62 82 65
rect 75 58 77 62
rect 81 58 82 62
rect 75 43 82 58
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect -2 69 90 78
rect -2 68 29 69
rect 28 65 29 68
rect 33 68 77 69
rect 33 65 34 68
rect 28 62 34 65
rect 76 65 77 68
rect 81 68 90 69
rect 81 65 82 68
rect 5 61 9 62
rect 28 58 29 62
rect 33 58 34 62
rect 53 62 57 63
rect 76 62 82 65
rect 76 58 77 62
rect 81 58 82 62
rect 5 55 9 57
rect 2 54 9 55
rect 53 55 57 58
rect 2 50 5 54
rect 9 51 53 54
rect 57 51 63 54
rect 9 50 63 51
rect 2 22 6 50
rect 10 42 63 46
rect 10 33 14 42
rect 57 39 63 42
rect 29 34 30 38
rect 34 34 53 38
rect 61 35 63 39
rect 57 34 63 35
rect 10 28 14 29
rect 20 33 24 34
rect 49 30 53 34
rect 24 29 45 30
rect 20 26 45 29
rect 49 26 74 30
rect 78 26 79 30
rect 41 22 45 26
rect 2 18 3 22
rect 7 18 23 22
rect 27 18 28 22
rect 32 18 33 22
rect 37 18 38 22
rect 41 18 43 22
rect 47 18 55 22
rect 32 15 38 18
rect 12 12 13 15
rect -2 11 13 12
rect 17 12 18 15
rect 32 12 33 15
rect 17 11 33 12
rect 37 12 38 15
rect 37 11 90 12
rect -2 2 90 11
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
<< ntransistor >>
rect 9 10 11 25
rect 19 10 21 25
rect 29 10 31 25
<< ptransistor >>
rect 11 43 13 70
rect 18 43 20 70
rect 25 43 27 70
rect 35 43 37 70
rect 42 43 44 70
rect 49 43 51 70
rect 59 43 61 70
rect 66 43 68 70
rect 73 43 75 70
<< polycontact >>
rect 30 34 34 38
rect 10 29 14 33
rect 20 29 24 33
rect 57 35 61 39
rect 74 26 78 30
rect 43 18 47 22
<< ndcontact >>
rect 3 18 7 22
rect 13 11 17 15
rect 23 18 27 22
rect 33 18 37 22
rect 33 11 37 15
<< pdcontact >>
rect 5 57 9 61
rect 5 50 9 54
rect 29 65 33 69
rect 29 58 33 62
rect 53 58 57 62
rect 53 51 57 55
rect 77 65 81 69
rect 77 58 81 62
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
<< psubstratepdiff >>
rect 0 2 88 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 88 2
rect 0 -3 88 -2
<< nsubstratendiff >>
rect 0 82 88 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 88 82
rect 0 77 88 78
<< labels >>
rlabel metal1 12 20 12 20 6 z
rlabel metal1 4 40 4 40 6 z
rlabel metal1 12 36 12 36 6 c
rlabel metal1 12 52 12 52 6 z
rlabel metal1 20 20 20 20 6 z
rlabel metal1 28 28 28 28 6 b
rlabel metal1 20 44 20 44 6 c
rlabel metal1 28 44 28 44 6 c
rlabel metal1 20 52 20 52 6 z
rlabel metal1 28 52 28 52 6 z
rlabel metal1 44 6 44 6 6 vss
rlabel metal1 36 28 36 28 6 b
rlabel polycontact 44 20 44 20 6 b
rlabel metal1 36 36 36 36 6 a
rlabel metal1 36 44 36 44 6 c
rlabel metal1 44 36 44 36 6 a
rlabel metal1 44 44 44 44 6 c
rlabel metal1 44 52 44 52 6 z
rlabel metal1 36 52 36 52 6 z
rlabel metal1 44 74 44 74 6 vdd
rlabel metal1 52 20 52 20 6 b
rlabel metal1 52 28 52 28 6 a
rlabel metal1 60 28 60 28 6 a
rlabel metal1 68 28 68 28 6 a
rlabel metal1 52 44 52 44 6 c
rlabel metal1 60 40 60 40 6 c
rlabel metal1 60 52 60 52 6 z
rlabel metal1 52 52 52 52 6 z
rlabel polycontact 76 28 76 28 6 a
<< end >>
