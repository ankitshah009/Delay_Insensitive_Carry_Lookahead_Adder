magic
tech scmos
timestamp 1170759784
<< checkpaint >>
rect -22 -26 54 114
<< ab >>
rect 0 0 32 88
<< pwell >>
rect -4 -8 36 40
<< nwell >>
rect -4 40 36 96
<< polysilicon >>
rect 2 77 11 83
rect 9 74 11 77
rect 21 77 30 83
rect 21 74 23 77
rect 9 43 11 46
rect 21 43 23 46
rect 2 42 14 43
rect 2 38 6 42
rect 10 38 14 42
rect 2 37 14 38
rect 18 42 30 43
rect 18 38 19 42
rect 23 38 30 42
rect 18 37 30 38
rect 9 34 11 37
rect 21 34 23 37
rect 9 11 11 14
rect 2 5 11 11
rect 21 11 23 14
rect 21 5 30 11
<< ndiffusion >>
rect 2 26 9 34
rect 2 22 3 26
rect 7 22 9 26
rect 2 19 9 22
rect 2 15 3 19
rect 7 15 9 19
rect 2 14 9 15
rect 11 29 21 34
rect 11 25 14 29
rect 18 25 21 29
rect 11 22 21 25
rect 11 18 14 22
rect 18 18 21 22
rect 11 14 21 18
rect 23 19 30 34
rect 23 15 25 19
rect 29 15 30 19
rect 23 14 30 15
rect 13 2 19 14
<< pdiffusion >>
rect 13 74 19 86
rect 2 73 9 74
rect 2 69 3 73
rect 7 69 9 73
rect 2 66 9 69
rect 2 62 3 66
rect 7 62 9 66
rect 2 46 9 62
rect 11 62 21 74
rect 11 58 14 62
rect 18 58 21 62
rect 11 55 21 58
rect 11 51 14 55
rect 18 51 21 55
rect 11 46 21 51
rect 23 73 30 74
rect 23 69 25 73
rect 29 69 30 73
rect 23 66 30 69
rect 23 62 25 66
rect 29 62 30 66
rect 23 46 30 62
<< metal1 >>
rect -2 86 2 90
rect 10 86 22 90
rect 30 86 34 90
rect 3 82 7 86
rect 3 73 7 78
rect 3 66 7 69
rect 25 82 29 86
rect 25 73 29 78
rect 25 66 29 69
rect 3 61 7 62
rect 14 62 18 63
rect 25 61 29 62
rect 14 55 18 58
rect 6 43 10 55
rect 18 51 30 54
rect 14 50 30 51
rect 6 42 23 43
rect 10 38 19 42
rect 6 37 23 38
rect 6 33 10 37
rect 26 30 30 50
rect 14 29 30 30
rect 3 26 7 27
rect 3 19 7 22
rect 18 26 30 29
rect 14 22 18 25
rect 14 17 18 18
rect 25 19 29 20
rect 3 10 7 15
rect 3 2 7 6
rect 25 10 29 15
rect 25 2 29 6
rect -2 -2 2 2
rect 10 -2 22 2
rect 30 -2 34 2
<< metal2 >>
rect -2 86 6 90
rect 10 86 22 90
rect 26 86 34 90
rect -2 82 34 86
rect -2 78 3 82
rect 7 78 25 82
rect 29 78 34 82
rect -2 76 34 78
rect -2 10 34 12
rect -2 6 3 10
rect 7 6 25 10
rect 29 6 34 10
rect -2 2 34 6
rect -2 -2 6 2
rect 10 -2 22 2
rect 26 -2 34 2
<< ntransistor >>
rect 9 14 11 34
rect 21 14 23 34
<< ptransistor >>
rect 9 46 11 74
rect 21 46 23 74
<< polycontact >>
rect 6 38 10 42
rect 19 38 23 42
<< ndcontact >>
rect 3 22 7 26
rect 3 15 7 19
rect 14 25 18 29
rect 14 18 18 22
rect 25 15 29 19
<< pdcontact >>
rect 3 69 7 73
rect 3 62 7 66
rect 14 58 18 62
rect 14 51 18 55
rect 25 69 29 73
rect 25 62 29 66
<< m2contact >>
rect 6 86 10 90
rect 22 86 26 90
rect 3 78 7 82
rect 25 78 29 82
rect 3 6 7 10
rect 25 6 29 10
rect 6 -2 10 2
rect 22 -2 26 2
<< psubstratepcontact >>
rect 2 -2 6 2
rect 26 -2 30 2
<< nsubstratencontact >>
rect 2 86 6 90
rect 26 86 30 90
<< psubstratepdiff >>
rect 0 2 7 3
rect 25 2 32 3
rect 0 -2 2 2
rect 6 -2 7 2
rect 0 -3 7 -2
rect 25 -2 26 2
rect 30 -2 32 2
rect 25 -3 32 -2
<< nsubstratendiff >>
rect 0 90 7 91
rect 0 86 2 90
rect 6 86 7 90
rect 25 90 32 91
rect 25 86 26 90
rect 30 86 32 90
rect 0 85 7 86
rect 25 85 32 86
<< labels >>
rlabel metal1 8 44 8 44 6 a
rlabel ndcontact 16 20 16 20 6 z
rlabel pdcontact 16 60 16 60 6 z
rlabel metal1 24 28 24 28 6 z
rlabel metal1 24 52 24 52 6 z
rlabel metal2 16 6 16 6 6 vss
rlabel metal2 16 6 16 6 6 vss
rlabel metal2 16 82 16 82 6 vdd
<< end >>
