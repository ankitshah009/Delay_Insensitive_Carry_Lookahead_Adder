.subckt nd2v0x2 a b vdd vss z
*   SPICE3 file   created from nd2v0x2.ext -      technology: scmos
m00 z      b      vdd    vdd p w=24u  l=2.3636u ad=96p      pd=32u      as=180p     ps=63u
m01 vdd    a      z      vdd p w=24u  l=2.3636u ad=180p     pd=63u      as=96p      ps=32u
m02 w1     b      z      vss n w=20u  l=2.3636u ad=50p      pd=25u      as=112p     ps=54u
m03 vss    a      w1     vss n w=20u  l=2.3636u ad=180p     pd=58u      as=50p      ps=25u
C0  b      vdd    0.014f
C1  vss    z      0.080f
C2  vss    b      0.036f
C3  z      b      0.142f
C4  a      vdd    0.035f
C5  vss    w1     0.005f
C6  vss    a      0.024f
C7  w1     b      0.008f
C8  z      a      0.029f
C9  vss    vdd    0.003f
C10 a      b      0.104f
C11 z      vdd    0.186f
C13 z      vss    0.014f
C14 a      vss    0.027f
C15 b      vss    0.017f
.ends
