magic
tech scmos
timestamp 1180600810
<< checkpaint >>
rect -22 -22 132 122
<< ab >>
rect 0 0 110 100
<< pwell >>
rect -4 -4 114 48
<< nwell >>
rect -4 48 114 104
<< polysilicon >>
rect 15 94 17 98
rect 27 85 29 89
rect 39 85 41 89
rect 51 85 53 89
rect 63 85 65 89
rect 77 85 79 89
rect 87 85 89 89
rect 97 85 99 89
rect 15 43 17 55
rect 27 43 29 63
rect 39 43 41 63
rect 51 43 53 63
rect 63 43 65 61
rect 15 42 23 43
rect 15 38 18 42
rect 22 38 23 42
rect 15 37 23 38
rect 27 42 33 43
rect 27 38 28 42
rect 32 38 33 42
rect 27 37 33 38
rect 37 42 43 43
rect 37 38 38 42
rect 42 38 43 42
rect 37 37 43 38
rect 47 42 53 43
rect 47 38 48 42
rect 52 38 53 42
rect 47 37 53 38
rect 57 42 65 43
rect 57 38 58 42
rect 62 38 65 42
rect 77 53 79 56
rect 87 53 89 56
rect 77 52 83 53
rect 77 48 78 52
rect 82 48 83 52
rect 77 47 83 48
rect 87 52 93 53
rect 87 48 88 52
rect 92 48 93 52
rect 87 47 93 48
rect 77 39 79 47
rect 87 39 89 47
rect 57 37 65 38
rect 73 37 79 39
rect 85 37 89 39
rect 97 43 99 55
rect 97 42 103 43
rect 97 38 98 42
rect 102 38 103 42
rect 97 37 103 38
rect 15 34 17 37
rect 29 33 31 37
rect 39 33 41 37
rect 49 33 51 37
rect 61 29 63 37
rect 73 25 75 37
rect 85 25 87 37
rect 97 25 99 37
rect 15 10 17 14
rect 29 13 31 17
rect 39 13 41 17
rect 49 13 51 17
rect 61 13 63 17
rect 73 13 75 17
rect 85 13 87 17
rect 97 13 99 17
<< ndiffusion >>
rect 7 32 15 34
rect 7 28 8 32
rect 12 28 15 32
rect 7 14 15 28
rect 17 33 27 34
rect 17 17 29 33
rect 31 17 39 33
rect 41 17 49 33
rect 51 29 56 33
rect 51 22 61 29
rect 51 18 54 22
rect 58 18 61 22
rect 51 17 61 18
rect 63 25 70 29
rect 63 22 73 25
rect 63 18 66 22
rect 70 18 73 22
rect 63 17 73 18
rect 75 17 85 25
rect 87 22 97 25
rect 87 18 90 22
rect 94 18 97 22
rect 87 17 97 18
rect 99 22 107 25
rect 99 18 102 22
rect 106 18 107 22
rect 99 17 107 18
rect 17 14 27 17
rect 21 12 27 14
rect 21 8 22 12
rect 26 8 27 12
rect 77 12 83 17
rect 21 7 27 8
rect 77 8 78 12
rect 82 8 83 12
rect 77 7 83 8
<< pdiffusion >>
rect 7 82 15 94
rect 7 78 8 82
rect 12 78 15 82
rect 7 72 15 78
rect 7 68 8 72
rect 12 68 15 72
rect 7 62 15 68
rect 7 58 8 62
rect 12 58 15 62
rect 7 55 15 58
rect 17 85 24 94
rect 43 92 49 93
rect 43 88 44 92
rect 48 88 49 92
rect 43 85 49 88
rect 17 82 27 85
rect 17 78 20 82
rect 24 78 27 82
rect 17 63 27 78
rect 29 82 39 85
rect 29 78 32 82
rect 36 78 39 82
rect 29 63 39 78
rect 41 63 51 85
rect 53 82 63 85
rect 53 78 56 82
rect 60 78 63 82
rect 53 63 63 78
rect 17 55 24 63
rect 56 61 63 63
rect 65 72 77 85
rect 65 68 68 72
rect 72 68 77 72
rect 65 62 77 68
rect 65 61 68 62
rect 67 58 68 61
rect 72 58 77 62
rect 67 57 77 58
rect 72 56 77 57
rect 79 56 87 85
rect 89 56 97 85
rect 92 55 97 56
rect 99 82 107 85
rect 99 78 102 82
rect 106 78 107 82
rect 99 55 107 78
<< metal1 >>
rect -2 96 112 100
rect -2 92 56 96
rect 60 92 68 96
rect 72 92 80 96
rect 84 92 92 96
rect 96 92 112 96
rect -2 88 44 92
rect 48 88 112 92
rect 8 82 12 83
rect 8 72 12 78
rect 20 82 24 88
rect 31 78 32 82
rect 36 78 56 82
rect 60 78 102 82
rect 106 78 107 82
rect 20 77 24 78
rect 8 62 12 68
rect 8 32 12 58
rect 8 17 12 28
rect 18 42 22 43
rect 18 22 22 38
rect 28 42 32 73
rect 28 27 32 38
rect 38 42 42 73
rect 38 27 42 38
rect 48 42 52 73
rect 48 37 52 38
rect 58 42 62 73
rect 58 37 62 38
rect 68 72 72 73
rect 68 62 72 68
rect 68 32 72 58
rect 54 28 72 32
rect 78 52 82 73
rect 54 22 58 28
rect 78 27 82 48
rect 88 52 92 73
rect 88 27 92 48
rect 98 42 102 73
rect 98 27 102 38
rect 102 22 106 23
rect 18 18 54 22
rect 65 18 66 22
rect 70 18 90 22
rect 94 18 95 22
rect 54 17 58 18
rect 102 12 106 18
rect -2 8 22 12
rect 26 10 78 12
rect 26 8 34 10
rect -2 6 34 8
rect 38 6 44 10
rect 48 6 54 10
rect 58 6 65 10
rect 69 8 78 10
rect 82 10 112 12
rect 82 8 92 10
rect 69 6 92 8
rect 96 6 100 10
rect 104 6 112 10
rect -2 0 112 6
<< ntransistor >>
rect 15 14 17 34
rect 29 17 31 33
rect 39 17 41 33
rect 49 17 51 33
rect 61 17 63 29
rect 73 17 75 25
rect 85 17 87 25
rect 97 17 99 25
<< ptransistor >>
rect 15 55 17 94
rect 27 63 29 85
rect 39 63 41 85
rect 51 63 53 85
rect 63 61 65 85
rect 77 56 79 85
rect 87 56 89 85
rect 97 55 99 85
<< polycontact >>
rect 18 38 22 42
rect 28 38 32 42
rect 38 38 42 42
rect 48 38 52 42
rect 58 38 62 42
rect 78 48 82 52
rect 88 48 92 52
rect 98 38 102 42
<< ndcontact >>
rect 8 28 12 32
rect 54 18 58 22
rect 66 18 70 22
rect 90 18 94 22
rect 102 18 106 22
rect 22 8 26 12
rect 78 8 82 12
<< pdcontact >>
rect 8 78 12 82
rect 8 68 12 72
rect 8 58 12 62
rect 44 88 48 92
rect 20 78 24 82
rect 32 78 36 82
rect 56 78 60 82
rect 68 68 72 72
rect 68 58 72 62
rect 102 78 106 82
<< psubstratepcontact >>
rect 34 6 38 10
rect 44 6 48 10
rect 54 6 58 10
rect 65 6 69 10
rect 92 6 96 10
rect 100 6 104 10
<< nsubstratencontact >>
rect 56 92 60 96
rect 68 92 72 96
rect 80 92 84 96
rect 92 92 96 96
<< psubstratepdiff >>
rect 33 10 70 11
rect 33 6 34 10
rect 38 6 44 10
rect 48 6 54 10
rect 58 6 65 10
rect 69 6 70 10
rect 91 10 105 11
rect 33 5 70 6
rect 91 6 92 10
rect 96 6 100 10
rect 104 6 105 10
rect 91 5 105 6
<< nsubstratendiff >>
rect 55 96 97 97
rect 55 92 56 96
rect 60 92 68 96
rect 72 92 80 96
rect 84 92 92 96
rect 96 92 97 96
rect 55 91 97 92
<< labels >>
rlabel metal1 10 50 10 50 6 q
rlabel metal1 30 50 30 50 6 i0
rlabel metal1 40 50 40 50 6 i1
rlabel metal1 55 6 55 6 6 vss
rlabel metal1 60 55 60 55 6 i6
rlabel metal1 50 55 50 55 6 i2
rlabel metal1 55 94 55 94 6 vdd
rlabel polycontact 80 50 80 50 6 i3
rlabel polycontact 90 50 90 50 6 i4
rlabel metal1 100 50 100 50 6 i5
<< end >>
