magic
tech scmos
timestamp 1179385048
<< checkpaint >>
rect -22 -22 102 94
<< ab >>
rect 0 0 80 72
<< pwell >>
rect -4 -4 84 32
<< nwell >>
rect -4 32 84 76
<< polysilicon >>
rect 19 66 21 70
rect 29 66 31 70
rect 39 66 41 70
rect 49 66 51 70
rect 59 66 61 70
rect 9 57 11 61
rect 9 35 11 38
rect 19 35 21 38
rect 29 35 31 38
rect 39 35 41 38
rect 9 34 41 35
rect 9 33 32 34
rect 9 26 11 33
rect 19 26 21 33
rect 29 30 32 33
rect 36 33 41 34
rect 36 30 37 33
rect 49 32 51 39
rect 59 36 61 39
rect 58 35 64 36
rect 29 29 37 30
rect 48 31 54 32
rect 29 26 31 29
rect 48 28 49 31
rect 41 27 49 28
rect 53 27 54 31
rect 41 26 54 27
rect 58 31 59 35
rect 63 31 64 35
rect 58 30 64 31
rect 9 11 11 15
rect 41 17 43 26
rect 58 22 60 30
rect 48 20 60 22
rect 48 17 50 20
rect 58 17 60 20
rect 65 25 71 26
rect 65 21 66 25
rect 70 21 71 25
rect 65 20 71 21
rect 65 17 67 20
rect 19 2 21 6
rect 29 2 31 6
rect 41 2 43 6
rect 48 2 50 6
rect 58 2 60 6
rect 65 2 67 6
<< ndiffusion >>
rect 2 25 9 26
rect 2 21 3 25
rect 7 21 9 25
rect 2 20 9 21
rect 4 15 9 20
rect 11 20 19 26
rect 11 16 13 20
rect 17 16 19 20
rect 11 15 19 16
rect 13 6 19 15
rect 21 25 29 26
rect 21 21 23 25
rect 27 21 29 25
rect 21 18 29 21
rect 21 14 23 18
rect 27 14 29 18
rect 21 6 29 14
rect 31 19 39 26
rect 31 15 33 19
rect 37 17 39 19
rect 37 15 41 17
rect 31 11 41 15
rect 31 7 33 11
rect 37 7 41 11
rect 31 6 41 7
rect 43 6 48 17
rect 50 16 58 17
rect 50 12 52 16
rect 56 12 58 16
rect 50 6 58 12
rect 60 6 65 17
rect 67 11 74 17
rect 67 7 69 11
rect 73 7 74 11
rect 67 6 74 7
<< pdiffusion >>
rect 14 57 19 66
rect 2 56 9 57
rect 2 52 3 56
rect 7 52 9 56
rect 2 49 9 52
rect 2 45 3 49
rect 7 45 9 49
rect 2 38 9 45
rect 11 56 19 57
rect 11 52 13 56
rect 17 52 19 56
rect 11 49 19 52
rect 11 45 13 49
rect 17 45 19 49
rect 11 38 19 45
rect 21 65 29 66
rect 21 61 23 65
rect 27 61 29 65
rect 21 58 29 61
rect 21 54 23 58
rect 27 54 29 58
rect 21 38 29 54
rect 31 58 39 66
rect 31 54 33 58
rect 37 54 39 58
rect 31 51 39 54
rect 31 47 33 51
rect 37 47 39 51
rect 31 38 39 47
rect 41 65 49 66
rect 41 61 43 65
rect 47 61 49 65
rect 41 58 49 61
rect 41 54 43 58
rect 47 54 49 58
rect 41 39 49 54
rect 51 58 59 66
rect 51 54 53 58
rect 57 54 59 58
rect 51 51 59 54
rect 51 47 53 51
rect 57 47 59 51
rect 51 39 59 47
rect 61 59 67 66
rect 61 58 69 59
rect 61 54 63 58
rect 67 54 69 58
rect 61 51 69 54
rect 61 47 63 51
rect 67 47 69 51
rect 61 39 69 47
rect 41 38 47 39
<< metal1 >>
rect -2 68 82 72
rect -2 64 4 68
rect 8 65 72 68
rect 8 64 23 65
rect 3 56 7 64
rect 22 61 23 64
rect 27 64 43 65
rect 27 61 28 64
rect 22 58 28 61
rect 42 61 43 64
rect 47 64 72 65
rect 76 64 82 68
rect 47 61 48 64
rect 3 49 7 52
rect 12 52 13 56
rect 17 52 18 56
rect 22 54 23 58
rect 27 54 28 58
rect 33 58 38 59
rect 37 54 38 58
rect 42 58 48 61
rect 42 54 43 58
rect 47 54 48 58
rect 53 58 57 59
rect 12 50 18 52
rect 33 51 38 54
rect 12 49 33 50
rect 12 45 13 49
rect 17 47 33 49
rect 37 47 38 51
rect 53 51 57 54
rect 17 46 38 47
rect 41 47 53 50
rect 41 46 57 47
rect 63 58 67 64
rect 63 51 67 54
rect 63 46 67 47
rect 17 45 22 46
rect 3 44 7 45
rect 18 35 22 45
rect 2 30 27 35
rect 41 34 45 46
rect 58 35 63 43
rect 31 30 32 34
rect 36 30 45 34
rect 2 25 7 30
rect 2 21 3 25
rect 23 25 27 30
rect 2 20 7 21
rect 13 20 17 21
rect 13 8 17 16
rect 23 18 27 21
rect 23 13 27 14
rect 33 19 37 20
rect 33 11 37 15
rect 41 17 45 30
rect 49 31 54 35
rect 53 27 54 31
rect 58 31 59 35
rect 63 31 71 34
rect 58 30 71 31
rect 49 26 54 27
rect 49 25 71 26
rect 49 21 66 25
rect 70 21 71 25
rect 41 16 57 17
rect 41 13 52 16
rect 51 12 52 13
rect 56 12 57 16
rect -2 4 4 8
rect 8 7 33 8
rect 69 11 73 12
rect 37 7 69 8
rect 73 7 82 8
rect 8 4 82 7
rect -2 0 82 4
<< ntransistor >>
rect 9 15 11 26
rect 19 6 21 26
rect 29 6 31 26
rect 41 6 43 17
rect 48 6 50 17
rect 58 6 60 17
rect 65 6 67 17
<< ptransistor >>
rect 9 38 11 57
rect 19 38 21 66
rect 29 38 31 66
rect 39 38 41 66
rect 49 39 51 66
rect 59 39 61 66
<< polycontact >>
rect 32 30 36 34
rect 49 27 53 31
rect 59 31 63 35
rect 66 21 70 25
<< ndcontact >>
rect 3 21 7 25
rect 13 16 17 20
rect 23 21 27 25
rect 23 14 27 18
rect 33 15 37 19
rect 33 7 37 11
rect 52 12 56 16
rect 69 7 73 11
<< pdcontact >>
rect 3 52 7 56
rect 3 45 7 49
rect 13 52 17 56
rect 13 45 17 49
rect 23 61 27 65
rect 23 54 27 58
rect 33 54 37 58
rect 33 47 37 51
rect 43 61 47 65
rect 43 54 47 58
rect 53 54 57 58
rect 53 47 57 51
rect 63 54 67 58
rect 63 47 67 51
<< psubstratepcontact >>
rect 4 4 8 8
<< nsubstratencontact >>
rect 4 64 8 68
rect 72 64 76 68
<< psubstratepdiff >>
rect 3 8 9 9
rect 3 4 4 8
rect 8 4 9 8
rect 3 3 9 4
<< nsubstratendiff >>
rect 3 68 9 69
rect 3 64 4 68
rect 8 64 9 68
rect 71 68 77 69
rect 3 63 9 64
rect 71 64 72 68
rect 76 64 77 68
rect 71 63 77 64
<< labels >>
rlabel metal1 4 28 4 28 6 z
rlabel metal1 12 32 12 32 6 z
rlabel metal1 20 40 20 40 6 z
rlabel metal1 28 48 28 48 6 z
rlabel metal1 40 4 40 4 6 vss
rlabel metal1 38 32 38 32 6 zn
rlabel pdcontact 36 56 36 56 6 z
rlabel metal1 40 68 40 68 6 vdd
rlabel ndcontact 54 14 54 14 6 zn
rlabel metal1 60 24 60 24 6 a
rlabel polycontact 52 28 52 28 6 a
rlabel metal1 60 40 60 40 6 b
rlabel metal1 55 52 55 52 6 zn
rlabel polycontact 68 24 68 24 6 a
rlabel metal1 68 32 68 32 6 b
<< end >>
