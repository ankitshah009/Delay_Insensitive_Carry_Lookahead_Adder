magic
tech scmos
timestamp 1179385577
<< checkpaint >>
rect -22 -22 54 94
<< ab >>
rect 0 0 32 72
<< pwell >>
rect -4 -4 36 32
<< nwell >>
rect -4 32 36 76
<< polysilicon >>
rect 9 56 11 61
rect 21 56 23 61
rect 9 35 11 38
rect 21 35 23 38
rect 9 34 15 35
rect 9 30 10 34
rect 14 30 15 34
rect 9 29 15 30
rect 21 34 27 35
rect 21 30 22 34
rect 26 30 27 34
rect 21 29 27 30
rect 9 22 11 29
rect 21 26 23 29
rect 9 8 11 13
rect 21 12 23 17
<< ndiffusion >>
rect 13 22 21 26
rect 4 19 9 22
rect 2 18 9 19
rect 2 14 3 18
rect 7 14 9 18
rect 2 13 9 14
rect 11 18 21 22
rect 11 14 14 18
rect 18 17 21 18
rect 23 25 30 26
rect 23 21 25 25
rect 29 21 30 25
rect 23 20 30 21
rect 23 17 28 20
rect 18 14 19 17
rect 11 13 19 14
<< pdiffusion >>
rect 13 68 19 69
rect 13 64 14 68
rect 18 64 19 68
rect 13 56 19 64
rect 2 55 9 56
rect 2 51 3 55
rect 7 51 9 55
rect 2 48 9 51
rect 2 44 3 48
rect 7 44 9 48
rect 2 43 9 44
rect 4 38 9 43
rect 11 38 21 56
rect 23 51 28 56
rect 23 50 30 51
rect 23 46 25 50
rect 29 46 30 50
rect 23 45 30 46
rect 23 38 28 45
<< metal1 >>
rect -2 68 34 72
rect -2 64 4 68
rect 8 64 14 68
rect 18 64 24 68
rect 28 64 34 68
rect 2 55 14 59
rect 2 51 3 55
rect 7 53 14 55
rect 2 48 7 51
rect 2 44 3 48
rect 2 43 7 44
rect 10 46 25 50
rect 29 46 30 50
rect 2 19 6 43
rect 10 34 14 46
rect 26 35 30 43
rect 10 25 14 30
rect 18 34 30 35
rect 18 30 22 34
rect 26 30 30 34
rect 18 29 30 30
rect 10 21 25 25
rect 29 21 30 25
rect 2 18 7 19
rect 2 14 3 18
rect 2 13 7 14
rect 13 14 14 18
rect 18 14 19 18
rect 13 8 19 14
rect -2 4 21 8
rect 25 4 34 8
rect -2 0 34 4
<< ntransistor >>
rect 9 13 11 22
rect 21 17 23 26
<< ptransistor >>
rect 9 38 11 56
rect 21 38 23 56
<< polycontact >>
rect 10 30 14 34
rect 22 30 26 34
<< ndcontact >>
rect 3 14 7 18
rect 14 14 18 18
rect 25 21 29 25
<< pdcontact >>
rect 14 64 18 68
rect 3 51 7 55
rect 3 44 7 48
rect 25 46 29 50
<< psubstratepcontact >>
rect 21 4 25 8
<< nsubstratencontact >>
rect 4 64 8 68
rect 24 64 28 68
<< psubstratepdiff >>
rect 17 8 29 9
rect 17 4 21 8
rect 25 4 29 8
rect 17 3 29 4
<< nsubstratendiff >>
rect 3 68 9 69
rect 3 64 4 68
rect 8 64 9 68
rect 3 63 9 64
rect 23 68 29 69
rect 23 64 24 68
rect 28 64 29 68
rect 23 63 29 64
<< labels >>
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 35 12 35 6 an
rlabel metal1 12 56 12 56 6 z
rlabel metal1 16 4 16 4 6 vss
rlabel metal1 20 32 20 32 6 a
rlabel metal1 16 68 16 68 6 vdd
rlabel metal1 20 23 20 23 6 an
rlabel metal1 28 36 28 36 6 a
rlabel metal1 20 48 20 48 6 an
<< end >>
