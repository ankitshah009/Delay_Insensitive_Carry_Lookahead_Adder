magic
tech scmos
timestamp 1179385590
<< checkpaint >>
rect -22 -25 54 105
<< ab >>
rect 0 0 32 80
<< pwell >>
rect -4 -7 36 36
<< nwell >>
rect -4 36 36 87
<< polysilicon >>
rect 9 70 11 74
rect 19 70 21 74
rect 9 39 11 42
rect 19 39 21 42
rect 9 38 15 39
rect 9 34 10 38
rect 14 34 15 38
rect 9 33 15 34
rect 19 38 25 39
rect 19 34 20 38
rect 24 34 25 38
rect 19 33 25 34
rect 9 30 11 33
rect 19 30 21 33
rect 9 11 11 16
rect 19 11 21 16
<< ndiffusion >>
rect 2 29 9 30
rect 2 25 3 29
rect 7 25 9 29
rect 2 22 9 25
rect 2 18 3 22
rect 7 18 9 22
rect 2 16 9 18
rect 11 21 19 30
rect 11 17 13 21
rect 17 17 19 21
rect 11 16 19 17
rect 21 29 28 30
rect 21 25 23 29
rect 27 25 28 29
rect 21 22 28 25
rect 21 18 23 22
rect 27 18 28 22
rect 21 16 28 18
<< pdiffusion >>
rect 4 55 9 70
rect 2 54 9 55
rect 2 50 3 54
rect 7 50 9 54
rect 2 47 9 50
rect 2 43 3 47
rect 7 43 9 47
rect 2 42 9 43
rect 11 69 19 70
rect 11 65 13 69
rect 17 65 19 69
rect 11 42 19 65
rect 21 55 26 70
rect 21 54 28 55
rect 21 50 23 54
rect 27 50 28 54
rect 21 49 28 50
rect 21 42 26 49
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect -2 69 34 78
rect -2 68 13 69
rect 12 65 13 68
rect 17 68 34 69
rect 17 65 18 68
rect 2 62 7 63
rect 2 58 15 62
rect 2 54 7 58
rect 2 50 3 54
rect 2 47 7 50
rect 2 43 3 47
rect 2 42 7 43
rect 10 50 23 54
rect 27 50 28 54
rect 2 30 6 42
rect 10 38 14 50
rect 26 39 30 47
rect 2 29 7 30
rect 2 25 3 29
rect 10 29 14 34
rect 18 38 30 39
rect 18 34 20 38
rect 24 34 30 38
rect 18 33 30 34
rect 10 25 23 29
rect 27 25 28 29
rect 2 22 7 25
rect 2 18 3 22
rect 23 22 28 25
rect 2 17 7 18
rect 12 17 13 21
rect 17 17 18 21
rect 27 18 28 22
rect 23 17 28 18
rect 12 12 18 17
rect -2 2 34 12
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
<< ntransistor >>
rect 9 16 11 30
rect 19 16 21 30
<< ptransistor >>
rect 9 42 11 70
rect 19 42 21 70
<< polycontact >>
rect 10 34 14 38
rect 20 34 24 38
<< ndcontact >>
rect 3 25 7 29
rect 3 18 7 22
rect 13 17 17 21
rect 23 25 27 29
rect 23 18 27 22
<< pdcontact >>
rect 3 50 7 54
rect 3 43 7 47
rect 13 65 17 69
rect 23 50 27 54
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
<< psubstratepdiff >>
rect 0 2 32 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 32 2
rect 0 -3 32 -2
<< nsubstratendiff >>
rect 0 82 32 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 32 82
rect 0 77 32 78
<< labels >>
rlabel polycontact 12 36 12 36 6 an
rlabel metal1 4 40 4 40 6 z
rlabel metal1 12 39 12 39 6 an
rlabel metal1 12 60 12 60 6 z
rlabel metal1 16 6 16 6 6 vss
rlabel metal1 20 36 20 36 6 a
rlabel metal1 16 74 16 74 6 vdd
rlabel metal1 25 23 25 23 6 an
rlabel metal1 28 40 28 40 6 a
rlabel metal1 19 52 19 52 6 an
<< end >>
