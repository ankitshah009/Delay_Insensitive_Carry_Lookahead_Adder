magic
tech scmos
timestamp 1182081803
<< checkpaint >>
rect -25 -26 57 114
<< ab >>
rect 0 0 32 88
<< pwell >>
rect -7 -8 39 40
<< nwell >>
rect -7 40 39 96
<< polysilicon >>
rect 5 80 14 86
rect 18 80 27 86
rect 9 77 11 80
rect 21 77 23 80
rect 9 48 11 51
rect 21 48 23 51
rect 2 47 11 48
rect 2 43 6 47
rect 10 43 11 47
rect 2 42 11 43
rect 15 47 30 48
rect 15 43 22 47
rect 26 43 30 47
rect 15 42 30 43
rect 2 37 17 38
rect 2 33 6 37
rect 10 33 17 37
rect 2 32 17 33
rect 21 37 30 38
rect 21 33 22 37
rect 26 33 30 37
rect 21 32 30 33
rect 9 29 11 32
rect 21 29 23 32
rect 9 8 11 11
rect 21 8 23 11
rect 5 2 14 8
rect 18 2 27 8
<< ndiffusion >>
rect 2 16 9 29
rect 2 12 3 16
rect 7 12 9 16
rect 2 11 9 12
rect 11 26 21 29
rect 11 22 14 26
rect 18 22 21 26
rect 11 18 21 22
rect 11 14 14 18
rect 18 14 21 18
rect 11 11 21 14
rect 23 24 30 29
rect 23 20 25 24
rect 29 20 30 24
rect 23 17 30 20
rect 23 13 25 17
rect 29 13 30 17
rect 23 11 30 13
<< pdiffusion >>
rect 2 75 9 77
rect 2 71 3 75
rect 7 71 9 75
rect 2 68 9 71
rect 2 64 3 68
rect 7 64 9 68
rect 2 51 9 64
rect 11 51 21 77
rect 23 67 30 77
rect 23 63 25 67
rect 29 63 30 67
rect 23 60 30 63
rect 23 56 25 60
rect 29 56 30 60
rect 23 51 30 56
<< metal1 >>
rect -2 86 2 90
rect 30 86 34 90
rect 2 82 7 85
rect -2 81 7 82
rect 30 81 34 82
rect 3 75 7 81
rect 3 68 7 71
rect 3 63 7 64
rect 22 67 29 68
rect 22 63 25 67
rect 22 60 29 63
rect 22 59 25 60
rect 14 56 25 59
rect 14 55 29 56
rect 6 47 10 48
rect 6 37 10 43
rect 6 21 10 33
rect 14 26 18 55
rect 22 47 26 51
rect 22 37 26 43
rect 22 29 26 33
rect 14 18 18 22
rect 3 16 7 17
rect 14 13 18 14
rect 25 24 29 25
rect 25 17 29 20
rect 3 7 7 12
rect -2 6 7 7
rect 2 3 7 6
rect 25 7 29 13
rect 25 6 34 7
rect 25 3 30 6
rect -2 -2 2 2
rect 30 -2 34 2
<< metal2 >>
rect -2 86 34 90
rect 2 82 30 86
rect -2 80 34 82
rect -2 6 34 8
rect 2 2 30 6
rect -2 -2 34 2
<< ntransistor >>
rect 9 11 11 29
rect 21 11 23 29
<< ptransistor >>
rect 9 51 11 77
rect 21 51 23 77
<< polycontact >>
rect 6 43 10 47
rect 22 43 26 47
rect 6 33 10 37
rect 22 33 26 37
<< ndcontact >>
rect 3 12 7 16
rect 14 22 18 26
rect 14 14 18 18
rect 25 20 29 24
rect 25 13 29 17
<< pdcontact >>
rect 3 71 7 75
rect 3 64 7 68
rect 25 63 29 67
rect 25 56 29 60
<< m2contact >>
rect -2 82 2 86
rect 30 82 34 86
rect -2 2 2 6
rect 30 2 34 6
<< psubstratepcontact >>
rect -2 2 2 6
rect 30 2 34 6
<< nsubstratencontact >>
rect -2 82 2 86
rect 30 82 34 86
<< psubstratepdiff >>
rect -3 6 3 7
rect -3 2 -2 6
rect 2 2 3 6
rect 29 6 35 7
rect 29 2 30 6
rect 34 2 35 6
rect -3 0 3 2
rect 29 0 35 2
<< nsubstratendiff >>
rect -3 86 3 88
rect 29 86 35 88
rect -3 82 -2 86
rect 2 82 3 86
rect -3 81 3 82
rect 29 82 30 86
rect 34 82 35 86
rect 29 81 35 82
<< labels >>
rlabel metal1 8 32 8 32 6 a
rlabel metal1 16 36 16 36 6 z
rlabel metal1 24 40 24 40 6 b
rlabel metal1 24 64 24 64 6 z
rlabel metal2 16 4 16 4 6 vss
rlabel metal2 16 84 16 84 6 vdd
<< end >>
