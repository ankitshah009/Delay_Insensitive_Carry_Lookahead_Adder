magic
tech scmos
timestamp 1185039163
<< checkpaint >>
rect -22 -24 152 124
<< ab >>
rect 0 0 130 100
<< pwell >>
rect -2 -4 132 49
<< nwell >>
rect -2 49 132 104
<< polysilicon >>
rect 17 95 19 98
rect 29 95 31 98
rect 41 95 43 98
rect 53 95 55 98
rect 65 95 67 98
rect 93 85 95 88
rect 105 85 107 88
rect 117 85 119 88
rect 65 63 67 75
rect 75 66 81 67
rect 65 62 71 63
rect 65 58 66 62
rect 70 58 71 62
rect 75 62 76 66
rect 80 63 81 66
rect 93 63 95 65
rect 80 62 95 63
rect 75 61 95 62
rect 65 57 71 58
rect 105 57 107 65
rect 117 63 119 65
rect 111 62 119 63
rect 111 58 112 62
rect 116 58 119 62
rect 111 57 119 58
rect 65 56 107 57
rect 65 55 96 56
rect 17 47 19 55
rect 29 47 31 55
rect 41 47 43 55
rect 53 47 55 55
rect 95 52 96 55
rect 100 55 107 56
rect 100 52 101 55
rect 95 51 101 52
rect 121 48 127 49
rect 121 47 122 48
rect 17 45 122 47
rect 121 44 122 45
rect 126 44 127 48
rect 121 43 127 44
rect 17 38 91 39
rect 17 37 86 38
rect 17 25 19 37
rect 29 25 31 37
rect 41 25 43 37
rect 53 25 55 37
rect 85 34 86 37
rect 90 34 91 38
rect 85 33 91 34
rect 95 38 119 39
rect 95 34 96 38
rect 100 37 119 38
rect 100 34 101 37
rect 95 33 101 34
rect 59 32 67 33
rect 59 28 60 32
rect 64 28 67 32
rect 59 27 67 28
rect 75 32 81 33
rect 75 28 76 32
rect 80 29 81 32
rect 105 32 113 33
rect 80 28 95 29
rect 75 27 95 28
rect 65 25 67 27
rect 93 25 95 27
rect 105 28 108 32
rect 112 28 113 32
rect 105 27 113 28
rect 105 25 107 27
rect 117 25 119 37
rect 65 12 67 15
rect 93 12 95 15
rect 105 12 107 15
rect 117 12 119 15
rect 17 2 19 5
rect 29 2 31 5
rect 41 2 43 5
rect 53 2 55 5
<< ndiffusion >>
rect 9 22 17 25
rect 9 18 10 22
rect 14 18 17 22
rect 9 12 17 18
rect 9 8 10 12
rect 14 8 17 12
rect 9 5 17 8
rect 19 22 29 25
rect 19 18 22 22
rect 26 18 29 22
rect 19 5 29 18
rect 31 22 41 25
rect 31 18 34 22
rect 38 18 41 22
rect 31 12 41 18
rect 31 8 34 12
rect 38 8 41 12
rect 31 5 41 8
rect 43 22 53 25
rect 43 18 46 22
rect 50 18 53 22
rect 43 5 53 18
rect 55 15 65 25
rect 67 22 75 25
rect 67 18 70 22
rect 74 18 75 22
rect 67 15 75 18
rect 85 22 93 25
rect 85 18 86 22
rect 90 18 93 22
rect 85 15 93 18
rect 95 15 105 25
rect 107 22 117 25
rect 107 18 110 22
rect 114 18 117 22
rect 107 15 117 18
rect 119 22 127 25
rect 119 18 122 22
rect 126 18 127 22
rect 119 15 127 18
rect 55 12 63 15
rect 97 12 103 15
rect 55 8 58 12
rect 62 8 63 12
rect 55 5 63 8
rect 97 8 98 12
rect 102 8 103 12
rect 97 7 103 8
<< pdiffusion >>
rect 9 92 17 95
rect 9 88 10 92
rect 14 88 17 92
rect 9 82 17 88
rect 9 78 10 82
rect 14 78 17 82
rect 9 72 17 78
rect 9 68 10 72
rect 14 68 17 72
rect 9 62 17 68
rect 9 58 10 62
rect 14 58 17 62
rect 9 55 17 58
rect 19 82 29 95
rect 19 78 22 82
rect 26 78 29 82
rect 19 72 29 78
rect 19 68 22 72
rect 26 68 29 72
rect 19 62 29 68
rect 19 58 22 62
rect 26 58 29 62
rect 19 55 29 58
rect 31 92 41 95
rect 31 88 34 92
rect 38 88 41 92
rect 31 82 41 88
rect 31 78 34 82
rect 38 78 41 82
rect 31 72 41 78
rect 31 68 34 72
rect 38 68 41 72
rect 31 62 41 68
rect 31 58 34 62
rect 38 58 41 62
rect 31 55 41 58
rect 43 82 53 95
rect 43 78 46 82
rect 50 78 53 82
rect 43 72 53 78
rect 43 68 46 72
rect 50 68 53 72
rect 43 62 53 68
rect 43 58 46 62
rect 50 58 53 62
rect 43 55 53 58
rect 55 92 65 95
rect 55 88 58 92
rect 62 88 65 92
rect 55 75 65 88
rect 67 82 75 95
rect 109 92 115 93
rect 109 88 110 92
rect 114 88 115 92
rect 109 85 115 88
rect 67 78 70 82
rect 74 78 75 82
rect 67 75 75 78
rect 85 82 93 85
rect 85 78 86 82
rect 90 78 93 82
rect 55 55 63 75
rect 85 72 93 78
rect 85 68 86 72
rect 90 68 93 72
rect 85 65 93 68
rect 95 82 105 85
rect 95 78 98 82
rect 102 78 105 82
rect 95 72 105 78
rect 95 68 98 72
rect 102 68 105 72
rect 95 65 105 68
rect 107 65 117 85
rect 119 82 127 85
rect 119 78 122 82
rect 126 78 127 82
rect 119 72 127 78
rect 119 68 122 72
rect 126 68 127 72
rect 119 65 127 68
<< metal1 >>
rect -2 96 132 101
rect -2 92 82 96
rect 86 92 98 96
rect 102 92 132 96
rect -2 88 10 92
rect 14 88 34 92
rect 38 88 58 92
rect 62 88 110 92
rect 114 88 132 92
rect -2 87 132 88
rect 9 82 15 87
rect 9 78 10 82
rect 14 78 15 82
rect 9 72 15 78
rect 9 68 10 72
rect 14 68 15 72
rect 9 62 15 68
rect 9 58 10 62
rect 14 58 15 62
rect 9 57 15 58
rect 21 82 27 83
rect 21 78 22 82
rect 26 78 27 82
rect 21 72 27 78
rect 21 68 22 72
rect 26 68 27 72
rect 21 62 27 68
rect 21 58 22 62
rect 26 58 27 62
rect 21 45 27 58
rect 33 82 39 87
rect 33 78 34 82
rect 38 78 39 82
rect 33 72 39 78
rect 45 82 53 83
rect 69 82 80 83
rect 45 78 46 82
rect 50 78 53 82
rect 45 77 53 78
rect 47 73 53 77
rect 33 68 34 72
rect 38 68 39 72
rect 33 62 39 68
rect 45 72 53 73
rect 45 68 46 72
rect 50 68 53 72
rect 45 67 53 68
rect 47 63 53 67
rect 33 58 34 62
rect 38 58 39 62
rect 33 57 39 58
rect 45 62 53 63
rect 45 58 46 62
rect 50 58 53 62
rect 45 57 53 58
rect 47 45 53 57
rect 21 39 53 45
rect 9 22 15 23
rect 9 18 10 22
rect 14 18 15 22
rect 9 13 15 18
rect 21 22 27 39
rect 47 23 53 39
rect 21 18 22 22
rect 26 18 27 22
rect 21 17 27 18
rect 33 22 39 23
rect 33 18 34 22
rect 38 18 39 22
rect 33 13 39 18
rect 45 22 53 23
rect 45 18 46 22
rect 50 18 53 22
rect 57 63 63 82
rect 69 78 70 82
rect 74 78 80 82
rect 69 77 80 78
rect 85 82 91 83
rect 85 78 86 82
rect 90 78 91 82
rect 85 77 91 78
rect 97 82 103 83
rect 121 82 127 83
rect 97 78 98 82
rect 102 78 122 82
rect 126 78 127 82
rect 97 77 103 78
rect 121 77 127 78
rect 76 67 80 77
rect 86 73 90 77
rect 98 73 102 77
rect 122 73 126 77
rect 85 72 91 73
rect 85 68 86 72
rect 90 68 91 72
rect 85 67 91 68
rect 97 72 103 73
rect 121 72 127 73
rect 97 68 98 72
rect 102 68 103 72
rect 97 67 103 68
rect 75 66 81 67
rect 57 62 71 63
rect 57 58 66 62
rect 70 58 71 62
rect 75 62 76 66
rect 80 62 81 66
rect 75 61 81 62
rect 57 57 71 58
rect 57 33 63 57
rect 76 33 80 61
rect 86 39 90 67
rect 107 63 113 72
rect 121 68 122 72
rect 126 68 127 72
rect 121 67 127 68
rect 107 62 117 63
rect 107 58 112 62
rect 116 58 117 62
rect 107 57 117 58
rect 95 56 101 57
rect 95 52 96 56
rect 100 52 101 56
rect 95 51 101 52
rect 96 39 100 51
rect 85 38 91 39
rect 85 34 86 38
rect 90 34 91 38
rect 85 33 91 34
rect 95 38 101 39
rect 95 34 96 38
rect 100 34 101 38
rect 95 33 101 34
rect 57 32 65 33
rect 57 28 60 32
rect 64 28 65 32
rect 57 27 65 28
rect 75 32 81 33
rect 75 28 76 32
rect 80 28 81 32
rect 75 27 81 28
rect 57 18 63 27
rect 76 23 80 27
rect 86 23 90 33
rect 107 32 113 57
rect 122 49 126 67
rect 121 48 127 49
rect 121 44 122 48
rect 126 44 127 48
rect 121 43 127 44
rect 107 28 108 32
rect 112 28 113 32
rect 107 27 113 28
rect 122 23 126 43
rect 69 22 80 23
rect 69 18 70 22
rect 74 18 80 22
rect 45 17 53 18
rect 69 17 80 18
rect 85 22 91 23
rect 109 22 115 23
rect 85 18 86 22
rect 90 18 110 22
rect 114 18 115 22
rect 85 17 91 18
rect 109 17 115 18
rect 121 22 127 23
rect 121 18 122 22
rect 126 18 127 22
rect 121 17 127 18
rect -2 12 132 13
rect -2 8 10 12
rect 14 8 34 12
rect 38 8 58 12
rect 62 8 98 12
rect 102 8 132 12
rect -2 4 70 8
rect 74 4 86 8
rect 90 4 110 8
rect 114 4 122 8
rect 126 4 132 8
rect -2 -1 132 4
<< ntransistor >>
rect 17 5 19 25
rect 29 5 31 25
rect 41 5 43 25
rect 53 5 55 25
rect 65 15 67 25
rect 93 15 95 25
rect 105 15 107 25
rect 117 15 119 25
<< ptransistor >>
rect 17 55 19 95
rect 29 55 31 95
rect 41 55 43 95
rect 53 55 55 95
rect 65 75 67 95
rect 93 65 95 85
rect 105 65 107 85
rect 117 65 119 85
<< polycontact >>
rect 66 58 70 62
rect 76 62 80 66
rect 112 58 116 62
rect 96 52 100 56
rect 122 44 126 48
rect 86 34 90 38
rect 96 34 100 38
rect 60 28 64 32
rect 76 28 80 32
rect 108 28 112 32
<< ndcontact >>
rect 10 18 14 22
rect 10 8 14 12
rect 22 18 26 22
rect 34 18 38 22
rect 34 8 38 12
rect 46 18 50 22
rect 70 18 74 22
rect 86 18 90 22
rect 110 18 114 22
rect 122 18 126 22
rect 58 8 62 12
rect 98 8 102 12
<< pdcontact >>
rect 10 88 14 92
rect 10 78 14 82
rect 10 68 14 72
rect 10 58 14 62
rect 22 78 26 82
rect 22 68 26 72
rect 22 58 26 62
rect 34 88 38 92
rect 34 78 38 82
rect 34 68 38 72
rect 34 58 38 62
rect 46 78 50 82
rect 46 68 50 72
rect 46 58 50 62
rect 58 88 62 92
rect 110 88 114 92
rect 70 78 74 82
rect 86 78 90 82
rect 86 68 90 72
rect 98 78 102 82
rect 98 68 102 72
rect 122 78 126 82
rect 122 68 126 72
<< psubstratepcontact >>
rect 70 4 74 8
rect 86 4 90 8
rect 110 4 114 8
rect 122 4 126 8
<< nsubstratencontact >>
rect 82 92 86 96
rect 98 92 102 96
<< psubstratepdiff >>
rect 69 8 91 9
rect 69 4 70 8
rect 74 4 86 8
rect 90 4 91 8
rect 109 8 127 9
rect 69 3 91 4
rect 109 4 110 8
rect 114 4 122 8
rect 126 4 127 8
rect 109 3 127 4
<< nsubstratendiff >>
rect 81 96 103 97
rect 81 92 82 96
rect 86 92 98 96
rect 102 92 103 96
rect 81 91 103 92
<< labels >>
rlabel metal1 50 50 50 50 6 q
rlabel metal1 60 50 60 50 6 cmd
rlabel metal1 60 50 60 50 6 cmd
rlabel metal1 50 50 50 50 6 q
rlabel metal1 65 6 65 6 6 vss
rlabel metal1 65 6 65 6 6 vss
rlabel metal1 65 94 65 94 6 vdd
rlabel metal1 65 94 65 94 6 vdd
rlabel metal1 110 50 110 50 6 i
rlabel metal1 110 50 110 50 6 i
<< end >>
