.subckt iv1v1x4 a vdd vss z
*   SPICE3 file   created from iv1v1x4.ext -      technology: scmos
m00 z      a      vdd    vdd p w=28u  l=2.3636u ad=112p     pd=36u      as=210p     ps=71u
m01 vdd    a      z      vdd p w=28u  l=2.3636u ad=210p     pd=71u      as=112p     ps=36u
m02 z      a      vss    vss n w=19u  l=2.3636u ad=76p      pd=27u      as=142.5p   ps=53u
m03 vss    a      z      vss n w=19u  l=2.3636u ad=142.5p   pd=53u      as=76p      ps=27u
C0  vss    a      0.036f
C1  z      vdd    0.187f
C2  vss    z      0.220f
C3  z      a      0.109f
C4  vss    vdd    0.010f
C5  a      vdd    0.037f
C7  z      vss    0.006f
C8  a      vss    0.035f
.ends
