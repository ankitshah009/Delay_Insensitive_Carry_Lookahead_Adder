.subckt bf1_y05 a vdd vss z
*   SPICE3 file   created from bf1_y05.ext -      technology: scmos
m00 vdd    an     z      vdd p w=12u  l=2.3636u ad=72p      pd=26u      as=78p      ps=40u
m01 an     a      vdd    vdd p w=12u  l=2.3636u ad=78p      pd=40u      as=72p      ps=26u
m02 vss    an     z      vss n w=6u   l=2.3636u ad=60p      pd=26u      as=48p      ps=28u
m03 an     a      vss    vss n w=6u   l=2.3636u ad=48p      pd=28u      as=60p      ps=26u
C0  vss    z      0.011f
C1  a      an     0.278f
C2  z      vdd    0.011f
C3  vss    a      0.005f
C4  vss    an     0.075f
C5  a      z      0.049f
C6  a      vdd    0.005f
C7  z      an     0.222f
C8  an     vdd    0.075f
C10 a      vss    0.031f
C11 z      vss    0.017f
C12 an     vss    0.040f
.ends
