magic
tech scmos
timestamp 1179387037
<< checkpaint >>
rect -22 -25 110 105
<< ab >>
rect 0 0 88 80
<< pwell >>
rect -4 -7 92 36
<< nwell >>
rect -4 36 92 87
<< polysilicon >>
rect 32 67 34 72
rect 39 67 41 72
rect 49 67 51 72
rect 56 67 58 72
rect 66 67 68 72
rect 73 67 75 72
rect 9 61 11 65
rect 22 63 24 67
rect 9 39 11 42
rect 22 39 24 42
rect 32 39 34 42
rect 39 39 41 42
rect 49 39 51 42
rect 56 39 58 42
rect 66 39 68 42
rect 9 38 24 39
rect 9 34 10 38
rect 14 34 24 38
rect 9 33 24 34
rect 29 38 35 39
rect 29 34 30 38
rect 34 34 35 38
rect 29 33 35 34
rect 39 38 52 39
rect 39 34 47 38
rect 51 34 52 38
rect 56 38 68 39
rect 56 37 60 38
rect 39 33 52 34
rect 59 34 60 37
rect 64 37 68 38
rect 73 39 75 42
rect 73 38 79 39
rect 64 34 65 37
rect 59 33 65 34
rect 73 34 74 38
rect 78 34 79 38
rect 73 33 79 34
rect 10 30 12 33
rect 20 30 22 33
rect 30 30 32 33
rect 40 30 42 33
rect 50 30 52 33
rect 62 30 64 33
rect 10 8 12 13
rect 20 8 22 13
rect 30 8 32 13
rect 40 8 42 13
rect 50 8 52 13
rect 62 8 64 13
<< ndiffusion >>
rect 5 22 10 30
rect 3 21 10 22
rect 3 17 4 21
rect 8 17 10 21
rect 3 16 10 17
rect 5 13 10 16
rect 12 29 20 30
rect 12 25 14 29
rect 18 25 20 29
rect 12 13 20 25
rect 22 21 30 30
rect 22 17 24 21
rect 28 17 30 21
rect 22 13 30 17
rect 32 18 40 30
rect 32 14 34 18
rect 38 14 40 18
rect 32 13 40 14
rect 42 21 50 30
rect 42 17 44 21
rect 48 17 50 21
rect 42 13 50 17
rect 52 13 62 30
rect 64 22 69 30
rect 64 21 71 22
rect 64 17 66 21
rect 70 17 71 21
rect 64 16 71 17
rect 64 13 69 16
rect 54 12 60 13
rect 54 8 55 12
rect 59 8 60 12
rect 54 7 60 8
<< pdiffusion >>
rect 27 63 32 67
rect 14 62 22 63
rect 14 61 15 62
rect 4 55 9 61
rect 2 54 9 55
rect 2 50 3 54
rect 7 50 9 54
rect 2 47 9 50
rect 2 43 3 47
rect 7 43 9 47
rect 2 42 9 43
rect 11 58 15 61
rect 19 58 22 62
rect 11 55 22 58
rect 11 51 15 55
rect 19 51 22 55
rect 11 42 22 51
rect 24 54 32 63
rect 24 50 26 54
rect 30 50 32 54
rect 24 47 32 50
rect 24 43 26 47
rect 30 43 32 47
rect 24 42 32 43
rect 34 42 39 67
rect 41 66 49 67
rect 41 62 43 66
rect 47 62 49 66
rect 41 42 49 62
rect 51 42 56 67
rect 58 62 66 67
rect 58 58 60 62
rect 64 58 66 62
rect 58 55 66 58
rect 58 51 60 55
rect 64 51 66 55
rect 58 42 66 51
rect 68 42 73 67
rect 75 66 82 67
rect 75 62 77 66
rect 81 62 82 66
rect 75 59 82 62
rect 75 55 77 59
rect 81 55 82 59
rect 75 42 82 55
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect -2 68 90 78
rect 14 62 20 68
rect 14 58 15 62
rect 19 58 20 62
rect 43 66 47 68
rect 77 66 81 68
rect 43 61 47 62
rect 58 62 64 63
rect 14 55 20 58
rect 2 54 7 55
rect 2 50 3 54
rect 14 51 15 55
rect 19 51 20 55
rect 58 58 60 62
rect 58 55 64 58
rect 58 54 60 55
rect 2 47 7 50
rect 25 50 26 54
rect 30 51 60 54
rect 77 59 81 62
rect 77 54 81 55
rect 64 51 71 54
rect 30 50 71 51
rect 25 47 30 50
rect 2 43 3 47
rect 7 43 26 47
rect 18 42 30 43
rect 34 42 71 46
rect 2 38 14 39
rect 2 34 10 38
rect 2 33 14 34
rect 2 25 6 33
rect 13 25 14 29
rect 18 25 22 42
rect 29 34 30 38
rect 34 34 39 42
rect 59 38 65 42
rect 46 34 47 38
rect 51 34 55 38
rect 59 34 60 38
rect 64 34 65 38
rect 73 34 74 38
rect 78 34 79 38
rect 49 30 55 34
rect 73 30 79 34
rect 26 23 46 27
rect 49 26 79 30
rect 26 21 30 23
rect 3 17 4 21
rect 8 17 24 21
rect 28 17 30 21
rect 42 21 46 23
rect 34 18 38 19
rect 42 17 44 21
rect 48 17 66 21
rect 70 17 71 21
rect 34 12 38 14
rect -2 8 55 12
rect 59 8 90 12
rect -2 2 90 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
<< ntransistor >>
rect 10 13 12 30
rect 20 13 22 30
rect 30 13 32 30
rect 40 13 42 30
rect 50 13 52 30
rect 62 13 64 30
<< ptransistor >>
rect 9 42 11 61
rect 22 42 24 63
rect 32 42 34 67
rect 39 42 41 67
rect 49 42 51 67
rect 56 42 58 67
rect 66 42 68 67
rect 73 42 75 67
<< polycontact >>
rect 10 34 14 38
rect 30 34 34 38
rect 47 34 51 38
rect 60 34 64 38
rect 74 34 78 38
<< ndcontact >>
rect 4 17 8 21
rect 14 25 18 29
rect 24 17 28 21
rect 34 14 38 18
rect 44 17 48 21
rect 66 17 70 21
rect 55 8 59 12
<< pdcontact >>
rect 3 50 7 54
rect 3 43 7 47
rect 15 58 19 62
rect 15 51 19 55
rect 26 50 30 54
rect 26 43 30 47
rect 43 62 47 66
rect 60 58 64 62
rect 60 51 64 55
rect 77 62 81 66
rect 77 55 81 59
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
<< psubstratepdiff >>
rect 0 2 88 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 88 2
rect 0 -3 88 -2
<< nsubstratendiff >>
rect 0 82 88 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 88 82
rect 0 77 88 78
<< labels >>
rlabel metal1 4 32 4 32 6 b
rlabel polycontact 12 36 12 36 6 b
rlabel pdcontact 4 52 4 52 6 z
rlabel metal1 16 19 16 19 6 n1
rlabel metal1 20 36 20 36 6 z
rlabel pdcontact 28 52 28 52 6 z
rlabel metal1 44 6 44 6 6 vss
rlabel metal1 36 36 36 36 6 a2
rlabel metal1 44 44 44 44 6 a2
rlabel metal1 44 52 44 52 6 z
rlabel metal1 36 52 36 52 6 z
rlabel metal1 44 74 44 74 6 vdd
rlabel metal1 60 28 60 28 6 a1
rlabel metal1 68 28 68 28 6 a1
rlabel metal1 52 32 52 32 6 a1
rlabel metal1 52 44 52 44 6 a2
rlabel metal1 60 44 60 44 6 a2
rlabel metal1 68 44 68 44 6 a2
rlabel metal1 68 52 68 52 6 z
rlabel metal1 52 52 52 52 6 z
rlabel metal1 60 56 60 56 6 z
rlabel metal1 56 19 56 19 6 n1
rlabel metal1 76 32 76 32 6 a1
<< end >>
