magic
tech scmos
timestamp 1179386503
<< checkpaint >>
rect -22 -22 78 94
<< ab >>
rect 0 0 56 72
<< pwell >>
rect -4 -4 60 32
<< nwell >>
rect -4 32 60 76
<< polysilicon >>
rect 9 59 11 65
rect 19 59 21 65
rect 31 57 33 61
rect 41 57 43 61
rect 9 35 11 40
rect 19 37 21 40
rect 31 37 33 40
rect 19 36 33 37
rect 9 34 15 35
rect 9 30 10 34
rect 14 30 15 34
rect 9 29 15 30
rect 19 32 26 36
rect 30 35 33 36
rect 41 35 43 40
rect 30 32 31 35
rect 19 31 31 32
rect 41 34 47 35
rect 41 31 42 34
rect 12 26 14 29
rect 19 26 21 31
rect 29 26 31 31
rect 36 30 42 31
rect 46 30 47 34
rect 36 29 47 30
rect 36 26 38 29
rect 12 4 14 9
rect 19 4 21 9
rect 29 8 31 13
rect 36 8 38 13
<< ndiffusion >>
rect 3 9 12 26
rect 14 9 19 26
rect 21 18 29 26
rect 21 14 23 18
rect 27 14 29 18
rect 21 13 29 14
rect 31 13 36 26
rect 38 18 46 26
rect 38 14 40 18
rect 44 14 46 18
rect 38 13 46 14
rect 21 9 26 13
rect 3 8 10 9
rect 3 4 5 8
rect 9 4 10 8
rect 3 3 10 4
<< pdiffusion >>
rect 2 58 9 59
rect 2 54 3 58
rect 7 54 9 58
rect 2 51 9 54
rect 2 47 3 51
rect 7 47 9 51
rect 2 40 9 47
rect 11 52 19 59
rect 11 48 13 52
rect 17 48 19 52
rect 11 45 19 48
rect 11 41 13 45
rect 17 41 19 45
rect 11 40 19 41
rect 21 58 29 59
rect 21 54 24 58
rect 28 57 29 58
rect 28 54 31 57
rect 21 40 31 54
rect 33 56 41 57
rect 33 52 35 56
rect 39 52 41 56
rect 33 49 41 52
rect 33 45 35 49
rect 39 45 41 49
rect 33 40 41 45
rect 43 56 50 57
rect 43 52 45 56
rect 49 52 50 56
rect 43 49 50 52
rect 43 45 45 49
rect 49 45 50 49
rect 43 40 50 45
<< metal1 >>
rect -2 68 58 72
rect -2 64 34 68
rect 38 64 44 68
rect 48 64 58 68
rect 2 58 8 64
rect 2 54 3 58
rect 7 54 8 58
rect 23 58 29 64
rect 23 54 24 58
rect 28 54 29 58
rect 34 56 40 59
rect 2 51 8 54
rect 2 47 3 51
rect 7 47 8 51
rect 13 52 17 54
rect 34 52 35 56
rect 39 52 40 56
rect 34 50 40 52
rect 17 49 40 50
rect 17 48 35 49
rect 13 46 35 48
rect 13 45 17 46
rect 34 45 35 46
rect 39 45 40 49
rect 44 56 50 64
rect 44 52 45 56
rect 49 52 50 56
rect 44 49 50 52
rect 44 45 45 49
rect 49 45 50 49
rect 2 41 13 43
rect 2 39 17 41
rect 2 18 6 39
rect 25 38 39 42
rect 25 36 31 38
rect 10 34 18 35
rect 14 30 18 34
rect 25 32 26 36
rect 30 32 31 36
rect 25 30 31 32
rect 41 30 42 34
rect 46 30 47 34
rect 10 29 18 30
rect 14 26 18 29
rect 41 26 47 30
rect 14 22 47 26
rect 2 14 23 18
rect 27 14 31 18
rect 39 14 40 18
rect 44 14 45 18
rect 39 8 45 14
rect -2 4 5 8
rect 9 4 45 8
rect 49 4 58 8
rect -2 0 58 4
<< ntransistor >>
rect 12 9 14 26
rect 19 9 21 26
rect 29 13 31 26
rect 36 13 38 26
<< ptransistor >>
rect 9 40 11 59
rect 19 40 21 59
rect 31 40 33 57
rect 41 40 43 57
<< polycontact >>
rect 10 30 14 34
rect 26 32 30 36
rect 42 30 46 34
<< ndcontact >>
rect 23 14 27 18
rect 40 14 44 18
rect 5 4 9 8
<< pdcontact >>
rect 3 54 7 58
rect 3 47 7 51
rect 13 48 17 52
rect 13 41 17 45
rect 24 54 28 58
rect 35 52 39 56
rect 35 45 39 49
rect 45 52 49 56
rect 45 45 49 49
<< psubstratepcontact >>
rect 45 4 49 8
<< nsubstratencontact >>
rect 34 64 38 68
rect 44 64 48 68
<< psubstratepdiff >>
rect 44 8 50 9
rect 44 4 45 8
rect 49 4 50 8
rect 44 3 50 4
<< nsubstratendiff >>
rect 33 68 49 69
rect 33 64 34 68
rect 38 64 44 68
rect 48 64 49 68
rect 33 63 49 64
<< labels >>
rlabel metal1 4 32 4 32 6 z
rlabel metal1 20 16 20 16 6 z
rlabel metal1 12 16 12 16 6 z
rlabel polycontact 12 32 12 32 6 a
rlabel metal1 20 24 20 24 6 a
rlabel metal1 20 48 20 48 6 z
rlabel metal1 28 4 28 4 6 vss
rlabel metal1 28 16 28 16 6 z
rlabel metal1 28 24 28 24 6 a
rlabel metal1 36 24 36 24 6 a
rlabel metal1 36 40 36 40 6 b
rlabel metal1 28 36 28 36 6 b
rlabel metal1 28 48 28 48 6 z
rlabel metal1 36 52 36 52 6 z
rlabel metal1 28 68 28 68 6 vdd
rlabel metal1 44 28 44 28 6 a
<< end >>
