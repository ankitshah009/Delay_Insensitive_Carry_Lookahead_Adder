magic
tech scmos
timestamp 1179386188
<< checkpaint >>
rect -22 -25 78 105
<< ab >>
rect 0 0 56 80
<< pwell >>
rect -4 -7 60 36
<< nwell >>
rect -4 36 60 87
<< polysilicon >>
rect 22 68 24 73
rect 32 68 34 73
rect 45 70 47 74
rect 9 61 11 65
rect 45 49 47 52
rect 41 48 47 49
rect 41 44 42 48
rect 46 44 47 48
rect 9 31 11 43
rect 22 41 24 44
rect 16 40 24 41
rect 16 36 17 40
rect 21 36 24 40
rect 32 41 34 44
rect 41 43 47 44
rect 32 39 37 41
rect 16 35 24 36
rect 35 38 41 39
rect 22 33 30 35
rect 9 30 16 31
rect 28 30 30 33
rect 35 34 36 38
rect 40 34 41 38
rect 35 33 41 34
rect 35 30 37 33
rect 45 30 47 43
rect 9 26 11 30
rect 15 26 16 30
rect 9 25 16 26
rect 9 22 11 25
rect 9 8 11 13
rect 45 16 47 21
rect 28 6 30 10
rect 35 6 37 10
<< ndiffusion >>
rect 21 29 28 30
rect 21 25 22 29
rect 26 25 28 29
rect 21 24 28 25
rect 2 21 9 22
rect 2 17 3 21
rect 7 17 9 21
rect 2 16 9 17
rect 4 13 9 16
rect 11 20 17 22
rect 11 13 19 20
rect 13 12 19 13
rect 13 8 14 12
rect 18 8 19 12
rect 23 10 28 24
rect 30 10 35 30
rect 37 26 45 30
rect 37 22 39 26
rect 43 22 45 26
rect 37 21 45 22
rect 47 29 54 30
rect 47 25 49 29
rect 53 25 54 29
rect 47 24 54 25
rect 47 21 52 24
rect 37 10 43 21
rect 13 7 19 8
<< pdiffusion >>
rect 36 69 45 70
rect 36 68 37 69
rect 14 62 22 68
rect 14 61 15 62
rect 4 56 9 61
rect 2 55 9 56
rect 2 51 3 55
rect 7 51 9 55
rect 2 48 9 51
rect 2 44 3 48
rect 7 44 9 48
rect 2 43 9 44
rect 11 58 15 61
rect 19 58 22 62
rect 11 44 22 58
rect 24 57 32 68
rect 24 53 26 57
rect 30 53 32 57
rect 24 49 32 53
rect 24 45 26 49
rect 30 45 32 49
rect 24 44 32 45
rect 34 65 37 68
rect 41 65 45 69
rect 34 62 45 65
rect 34 58 37 62
rect 41 58 45 62
rect 34 52 45 58
rect 47 58 52 70
rect 47 57 54 58
rect 47 53 49 57
rect 53 53 54 57
rect 47 52 54 53
rect 34 44 39 52
rect 11 43 16 44
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect -2 69 58 78
rect -2 68 37 69
rect 14 62 20 68
rect 14 58 15 62
rect 19 58 20 62
rect 36 65 37 68
rect 41 68 58 69
rect 41 65 42 68
rect 36 62 42 65
rect 36 58 37 62
rect 41 58 42 62
rect 26 57 30 58
rect 3 55 7 56
rect 3 48 7 51
rect 17 53 26 54
rect 49 57 53 58
rect 17 50 30 53
rect 3 40 7 44
rect 26 49 30 50
rect 34 49 46 55
rect 2 36 17 40
rect 21 36 22 40
rect 2 21 6 36
rect 26 30 30 45
rect 42 48 46 49
rect 42 41 46 44
rect 49 38 53 53
rect 35 34 36 38
rect 40 34 53 38
rect 9 26 11 30
rect 15 26 18 30
rect 14 22 18 26
rect 21 29 30 30
rect 21 25 22 29
rect 26 26 30 29
rect 49 29 53 34
rect 39 26 43 27
rect 26 25 27 26
rect 49 24 53 25
rect 2 17 3 21
rect 7 17 8 21
rect 14 18 31 22
rect 39 12 43 22
rect -2 8 14 12
rect 18 8 58 12
rect -2 2 58 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
<< ntransistor >>
rect 9 13 11 22
rect 28 10 30 30
rect 35 10 37 30
rect 45 21 47 30
<< ptransistor >>
rect 9 43 11 61
rect 22 44 24 68
rect 32 44 34 68
rect 45 52 47 70
<< polycontact >>
rect 42 44 46 48
rect 17 36 21 40
rect 36 34 40 38
rect 11 26 15 30
<< ndcontact >>
rect 22 25 26 29
rect 3 17 7 21
rect 14 8 18 12
rect 39 22 43 26
rect 49 25 53 29
<< pdcontact >>
rect 3 51 7 55
rect 3 44 7 48
rect 15 58 19 62
rect 26 53 30 57
rect 26 45 30 49
rect 37 65 41 69
rect 37 58 41 62
rect 49 53 53 57
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
<< psubstratepdiff >>
rect 0 2 56 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 56 2
rect 0 -3 56 -2
<< nsubstratendiff >>
rect 0 82 56 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 56 82
rect 0 77 56 78
<< labels >>
rlabel polycontact 20 38 20 38 6 bn
rlabel polycontact 38 36 38 36 6 an
rlabel pdcontact 5 46 5 46 6 bn
rlabel metal1 4 28 4 28 6 bn
rlabel metal1 20 20 20 20 6 b
rlabel polycontact 12 28 12 28 6 b
rlabel metal1 12 38 12 38 6 bn
rlabel metal1 20 52 20 52 6 z
rlabel metal1 28 6 28 6 6 vss
rlabel metal1 28 20 28 20 6 b
rlabel metal1 28 44 28 44 6 z
rlabel metal1 36 52 36 52 6 a
rlabel metal1 28 74 28 74 6 vdd
rlabel metal1 44 36 44 36 6 an
rlabel metal1 51 41 51 41 6 an
rlabel metal1 44 48 44 48 6 a
<< end >>
