.subckt noa2a22_x4 i0 i1 i2 i3 nq vdd vss
*   SPICE3 file   created from noa2a22_x4.ext -      technology: scmos
m00 w1     i0     w2     vdd p w=20u  l=2.3636u ad=100p     pd=30u      as=130p     ps=43u
m01 w2     i1     w1     vdd p w=20u  l=2.3636u ad=130p     pd=43u      as=100p     ps=30u
m02 vdd    i3     w2     vdd p w=20u  l=2.3636u ad=132.571p pd=38.8571u as=130p     ps=43u
m03 w2     i2     vdd    vdd p w=20u  l=2.3636u ad=130p     pd=43u      as=132.571p ps=38.8571u
m04 vdd    w1     w3     vdd p w=20u  l=2.3636u ad=132.571p pd=38.8571u as=160p     ps=56u
m05 nq     w3     vdd    vdd p w=40u  l=2.3636u ad=200p     pd=50u      as=265.143p ps=77.7143u
m06 vdd    w3     nq     vdd p w=40u  l=2.3636u ad=265.143p pd=77.7143u as=200p     ps=50u
m07 w4     i0     vss    vss n w=10u  l=2.3636u ad=50p      pd=20u      as=85.1429p ps=31.4286u
m08 w1     i1     w4     vss n w=10u  l=2.3636u ad=50p      pd=20u      as=50p      ps=20u
m09 w5     i3     w1     vss n w=10u  l=2.3636u ad=50p      pd=20u      as=50p      ps=20u
m10 vss    i2     w5     vss n w=10u  l=2.3636u ad=85.1429p pd=31.4286u as=50p      ps=20u
m11 vss    w1     w3     vss n w=10u  l=2.3636u ad=85.1429p pd=31.4286u as=80p      ps=36u
m12 nq     w3     vss    vss n w=20u  l=2.3636u ad=100p     pd=30u      as=170.286p ps=62.8571u
m13 vss    w3     nq     vss n w=20u  l=2.3636u ad=170.286p pd=62.8571u as=100p     ps=30u
C0  nq     w1     0.087f
C1  w5     i3     0.016f
C2  i1     w3     0.033f
C3  i3     vdd    0.010f
C4  w4     i1     0.016f
C5  w1     w2     0.289f
C6  vss    i3     0.047f
C7  nq     i2     0.039f
C8  i0     vdd    0.010f
C9  vss    i0     0.051f
C10 w2     i2     0.017f
C11 w1     i3     0.342f
C12 w2     i1     0.017f
C13 i2     i3     0.425f
C14 w1     i0     0.090f
C15 nq     w3     0.132f
C16 vss    vdd    0.005f
C17 w1     vdd    0.229f
C18 i2     i0     0.062f
C19 i3     i1     0.172f
C20 vss    w1     0.064f
C21 w5     i2     0.004f
C22 i3     w3     0.069f
C23 i2     vdd    0.010f
C24 i1     i0     0.425f
C25 vss    i2     0.058f
C26 nq     w2     0.006f
C27 i1     vdd    0.011f
C28 w1     i2     0.173f
C29 w4     i0     0.004f
C30 vss    i1     0.042f
C31 w3     vdd    0.031f
C32 w2     i3     0.017f
C33 w1     i1     0.314f
C34 vss    w3     0.116f
C35 i2     i1     0.090f
C36 w2     i0     0.017f
C37 w1     w3     0.349f
C38 nq     vdd    0.231f
C39 vss    nq     0.130f
C40 w2     vdd    0.409f
C41 i2     w3     0.142f
C42 i3     i0     0.090f
C44 nq     vss    0.018f
C45 w1     vss    0.046f
C46 i2     vss    0.040f
C47 i3     vss    0.050f
C48 i1     vss    0.050f
C49 i0     vss    0.040f
C50 w3     vss    0.069f
.ends
