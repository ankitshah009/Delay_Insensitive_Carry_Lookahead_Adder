magic
tech scmos
timestamp 1179387279
<< checkpaint >>
rect -22 -22 110 94
<< ab >>
rect 0 0 88 72
<< pwell >>
rect -4 -4 92 32
<< nwell >>
rect -4 32 92 76
<< polysilicon >>
rect 21 64 23 69
rect 28 64 30 69
rect 35 64 37 69
rect 42 64 44 69
rect 52 64 54 69
rect 59 64 61 69
rect 66 64 68 69
rect 73 64 75 69
rect 9 56 11 61
rect 21 41 23 46
rect 18 40 24 41
rect 9 30 11 38
rect 18 36 19 40
rect 23 36 24 40
rect 18 35 24 36
rect 9 29 15 30
rect 9 25 10 29
rect 14 25 15 29
rect 9 24 15 25
rect 9 21 11 24
rect 21 18 23 35
rect 28 31 30 46
rect 35 37 37 46
rect 42 43 44 46
rect 52 43 54 46
rect 42 42 55 43
rect 42 41 50 42
rect 49 38 50 41
rect 54 38 55 42
rect 49 37 55 38
rect 35 35 45 37
rect 28 30 39 31
rect 28 29 34 30
rect 31 26 34 29
rect 38 26 39 30
rect 31 25 39 26
rect 43 27 45 35
rect 43 26 49 27
rect 31 18 33 25
rect 43 22 44 26
rect 48 22 49 26
rect 43 21 49 22
rect 43 18 45 21
rect 53 18 55 37
rect 59 27 61 46
rect 66 37 68 46
rect 73 43 75 46
rect 73 42 81 43
rect 73 41 76 42
rect 75 38 76 41
rect 80 38 81 42
rect 75 37 81 38
rect 65 36 71 37
rect 65 32 66 36
rect 70 32 71 36
rect 65 31 71 32
rect 59 26 65 27
rect 59 22 60 26
rect 64 22 65 26
rect 59 21 65 22
rect 9 7 11 12
rect 21 7 23 12
rect 31 7 33 12
rect 43 7 45 12
rect 53 7 55 12
<< ndiffusion >>
rect 4 18 9 21
rect 2 17 9 18
rect 2 13 3 17
rect 7 13 9 17
rect 2 12 9 13
rect 11 18 19 21
rect 11 12 21 18
rect 23 17 31 18
rect 23 13 25 17
rect 29 13 31 17
rect 23 12 31 13
rect 33 12 43 18
rect 45 17 53 18
rect 45 13 47 17
rect 51 13 53 17
rect 45 12 53 13
rect 55 12 63 18
rect 13 8 19 12
rect 13 4 14 8
rect 18 4 19 8
rect 35 8 41 12
rect 13 3 19 4
rect 35 4 36 8
rect 40 4 41 8
rect 57 8 63 12
rect 35 3 41 4
rect 57 4 58 8
rect 62 4 63 8
rect 57 3 63 4
<< pdiffusion >>
rect 13 65 19 66
rect 13 61 14 65
rect 18 64 19 65
rect 18 61 21 64
rect 13 56 21 61
rect 4 51 9 56
rect 2 50 9 51
rect 2 46 3 50
rect 7 46 9 50
rect 2 43 9 46
rect 2 39 3 43
rect 7 39 9 43
rect 2 38 9 39
rect 11 46 21 56
rect 23 46 28 64
rect 30 46 35 64
rect 37 46 42 64
rect 44 58 52 64
rect 44 54 46 58
rect 50 54 52 58
rect 44 46 52 54
rect 54 46 59 64
rect 61 46 66 64
rect 68 46 73 64
rect 75 63 82 64
rect 75 59 77 63
rect 81 59 82 63
rect 75 46 82 59
rect 11 38 16 46
<< metal1 >>
rect -2 68 90 72
rect -2 64 4 68
rect 8 65 90 68
rect 8 64 14 65
rect 13 61 14 64
rect 18 64 90 65
rect 18 61 19 64
rect 77 63 81 64
rect 2 51 6 59
rect 10 54 46 58
rect 50 54 51 58
rect 2 50 7 51
rect 2 46 3 50
rect 2 43 7 46
rect 2 39 3 43
rect 2 38 7 39
rect 2 18 6 38
rect 10 29 14 54
rect 58 50 62 59
rect 77 58 81 59
rect 18 46 81 50
rect 18 40 23 46
rect 75 42 81 46
rect 18 36 19 40
rect 18 35 23 36
rect 26 38 50 42
rect 54 38 55 42
rect 26 29 30 38
rect 65 36 71 42
rect 75 38 76 42
rect 80 38 81 42
rect 65 34 66 36
rect 34 32 66 34
rect 70 32 71 36
rect 34 30 71 32
rect 14 25 23 28
rect 10 24 23 25
rect 2 17 16 18
rect 2 13 3 17
rect 7 13 16 17
rect 19 17 23 24
rect 34 21 38 26
rect 43 22 44 26
rect 48 22 60 26
rect 64 22 65 26
rect 19 13 25 17
rect 29 13 47 17
rect 51 13 52 17
rect 58 13 62 22
rect -2 4 14 8
rect 18 4 36 8
rect 40 4 58 8
rect 62 4 68 8
rect 72 4 76 8
rect 80 4 90 8
rect -2 0 90 4
<< ntransistor >>
rect 9 12 11 21
rect 21 12 23 18
rect 31 12 33 18
rect 43 12 45 18
rect 53 12 55 18
<< ptransistor >>
rect 9 38 11 56
rect 21 46 23 64
rect 28 46 30 64
rect 35 46 37 64
rect 42 46 44 64
rect 52 46 54 64
rect 59 46 61 64
rect 66 46 68 64
rect 73 46 75 64
<< polycontact >>
rect 19 36 23 40
rect 10 25 14 29
rect 50 38 54 42
rect 34 26 38 30
rect 44 22 48 26
rect 76 38 80 42
rect 66 32 70 36
rect 60 22 64 26
<< ndcontact >>
rect 3 13 7 17
rect 25 13 29 17
rect 47 13 51 17
rect 14 4 18 8
rect 36 4 40 8
rect 58 4 62 8
<< pdcontact >>
rect 14 61 18 65
rect 3 46 7 50
rect 3 39 7 43
rect 46 54 50 58
rect 77 59 81 63
<< psubstratepcontact >>
rect 68 4 72 8
rect 76 4 80 8
<< nsubstratencontact >>
rect 4 64 8 68
<< psubstratepdiff >>
rect 67 8 81 24
rect 67 4 68 8
rect 72 4 76 8
rect 80 4 81 8
rect 67 3 81 4
<< nsubstratendiff >>
rect 3 68 9 69
rect 3 64 4 68
rect 8 64 9 68
rect 3 63 9 64
<< labels >>
rlabel polycontact 12 27 12 27 6 zn
rlabel metal1 12 16 12 16 6 z
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 41 12 41 6 zn
rlabel metal1 28 32 28 32 6 d
rlabel metal1 20 40 20 40 6 a
rlabel metal1 28 48 28 48 6 a
rlabel metal1 44 4 44 4 6 vss
rlabel metal1 35 15 35 15 6 zn
rlabel metal1 36 24 36 24 6 b
rlabel metal1 44 32 44 32 6 b
rlabel metal1 36 40 36 40 6 d
rlabel metal1 44 40 44 40 6 d
rlabel metal1 36 48 36 48 6 a
rlabel metal1 44 48 44 48 6 a
rlabel metal1 30 56 30 56 6 zn
rlabel metal1 44 68 44 68 6 vdd
rlabel metal1 52 24 52 24 6 c
rlabel metal1 60 20 60 20 6 c
rlabel metal1 60 32 60 32 6 b
rlabel metal1 52 32 52 32 6 b
rlabel polycontact 52 40 52 40 6 d
rlabel metal1 68 36 68 36 6 b
rlabel metal1 52 48 52 48 6 a
rlabel metal1 60 52 60 52 6 a
rlabel metal1 68 48 68 48 6 a
rlabel metal1 76 48 76 48 6 a
<< end >>
