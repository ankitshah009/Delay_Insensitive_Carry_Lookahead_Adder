magic
tech scmos
timestamp 1179386557
<< checkpaint >>
rect -22 -25 94 105
<< ab >>
rect 0 0 72 80
<< pwell >>
rect -4 -7 76 36
<< nwell >>
rect -4 36 76 87
<< polysilicon >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 39 70 41 74
rect 49 70 51 74
rect 59 70 61 74
rect 9 39 11 50
rect 19 47 21 50
rect 19 46 25 47
rect 19 42 20 46
rect 24 42 25 46
rect 19 41 25 42
rect 9 38 15 39
rect 9 34 10 38
rect 14 36 15 38
rect 14 34 16 36
rect 9 33 16 34
rect 14 30 16 33
rect 21 30 23 41
rect 29 39 31 50
rect 39 39 41 50
rect 49 47 51 50
rect 29 38 41 39
rect 29 36 32 38
rect 28 34 32 36
rect 36 34 41 38
rect 28 33 41 34
rect 45 46 51 47
rect 45 42 46 46
rect 50 42 51 46
rect 45 41 51 42
rect 28 30 30 33
rect 38 30 40 33
rect 45 30 47 41
rect 59 39 61 50
rect 55 38 61 39
rect 55 36 56 38
rect 52 34 56 36
rect 60 34 61 38
rect 52 33 61 34
rect 52 30 54 33
rect 14 6 16 10
rect 21 6 23 10
rect 28 6 30 10
rect 38 6 40 10
rect 45 6 47 10
rect 52 6 54 10
<< ndiffusion >>
rect 6 15 14 30
rect 6 11 8 15
rect 12 11 14 15
rect 6 10 14 11
rect 16 10 21 30
rect 23 10 28 30
rect 30 22 38 30
rect 30 18 32 22
rect 36 18 38 22
rect 30 10 38 18
rect 40 10 45 30
rect 47 10 52 30
rect 54 29 62 30
rect 54 25 56 29
rect 60 25 62 29
rect 54 22 62 25
rect 54 18 56 22
rect 60 18 62 22
rect 54 17 62 18
rect 54 10 59 17
<< pdiffusion >>
rect 2 69 9 70
rect 2 65 3 69
rect 7 65 9 69
rect 2 62 9 65
rect 2 58 3 62
rect 7 58 9 62
rect 2 50 9 58
rect 11 62 19 70
rect 11 58 13 62
rect 17 58 19 62
rect 11 55 19 58
rect 11 51 13 55
rect 17 51 19 55
rect 11 50 19 51
rect 21 69 29 70
rect 21 65 23 69
rect 27 65 29 69
rect 21 62 29 65
rect 21 58 23 62
rect 27 58 29 62
rect 21 50 29 58
rect 31 62 39 70
rect 31 58 33 62
rect 37 58 39 62
rect 31 55 39 58
rect 31 51 33 55
rect 37 51 39 55
rect 31 50 39 51
rect 41 69 49 70
rect 41 65 43 69
rect 47 65 49 69
rect 41 50 49 65
rect 51 62 59 70
rect 51 58 53 62
rect 57 58 59 62
rect 51 55 59 58
rect 51 51 53 55
rect 57 51 59 55
rect 51 50 59 51
rect 61 69 68 70
rect 61 65 63 69
rect 67 65 68 69
rect 61 62 68 65
rect 61 58 63 62
rect 67 58 68 62
rect 61 50 68 58
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect -2 69 74 78
rect -2 68 3 69
rect 2 65 3 68
rect 7 68 23 69
rect 7 65 8 68
rect 2 62 8 65
rect 22 65 23 68
rect 27 68 43 69
rect 27 65 28 68
rect 42 65 43 68
rect 47 68 63 69
rect 47 65 48 68
rect 62 65 63 68
rect 67 68 74 69
rect 67 65 68 68
rect 2 58 3 62
rect 7 58 8 62
rect 13 62 17 63
rect 22 62 28 65
rect 62 62 68 65
rect 22 58 23 62
rect 27 58 28 62
rect 32 58 33 62
rect 37 58 53 62
rect 57 58 58 62
rect 62 58 63 62
rect 67 58 68 62
rect 13 55 17 58
rect 2 51 13 54
rect 32 55 37 58
rect 32 54 33 55
rect 17 51 33 54
rect 53 55 58 58
rect 2 50 37 51
rect 2 22 6 50
rect 41 46 47 54
rect 57 54 58 55
rect 57 51 63 54
rect 53 50 63 51
rect 19 42 20 46
rect 24 42 46 46
rect 50 42 55 46
rect 10 38 14 39
rect 25 34 32 38
rect 36 34 39 38
rect 44 34 56 38
rect 60 34 63 38
rect 10 30 14 34
rect 44 30 48 34
rect 10 26 48 30
rect 2 18 32 22
rect 36 18 37 22
rect 42 17 46 26
rect 55 25 56 29
rect 60 25 61 29
rect 55 22 61 25
rect 55 18 56 22
rect 60 18 61 22
rect 7 12 8 15
rect -2 11 8 12
rect 12 12 13 15
rect 55 12 61 18
rect 12 11 74 12
rect -2 2 74 11
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
<< ntransistor >>
rect 14 10 16 30
rect 21 10 23 30
rect 28 10 30 30
rect 38 10 40 30
rect 45 10 47 30
rect 52 10 54 30
<< ptransistor >>
rect 9 50 11 70
rect 19 50 21 70
rect 29 50 31 70
rect 39 50 41 70
rect 49 50 51 70
rect 59 50 61 70
<< polycontact >>
rect 20 42 24 46
rect 10 34 14 38
rect 32 34 36 38
rect 46 42 50 46
rect 56 34 60 38
<< ndcontact >>
rect 8 11 12 15
rect 32 18 36 22
rect 56 25 60 29
rect 56 18 60 22
<< pdcontact >>
rect 3 65 7 69
rect 3 58 7 62
rect 13 58 17 62
rect 13 51 17 55
rect 23 65 27 69
rect 23 58 27 62
rect 33 58 37 62
rect 33 51 37 55
rect 43 65 47 69
rect 53 58 57 62
rect 53 51 57 55
rect 63 65 67 69
rect 63 58 67 62
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
<< psubstratepdiff >>
rect 0 2 72 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 72 2
rect 0 -3 72 -2
<< nsubstratendiff >>
rect 0 82 72 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 72 82
rect 0 77 72 78
<< labels >>
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 20 12 20 6 z
rlabel metal1 20 20 20 20 6 z
rlabel metal1 20 28 20 28 6 a
rlabel polycontact 12 36 12 36 6 a
rlabel metal1 20 52 20 52 6 z
rlabel metal1 12 52 12 52 6 z
rlabel metal1 36 6 36 6 6 vss
rlabel metal1 28 20 28 20 6 z
rlabel metal1 28 28 28 28 6 a
rlabel metal1 36 28 36 28 6 a
rlabel metal1 28 36 28 36 6 c
rlabel metal1 28 44 28 44 6 b
rlabel metal1 36 36 36 36 6 c
rlabel metal1 36 44 36 44 6 b
rlabel metal1 28 52 28 52 6 z
rlabel pdcontact 36 60 36 60 6 z
rlabel metal1 36 74 36 74 6 vdd
rlabel metal1 44 24 44 24 6 a
rlabel metal1 52 36 52 36 6 a
rlabel metal1 52 44 52 44 6 b
rlabel metal1 44 48 44 48 6 b
rlabel metal1 44 60 44 60 6 z
rlabel metal1 52 60 52 60 6 z
rlabel metal1 60 36 60 36 6 a
rlabel metal1 60 52 60 52 6 z
<< end >>
