magic
tech scmos
timestamp 1179386296
<< checkpaint >>
rect -22 -25 54 105
<< ab >>
rect 0 0 32 80
<< pwell >>
rect -4 -7 36 36
<< nwell >>
rect -4 36 36 87
<< polysilicon >>
rect 10 61 12 66
rect 20 61 22 65
rect 10 39 12 47
rect 9 38 15 39
rect 9 34 10 38
rect 14 34 15 38
rect 9 33 15 34
rect 9 23 11 33
rect 20 32 22 47
rect 20 31 26 32
rect 20 28 21 31
rect 16 27 21 28
rect 25 27 26 31
rect 16 26 26 27
rect 16 23 18 26
rect 9 6 11 11
rect 16 6 18 11
<< ndiffusion >>
rect 2 22 9 23
rect 2 18 3 22
rect 7 18 9 22
rect 2 17 9 18
rect 4 11 9 17
rect 11 11 16 23
rect 18 16 30 23
rect 18 12 25 16
rect 29 12 30 16
rect 18 11 30 12
<< pdiffusion >>
rect 2 62 8 63
rect 2 58 3 62
rect 7 61 8 62
rect 7 58 10 61
rect 2 47 10 58
rect 12 60 20 61
rect 12 56 14 60
rect 18 56 20 60
rect 12 53 20 56
rect 12 49 14 53
rect 18 49 20 53
rect 12 47 20 49
rect 22 60 30 61
rect 22 56 25 60
rect 29 56 30 60
rect 22 53 30 56
rect 22 49 25 53
rect 29 49 30 53
rect 22 47 30 49
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect -2 68 34 78
rect 2 62 8 68
rect 2 58 3 62
rect 7 58 8 62
rect 24 60 30 68
rect 13 56 14 60
rect 18 56 19 60
rect 13 54 19 56
rect 2 53 19 54
rect 2 49 14 53
rect 18 49 19 53
rect 24 56 25 60
rect 29 56 30 60
rect 24 53 30 56
rect 24 49 25 53
rect 29 49 30 53
rect 2 23 6 49
rect 17 42 23 46
rect 10 38 23 42
rect 10 33 14 34
rect 18 27 21 31
rect 25 27 30 31
rect 18 25 30 27
rect 2 22 7 23
rect 2 18 3 22
rect 2 17 7 18
rect 18 17 22 25
rect 25 16 29 17
rect -2 2 34 12
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
<< ntransistor >>
rect 9 11 11 23
rect 16 11 18 23
<< ptransistor >>
rect 10 47 12 61
rect 20 47 22 61
<< polycontact >>
rect 10 34 14 38
rect 21 27 25 31
<< ndcontact >>
rect 3 18 7 22
rect 25 12 29 16
<< pdcontact >>
rect 3 58 7 62
rect 14 56 18 60
rect 14 49 18 53
rect 25 56 29 60
rect 25 49 29 53
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
<< psubstratepdiff >>
rect 0 2 32 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 32 2
rect 0 -3 32 -2
<< nsubstratendiff >>
rect 0 82 32 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 32 82
rect 0 77 32 78
<< labels >>
rlabel metal1 4 32 4 32 6 z
rlabel polycontact 12 36 12 36 6 b
rlabel metal1 12 52 12 52 6 z
rlabel metal1 16 6 16 6 6 vss
rlabel metal1 20 24 20 24 6 a
rlabel metal1 20 44 20 44 6 b
rlabel metal1 16 74 16 74 6 vdd
rlabel metal1 28 28 28 28 6 a
<< end >>
