magic
tech scmos
timestamp 1182081815
<< checkpaint >>
rect -25 -26 57 114
<< ab >>
rect 0 0 32 88
<< pwell >>
rect -7 -8 39 40
<< nwell >>
rect -7 40 39 96
<< polysilicon >>
rect 5 85 14 86
rect 5 81 6 85
rect 10 81 14 85
rect 5 80 14 81
rect 18 85 27 86
rect 18 81 22 85
rect 26 81 27 85
rect 18 80 27 81
rect 9 77 11 80
rect 21 77 23 80
rect 9 48 11 51
rect 21 48 23 51
rect 2 42 11 48
rect 15 42 30 48
rect 2 32 17 38
rect 21 32 30 38
rect 9 29 11 32
rect 21 29 23 32
rect 9 8 11 11
rect 21 8 23 11
rect 5 7 14 8
rect 5 3 6 7
rect 10 3 14 7
rect 5 2 14 3
rect 18 7 27 8
rect 18 3 22 7
rect 26 3 27 7
rect 18 2 27 3
<< ndiffusion >>
rect 2 11 9 29
rect 11 11 21 29
rect 23 11 30 29
<< pdiffusion >>
rect 2 51 9 77
rect 11 51 21 77
rect 23 51 30 77
<< metal1 >>
rect -2 86 2 90
rect 30 86 34 90
rect 2 82 6 85
rect -2 81 6 82
rect 10 81 22 85
rect 26 82 30 85
rect 26 81 34 82
rect -2 6 6 7
rect 2 3 6 6
rect 10 3 22 7
rect 26 6 34 7
rect 26 3 30 6
rect -2 -2 2 2
rect 30 -2 34 2
<< metal2 >>
rect -2 86 34 90
rect 2 82 30 86
rect -2 80 34 82
rect -2 6 34 8
rect 2 2 30 6
rect -2 -2 34 2
<< ntransistor >>
rect 9 11 11 29
rect 21 11 23 29
<< ptransistor >>
rect 9 51 11 77
rect 21 51 23 77
<< polycontact >>
rect 6 81 10 85
rect 22 81 26 85
rect 6 3 10 7
rect 22 3 26 7
<< m2contact >>
rect -2 82 2 86
rect 30 82 34 86
rect -2 2 2 6
rect 30 2 34 6
<< psubstratepcontact >>
rect -2 2 2 6
rect 30 2 34 6
<< nsubstratencontact >>
rect -2 82 2 86
rect 30 82 34 86
<< psubstratepdiff >>
rect -3 6 3 7
rect -3 2 -2 6
rect 2 2 3 6
rect 29 6 35 7
rect 29 2 30 6
rect 34 2 35 6
rect -3 0 3 2
rect 29 0 35 2
<< nsubstratendiff >>
rect -3 86 3 88
rect 29 86 35 88
rect -3 82 -2 86
rect 2 82 3 86
rect -3 81 3 82
rect 29 82 30 86
rect 34 82 35 86
rect 29 81 35 82
<< labels >>
rlabel metal2 16 4 16 4 6 vss
rlabel metal2 16 84 16 84 6 vdd
<< end >>
