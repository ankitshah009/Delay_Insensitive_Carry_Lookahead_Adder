.subckt oa2ao222_x2 i0 i1 i2 i3 i4 q vdd vss
*   SPICE3 file   created from oa2ao222_x2.ext -      technology: scmos
m00 vdd    i0     w1     vdd p w=29u  l=2.3636u ad=196.49p  pd=56.8163u as=193.123p ps=56.7391u
m01 w1     i1     vdd    vdd p w=29u  l=2.3636u ad=193.123p pd=56.7391u as=196.49p  ps=56.8163u
m02 w2     i4     w1     vdd p w=40u  l=2.3636u ad=200p     pd=50u      as=266.377p ps=78.2609u
m03 w3     i2     w2     vdd p w=40u  l=2.3636u ad=160p     pd=48u      as=200p     ps=50u
m04 w1     i3     w3     vdd p w=40u  l=2.3636u ad=266.377p pd=78.2609u as=160p     ps=48u
m05 q      w2     vdd    vdd p w=40u  l=2.3636u ad=320p     pd=96u      as=271.02p  ps=78.3673u
m06 w4     i0     vss    vss n w=18u  l=2.3636u ad=72p      pd=26u      as=168.387p ps=59.2258u
m07 w2     i1     w4     vss n w=18u  l=2.3636u ad=100.8p   pd=33.6u    as=72p      ps=26u
m08 w5     i4     w2     vss n w=12u  l=2.3636u ad=96p      pd=36u      as=67.2p    ps=22.4u
m09 vss    i2     w5     vss n w=12u  l=2.3636u ad=112.258p pd=39.4839u as=96p      ps=36u
m10 w5     i3     vss    vss n w=12u  l=2.3636u ad=96p      pd=36u      as=112.258p ps=39.4839u
m11 q      w2     vss    vss n w=20u  l=2.3636u ad=160p     pd=56u      as=187.097p ps=65.8064u
C0  vss    q      0.144f
C1  i0     w2     0.079f
C2  i1     i3     0.040f
C3  w1     i2     0.017f
C4  w5     i0     0.006f
C5  w4     i1     0.012f
C6  i1     i4     0.314f
C7  i0     i2     0.040f
C8  vdd    i3     0.012f
C9  w3     w1     0.016f
C10 w5     w2     0.087f
C11 vss    i0     0.063f
C12 vdd    i4     0.017f
C13 w2     i2     0.279f
C14 vss    w2     0.109f
C15 w5     i2     0.033f
C16 w1     i1     0.036f
C17 q      vdd    0.114f
C18 i3     i4     0.052f
C19 w5     vss    0.250f
C20 q      i3     0.044f
C21 i1     i0     0.398f
C22 vss    i2     0.036f
C23 w1     vdd    0.502f
C24 w3     w2     0.016f
C25 i1     w2     0.109f
C26 i0     vdd    0.023f
C27 w1     i3     0.029f
C28 w3     i2     0.012f
C29 i1     i2     0.057f
C30 w1     i4     0.086f
C31 vdd    w2     0.180f
C32 q      w1     0.010f
C33 vss    i1     0.013f
C34 w4     i0     0.009f
C35 vdd    i2     0.012f
C36 i0     i4     0.094f
C37 w2     i3     0.161f
C38 w5     i3     0.047f
C39 i3     i2     0.322f
C40 w2     i4     0.268f
C41 w1     i0     0.064f
C42 vss    i3     0.031f
C43 w3     vdd    0.019f
C44 q      w2     0.141f
C45 i2     i4     0.094f
C46 w5     q      0.012f
C47 w3     i3     0.004f
C48 i1     vdd    0.050f
C49 vss    i4     0.009f
C50 w1     w2     0.194f
C51 q      i2     0.031f
C52 w5     vss    0.005f
C54 q      vss    0.025f
C55 i1     vss    0.024f
C56 i0     vss    0.023f
C58 w2     vss    0.033f
C59 i3     vss    0.023f
C60 i2     vss    0.024f
C61 i4     vss    0.028f
.ends
