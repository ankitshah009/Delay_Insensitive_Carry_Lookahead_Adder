magic
tech scmos
timestamp 1171447631
<< checkpaint >>
rect -22 -26 118 114
<< ab >>
rect 0 0 96 88
<< pwell >>
rect -4 -8 100 40
<< nwell >>
rect -4 40 100 96
<< polysilicon >>
rect 2 82 11 83
rect 2 78 6 82
rect 10 78 11 82
rect 2 77 11 78
rect 9 74 11 77
rect 21 82 30 83
rect 21 78 25 82
rect 29 78 30 82
rect 21 77 30 78
rect 34 77 43 83
rect 21 74 23 77
rect 41 74 43 77
rect 53 77 62 83
rect 66 82 75 83
rect 66 78 67 82
rect 71 78 75 82
rect 66 77 75 78
rect 53 74 55 77
rect 73 74 75 77
rect 85 77 94 83
rect 85 74 87 77
rect 9 43 11 46
rect 21 43 23 46
rect 41 43 43 46
rect 53 43 55 46
rect 73 43 75 46
rect 85 43 87 46
rect 2 37 14 43
rect 18 42 30 43
rect 18 38 19 42
rect 23 38 30 42
rect 18 37 30 38
rect 34 42 46 43
rect 34 38 38 42
rect 42 38 46 42
rect 34 37 46 38
rect 50 37 62 43
rect 66 37 78 43
rect 82 42 94 43
rect 82 38 86 42
rect 90 38 94 42
rect 82 37 94 38
rect 9 34 11 37
rect 21 34 23 37
rect 41 34 43 37
rect 53 34 55 37
rect 73 34 75 37
rect 85 34 87 37
rect 9 11 11 14
rect 2 5 11 11
rect 21 11 23 14
rect 41 11 43 14
rect 21 5 30 11
rect 34 5 43 11
rect 53 11 55 14
rect 73 11 75 14
rect 53 10 62 11
rect 53 6 54 10
rect 58 6 62 10
rect 53 5 62 6
rect 66 5 75 11
rect 85 11 87 14
rect 85 5 94 11
<< ndiffusion >>
rect 2 14 9 34
rect 11 26 21 34
rect 11 22 14 26
rect 18 22 21 26
rect 11 19 21 22
rect 11 15 14 19
rect 18 15 21 19
rect 11 14 21 15
rect 23 33 30 34
rect 23 29 25 33
rect 29 29 30 33
rect 23 26 30 29
rect 23 22 25 26
rect 29 22 30 26
rect 23 14 30 22
rect 34 30 41 34
rect 34 26 35 30
rect 39 26 41 30
rect 34 23 41 26
rect 34 19 35 23
rect 39 19 41 23
rect 34 14 41 19
rect 43 33 53 34
rect 43 29 46 33
rect 50 29 53 33
rect 43 14 53 29
rect 55 30 62 34
rect 55 26 57 30
rect 61 26 62 30
rect 55 14 62 26
rect 66 22 73 34
rect 66 18 67 22
rect 71 18 73 22
rect 66 14 73 18
rect 75 22 85 34
rect 75 18 78 22
rect 82 18 85 22
rect 75 15 85 18
rect 75 14 78 15
rect 13 2 19 14
rect 45 2 51 14
rect 77 11 78 14
rect 82 14 85 15
rect 87 29 94 34
rect 87 25 89 29
rect 93 25 94 29
rect 87 22 94 25
rect 87 18 89 22
rect 93 18 94 22
rect 87 14 94 18
rect 82 11 83 14
rect 77 2 83 11
<< pdiffusion >>
rect 13 74 19 86
rect 45 74 51 86
rect 77 74 83 86
rect 2 46 9 74
rect 11 73 21 74
rect 11 69 14 73
rect 18 69 21 73
rect 11 66 21 69
rect 11 62 14 66
rect 18 62 21 66
rect 11 46 21 62
rect 23 58 30 74
rect 23 54 25 58
rect 29 54 30 58
rect 23 51 30 54
rect 23 47 25 51
rect 29 47 30 51
rect 23 46 30 47
rect 34 70 41 74
rect 34 66 35 70
rect 39 66 41 70
rect 34 46 41 66
rect 43 46 53 74
rect 55 70 62 74
rect 55 66 57 70
rect 61 66 62 70
rect 55 54 62 66
rect 55 50 57 54
rect 61 50 62 54
rect 55 46 62 50
rect 66 70 73 74
rect 66 66 67 70
rect 71 66 73 70
rect 66 54 73 66
rect 66 50 67 54
rect 71 50 73 54
rect 66 46 73 50
rect 75 59 85 74
rect 75 55 78 59
rect 82 55 85 59
rect 75 51 85 55
rect 75 47 78 51
rect 82 47 85 51
rect 75 46 85 47
rect 87 73 94 74
rect 87 69 89 73
rect 93 69 94 73
rect 87 66 94 69
rect 87 62 89 66
rect 93 62 94 66
rect 87 46 94 62
<< metal1 >>
rect -2 86 2 90
rect 10 86 22 90
rect 30 86 34 90
rect 42 86 54 90
rect 62 86 66 90
rect 74 86 86 90
rect 94 86 98 90
rect 6 82 10 86
rect 6 77 10 78
rect 14 82 18 86
rect 89 82 93 86
rect 24 78 25 82
rect 29 78 67 82
rect 71 78 72 82
rect 14 73 18 78
rect 89 73 93 78
rect 18 69 35 70
rect 14 66 35 69
rect 39 66 40 70
rect 56 66 57 70
rect 61 66 67 70
rect 71 66 72 70
rect 89 66 93 69
rect 14 61 18 62
rect 38 59 82 62
rect 89 61 93 62
rect 25 58 29 59
rect 14 42 18 55
rect 25 51 29 54
rect 38 58 78 59
rect 29 47 34 50
rect 25 46 34 47
rect 14 38 19 42
rect 23 38 24 42
rect 14 33 18 38
rect 30 34 34 46
rect 38 42 42 58
rect 38 37 42 38
rect 46 50 57 54
rect 61 50 67 54
rect 71 50 72 54
rect 78 51 82 55
rect 25 33 39 34
rect 29 30 39 33
rect 14 26 18 27
rect 14 19 18 22
rect 25 26 29 29
rect 25 21 29 22
rect 35 23 39 26
rect 46 33 50 50
rect 78 30 82 47
rect 86 42 90 55
rect 86 33 90 38
rect 46 25 50 29
rect 56 26 57 30
rect 61 29 93 30
rect 61 26 89 29
rect 78 22 82 23
rect 39 19 67 22
rect 35 18 67 19
rect 71 18 72 22
rect 14 10 18 15
rect 14 2 18 6
rect 54 10 58 18
rect 54 5 58 6
rect 78 15 82 18
rect 89 22 93 25
rect 89 17 93 18
rect 78 10 82 11
rect 78 2 82 6
rect -2 -2 2 2
rect 10 -2 22 2
rect 30 -2 34 2
rect 42 -2 54 2
rect 62 -2 66 2
rect 74 -2 86 2
rect 94 -2 98 2
<< metal2 >>
rect -2 86 6 90
rect 10 86 22 90
rect 26 86 38 90
rect 42 86 54 90
rect 58 86 70 90
rect 74 86 86 90
rect 90 86 98 90
rect -2 82 98 86
rect -2 78 14 82
rect 18 78 89 82
rect 93 78 98 82
rect -2 76 98 78
rect -2 10 98 12
rect -2 6 14 10
rect 18 6 78 10
rect 82 6 98 10
rect -2 2 98 6
rect -2 -2 6 2
rect 10 -2 22 2
rect 26 -2 38 2
rect 42 -2 54 2
rect 58 -2 70 2
rect 74 -2 86 2
rect 90 -2 98 2
<< ntransistor >>
rect 9 14 11 34
rect 21 14 23 34
rect 41 14 43 34
rect 53 14 55 34
rect 73 14 75 34
rect 85 14 87 34
<< ptransistor >>
rect 9 46 11 74
rect 21 46 23 74
rect 41 46 43 74
rect 53 46 55 74
rect 73 46 75 74
rect 85 46 87 74
<< polycontact >>
rect 6 78 10 82
rect 25 78 29 82
rect 67 78 71 82
rect 19 38 23 42
rect 38 38 42 42
rect 86 38 90 42
rect 54 6 58 10
<< ndcontact >>
rect 14 22 18 26
rect 14 15 18 19
rect 25 29 29 33
rect 25 22 29 26
rect 35 26 39 30
rect 35 19 39 23
rect 46 29 50 33
rect 57 26 61 30
rect 67 18 71 22
rect 78 18 82 22
rect 78 11 82 15
rect 89 25 93 29
rect 89 18 93 22
<< pdcontact >>
rect 14 69 18 73
rect 14 62 18 66
rect 25 54 29 58
rect 25 47 29 51
rect 35 66 39 70
rect 57 66 61 70
rect 57 50 61 54
rect 67 66 71 70
rect 67 50 71 54
rect 78 55 82 59
rect 78 47 82 51
rect 89 69 93 73
rect 89 62 93 66
<< m2contact >>
rect 6 86 10 90
rect 22 86 26 90
rect 38 86 42 90
rect 54 86 58 90
rect 70 86 74 90
rect 86 86 90 90
rect 14 78 18 82
rect 89 78 93 82
rect 14 6 18 10
rect 78 6 82 10
rect 6 -2 10 2
rect 22 -2 26 2
rect 38 -2 42 2
rect 54 -2 58 2
rect 70 -2 74 2
rect 86 -2 90 2
<< psubstratepcontact >>
rect 2 -2 6 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 90 -2 94 2
<< nsubstratencontact >>
rect 2 86 6 90
rect 26 86 30 90
rect 34 86 38 90
rect 58 86 62 90
rect 66 86 70 90
rect 90 86 94 90
<< psubstratepdiff >>
rect 0 2 7 3
rect 25 2 39 3
rect 57 2 71 3
rect 89 2 96 3
rect 0 -2 2 2
rect 6 -2 7 2
rect 0 -3 7 -2
rect 25 -2 26 2
rect 30 -2 34 2
rect 38 -2 39 2
rect 25 -3 39 -2
rect 57 -2 58 2
rect 62 -2 66 2
rect 70 -2 71 2
rect 57 -3 71 -2
rect 89 -2 90 2
rect 94 -2 96 2
rect 89 -3 96 -2
<< nsubstratendiff >>
rect 0 90 7 91
rect 0 86 2 90
rect 6 86 7 90
rect 25 90 39 91
rect 25 86 26 90
rect 30 86 34 90
rect 38 86 39 90
rect 57 90 71 91
rect 57 86 58 90
rect 62 86 66 90
rect 70 86 71 90
rect 89 90 96 91
rect 89 86 90 90
rect 94 86 96 90
rect 0 85 7 86
rect 25 85 39 86
rect 57 85 71 86
rect 89 85 96 86
<< labels >>
rlabel metal1 16 44 16 44 6 b
rlabel metal1 48 36 48 36 6 z
rlabel metal1 64 52 64 52 6 z
rlabel metal1 56 52 56 52 6 z
rlabel metal1 88 44 88 44 6 a
rlabel metal2 48 6 48 6 6 vss
rlabel metal2 48 82 48 82 6 vdd
<< end >>
