.subckt iv1v2x2 a vdd vss z
*   SPICE3 file   created from iv1v2x2.ext -      technology: scmos
m00 vdd    a      z      vdd p w=27u  l=2.3636u ad=216p     pd=70u      as=161p     ps=68u
m01 vss    a      z      vss n w=12u  l=2.3636u ad=96p      pd=40u      as=72p      ps=38u
C0  z      a      0.085f
C1  vss    z      0.022f
C2  vdd    a      0.025f
C3  vss    vdd    0.004f
C4  vdd    z      0.060f
C5  vss    a      0.025f
C8  z      vss    0.006f
C9  a      vss    0.023f
.ends
