magic
tech scmos
timestamp 1170759820
<< checkpaint >>
rect -22 -26 86 114
<< ab >>
rect 0 0 64 88
<< pwell >>
rect -4 -8 68 40
<< nwell >>
rect -4 40 68 96
<< polysilicon >>
rect 2 77 11 83
rect 9 74 11 77
rect 21 77 30 83
rect 34 82 43 83
rect 34 78 38 82
rect 42 78 43 82
rect 34 77 43 78
rect 21 74 23 77
rect 41 74 43 77
rect 53 82 62 83
rect 53 78 54 82
rect 58 78 62 82
rect 53 77 62 78
rect 53 74 55 77
rect 9 43 11 46
rect 21 43 23 46
rect 41 43 43 46
rect 53 43 55 46
rect 2 42 14 43
rect 2 38 6 42
rect 10 38 14 42
rect 2 37 14 38
rect 18 42 30 43
rect 18 38 22 42
rect 26 38 30 42
rect 18 37 30 38
rect 34 37 46 43
rect 50 42 62 43
rect 50 38 54 42
rect 58 38 62 42
rect 50 37 62 38
rect 9 34 11 37
rect 21 34 23 37
rect 41 34 43 37
rect 53 34 55 37
rect 9 11 11 14
rect 2 5 11 11
rect 21 11 23 14
rect 41 11 43 14
rect 21 5 30 11
rect 34 5 43 11
rect 53 11 55 14
rect 53 5 62 11
<< ndiffusion >>
rect 2 26 9 34
rect 2 22 3 26
rect 7 22 9 26
rect 2 19 9 22
rect 2 15 3 19
rect 7 15 9 19
rect 2 14 9 15
rect 11 29 21 34
rect 11 25 14 29
rect 18 25 21 29
rect 11 22 21 25
rect 11 18 14 22
rect 18 18 21 22
rect 11 14 21 18
rect 23 19 30 34
rect 23 15 25 19
rect 29 15 30 19
rect 23 14 30 15
rect 34 19 41 34
rect 34 15 35 19
rect 39 15 41 19
rect 34 14 41 15
rect 43 29 53 34
rect 43 25 46 29
rect 50 25 53 29
rect 43 22 53 25
rect 43 18 46 22
rect 50 18 53 22
rect 43 14 53 18
rect 55 19 62 34
rect 55 15 57 19
rect 61 15 62 19
rect 55 14 62 15
rect 13 2 19 14
rect 45 2 51 14
<< pdiffusion >>
rect 13 74 19 86
rect 45 74 51 86
rect 2 73 9 74
rect 2 69 3 73
rect 7 69 9 73
rect 2 66 9 69
rect 2 62 3 66
rect 7 62 9 66
rect 2 46 9 62
rect 11 66 21 74
rect 11 62 14 66
rect 18 62 21 66
rect 11 59 21 62
rect 11 55 14 59
rect 18 55 21 59
rect 11 46 21 55
rect 23 73 30 74
rect 23 69 25 73
rect 29 69 30 73
rect 23 66 30 69
rect 23 62 25 66
rect 29 62 30 66
rect 23 46 30 62
rect 34 66 41 74
rect 34 62 35 66
rect 39 62 41 66
rect 34 59 41 62
rect 34 55 35 59
rect 39 55 41 59
rect 34 46 41 55
rect 43 58 53 74
rect 43 54 46 58
rect 50 54 53 58
rect 43 51 53 54
rect 43 47 46 51
rect 50 47 53 51
rect 43 46 53 47
rect 55 66 62 74
rect 55 62 57 66
rect 61 62 62 66
rect 55 59 62 62
rect 55 55 57 59
rect 61 55 62 59
rect 55 46 62 55
<< metal1 >>
rect -2 86 2 90
rect 10 86 22 90
rect 30 86 34 90
rect 42 86 54 90
rect 62 86 66 90
rect 3 82 7 86
rect 3 73 7 78
rect 3 66 7 69
rect 25 82 29 86
rect 37 78 38 82
rect 42 78 54 82
rect 58 78 59 82
rect 25 73 29 78
rect 3 61 7 62
rect 14 66 18 67
rect 14 59 18 62
rect 25 66 29 69
rect 25 61 29 62
rect 35 66 61 67
rect 39 63 57 66
rect 35 59 39 62
rect 57 59 61 62
rect 18 55 35 58
rect 6 42 10 55
rect 14 54 39 55
rect 46 58 50 59
rect 57 54 61 55
rect 46 51 50 54
rect 21 42 27 46
rect 21 38 22 42
rect 26 38 27 42
rect 6 34 27 38
rect 6 33 10 34
rect 46 30 50 47
rect 14 29 50 30
rect 3 26 7 27
rect 3 19 7 22
rect 18 26 46 29
rect 14 22 18 25
rect 54 42 58 47
rect 54 25 58 38
rect 46 22 50 25
rect 14 17 18 18
rect 25 19 29 20
rect 3 10 7 15
rect 3 2 7 6
rect 25 10 29 15
rect 25 2 29 6
rect 35 19 39 20
rect 46 17 50 18
rect 57 19 61 20
rect 35 10 39 15
rect 35 2 39 6
rect 57 10 61 15
rect 57 2 61 6
rect -2 -2 2 2
rect 10 -2 22 2
rect 30 -2 34 2
rect 42 -2 54 2
rect 62 -2 66 2
<< metal2 >>
rect -2 86 6 90
rect 10 86 22 90
rect 26 86 38 90
rect 42 86 54 90
rect 58 86 66 90
rect -2 82 66 86
rect -2 78 3 82
rect 7 78 25 82
rect 29 78 66 82
rect -2 76 66 78
rect -2 10 66 12
rect -2 6 3 10
rect 7 6 25 10
rect 29 6 35 10
rect 39 6 57 10
rect 61 6 66 10
rect -2 2 66 6
rect -2 -2 6 2
rect 10 -2 22 2
rect 26 -2 38 2
rect 42 -2 54 2
rect 58 -2 66 2
<< ntransistor >>
rect 9 14 11 34
rect 21 14 23 34
rect 41 14 43 34
rect 53 14 55 34
<< ptransistor >>
rect 9 46 11 74
rect 21 46 23 74
rect 41 46 43 74
rect 53 46 55 74
<< polycontact >>
rect 38 78 42 82
rect 54 78 58 82
rect 6 38 10 42
rect 22 38 26 42
rect 54 38 58 42
<< ndcontact >>
rect 3 22 7 26
rect 3 15 7 19
rect 14 25 18 29
rect 14 18 18 22
rect 25 15 29 19
rect 35 15 39 19
rect 46 25 50 29
rect 46 18 50 22
rect 57 15 61 19
<< pdcontact >>
rect 3 69 7 73
rect 3 62 7 66
rect 14 62 18 66
rect 14 55 18 59
rect 25 69 29 73
rect 25 62 29 66
rect 35 62 39 66
rect 35 55 39 59
rect 46 54 50 58
rect 46 47 50 51
rect 57 62 61 66
rect 57 55 61 59
<< m2contact >>
rect 6 86 10 90
rect 22 86 26 90
rect 38 86 42 90
rect 54 86 58 90
rect 3 78 7 82
rect 25 78 29 82
rect 3 6 7 10
rect 25 6 29 10
rect 35 6 39 10
rect 57 6 61 10
rect 6 -2 10 2
rect 22 -2 26 2
rect 38 -2 42 2
rect 54 -2 58 2
<< psubstratepcontact >>
rect 2 -2 6 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 58 -2 62 2
<< nsubstratencontact >>
rect 2 86 6 90
rect 26 86 30 90
rect 34 86 38 90
rect 58 86 62 90
<< psubstratepdiff >>
rect 0 2 7 3
rect 25 2 39 3
rect 57 2 64 3
rect 0 -2 2 2
rect 6 -2 7 2
rect 0 -3 7 -2
rect 25 -2 26 2
rect 30 -2 34 2
rect 38 -2 39 2
rect 25 -3 39 -2
rect 57 -2 58 2
rect 62 -2 64 2
rect 57 -3 64 -2
<< nsubstratendiff >>
rect 0 90 7 91
rect 0 86 2 90
rect 6 86 7 90
rect 25 90 39 91
rect 25 86 26 90
rect 30 86 34 90
rect 38 86 39 90
rect 57 90 64 91
rect 57 86 58 90
rect 62 86 64 90
rect 0 85 7 86
rect 25 85 39 86
rect 57 85 64 86
<< labels >>
rlabel metal1 8 44 8 44 6 a
rlabel ndcontact 16 20 16 20 6 z
rlabel metal1 16 36 16 36 6 a
rlabel metal1 24 28 24 28 6 z
rlabel metal1 32 28 32 28 6 z
rlabel polycontact 24 40 24 40 6 a
rlabel metal1 40 28 40 28 6 z
rlabel metal1 48 36 48 36 6 z
rlabel metal1 56 36 56 36 6 b
rlabel metal2 32 6 32 6 6 vss
rlabel metal2 32 82 32 82 6 vdd
<< end >>
