magic
tech scmos
timestamp 1179385040
<< checkpaint >>
rect -22 -22 78 94
<< ab >>
rect 0 0 56 72
<< pwell >>
rect -4 -4 60 32
<< nwell >>
rect -4 32 60 76
<< polysilicon >>
rect 9 66 11 70
rect 19 66 21 70
rect 29 57 31 62
rect 39 57 41 61
rect 9 35 11 38
rect 19 35 21 38
rect 29 35 31 42
rect 39 39 41 42
rect 39 38 47 39
rect 9 34 22 35
rect 9 30 17 34
rect 21 30 22 34
rect 9 29 22 30
rect 28 34 34 35
rect 28 30 29 34
rect 33 30 34 34
rect 28 29 34 30
rect 10 26 12 29
rect 20 26 22 29
rect 32 26 34 29
rect 39 34 42 38
rect 46 34 47 38
rect 39 33 47 34
rect 39 26 41 33
rect 10 7 12 12
rect 20 7 22 12
rect 32 9 34 14
rect 39 9 41 14
<< ndiffusion >>
rect 2 12 10 26
rect 12 18 20 26
rect 12 14 14 18
rect 18 14 20 18
rect 12 12 20 14
rect 22 14 32 26
rect 34 14 39 26
rect 41 20 46 26
rect 41 19 48 20
rect 41 15 43 19
rect 47 15 48 19
rect 41 14 48 15
rect 22 12 30 14
rect 2 8 8 12
rect 2 4 3 8
rect 7 4 8 8
rect 24 8 30 12
rect 2 3 8 4
rect 24 4 25 8
rect 29 4 30 8
rect 24 3 30 4
<< pdiffusion >>
rect 2 65 9 66
rect 2 61 3 65
rect 7 61 9 65
rect 2 58 9 61
rect 2 54 3 58
rect 7 54 9 58
rect 2 38 9 54
rect 11 58 19 66
rect 11 54 13 58
rect 17 54 19 58
rect 11 51 19 54
rect 11 47 13 51
rect 17 47 19 51
rect 11 38 19 47
rect 21 57 27 66
rect 21 56 29 57
rect 21 52 23 56
rect 27 52 29 56
rect 21 42 29 52
rect 31 56 39 57
rect 31 52 33 56
rect 37 52 39 56
rect 31 49 39 52
rect 31 45 33 49
rect 37 45 39 49
rect 31 42 39 45
rect 41 56 48 57
rect 41 52 43 56
rect 47 52 48 56
rect 41 49 48 52
rect 41 45 43 49
rect 47 45 48 49
rect 41 42 48 45
rect 21 38 27 42
<< metal1 >>
rect -2 68 58 72
rect -2 65 34 68
rect -2 64 3 65
rect 2 61 3 64
rect 7 64 34 65
rect 38 64 42 68
rect 46 64 58 68
rect 7 61 8 64
rect 2 58 8 61
rect 2 54 3 58
rect 7 54 8 58
rect 13 58 17 59
rect 13 51 17 54
rect 22 56 28 64
rect 42 56 48 64
rect 22 52 23 56
rect 27 52 28 56
rect 32 52 33 56
rect 37 52 38 56
rect 2 47 13 50
rect 32 49 38 52
rect 2 46 17 47
rect 2 18 6 46
rect 23 45 33 49
rect 37 45 38 49
rect 42 52 43 56
rect 47 52 48 56
rect 42 49 48 52
rect 42 45 43 49
rect 47 45 48 49
rect 23 42 27 45
rect 17 38 27 42
rect 33 38 46 42
rect 17 34 21 38
rect 25 30 29 34
rect 33 30 38 34
rect 17 26 21 30
rect 17 22 28 26
rect 2 14 14 18
rect 18 14 19 18
rect 2 13 19 14
rect 24 17 28 22
rect 34 21 38 30
rect 42 29 46 34
rect 43 19 47 20
rect 24 15 43 17
rect 24 13 47 15
rect -2 4 3 8
rect 7 4 25 8
rect 29 4 48 8
rect 52 4 58 8
rect -2 0 58 4
<< ntransistor >>
rect 10 12 12 26
rect 20 12 22 26
rect 32 14 34 26
rect 39 14 41 26
<< ptransistor >>
rect 9 38 11 66
rect 19 38 21 66
rect 29 42 31 57
rect 39 42 41 57
<< polycontact >>
rect 17 30 21 34
rect 29 30 33 34
rect 42 34 46 38
<< ndcontact >>
rect 14 14 18 18
rect 43 15 47 19
rect 3 4 7 8
rect 25 4 29 8
<< pdcontact >>
rect 3 61 7 65
rect 3 54 7 58
rect 13 54 17 58
rect 13 47 17 51
rect 23 52 27 56
rect 33 52 37 56
rect 33 45 37 49
rect 43 52 47 56
rect 43 45 47 49
<< psubstratepcontact >>
rect 48 4 52 8
<< nsubstratencontact >>
rect 34 64 38 68
rect 42 64 46 68
<< psubstratepdiff >>
rect 47 8 53 9
rect 47 4 48 8
rect 52 4 53 8
rect 47 3 53 4
<< nsubstratendiff >>
rect 33 68 47 69
rect 33 64 34 68
rect 38 64 42 68
rect 46 64 47 68
rect 33 63 47 64
<< labels >>
rlabel polysilicon 15 32 15 32 6 zn
rlabel metal1 4 28 4 28 6 z
rlabel metal1 12 16 12 16 6 z
rlabel polycontact 19 32 19 32 6 zn
rlabel metal1 12 48 12 48 6 z
rlabel metal1 28 4 28 4 6 vss
rlabel metal1 28 32 28 32 6 a
rlabel metal1 36 24 36 24 6 a
rlabel metal1 36 40 36 40 6 b
rlabel metal1 30 47 30 47 6 zn
rlabel metal1 35 50 35 50 6 zn
rlabel metal1 28 68 28 68 6 vdd
rlabel ndcontact 45 16 45 16 6 zn
rlabel metal1 44 32 44 32 6 b
<< end >>
