.subckt nr3_x1 a b c vdd vss z
*   SPICE3 file   created from nr3_x1.ext -      technology: scmos
m00 w1     a      vdd    vdd p w=39u  l=2.3636u ad=117p     pd=45u      as=331.5p   ps=95u
m01 w2     b      w1     vdd p w=39u  l=2.3636u ad=117p     pd=45u      as=117p     ps=45u
m02 z      c      w2     vdd p w=39u  l=2.3636u ad=195p     pd=49u      as=117p     ps=45u
m03 w3     c      z      vdd p w=39u  l=2.3636u ad=117p     pd=45u      as=195p     ps=49u
m04 w4     b      w3     vdd p w=39u  l=2.3636u ad=117p     pd=45u      as=117p     ps=45u
m05 vdd    a      w4     vdd p w=39u  l=2.3636u ad=331.5p   pd=95u      as=117p     ps=45u
m06 vss    a      z      vss n w=15u  l=2.3636u ad=95p      pd=32.6667u as=81p      ps=32u
m07 z      b      vss    vss n w=15u  l=2.3636u ad=81p      pd=32u      as=95p      ps=32.6667u
m08 vss    c      z      vss n w=15u  l=2.3636u ad=95p      pd=32.6667u as=81p      ps=32u
C0  z      vdd    0.159f
C1  vss    a      0.024f
C2  z      b      0.113f
C3  w3     a      0.012f
C4  w1     vdd    0.011f
C5  w2     a      0.012f
C6  vdd    c      0.010f
C7  vdd    a      0.076f
C8  c      b      0.246f
C9  b      a      0.510f
C10 z      w1     0.013f
C11 vss    b      0.032f
C12 w3     vdd    0.011f
C13 w2     vdd    0.011f
C14 w4     a      0.013f
C15 z      c      0.027f
C16 z      a      0.394f
C17 vss    z      0.247f
C18 vdd    b      0.031f
C19 w1     a      0.012f
C20 c      a      0.146f
C21 w4     vdd    0.011f
C22 vss    c      0.099f
C23 z      w2     0.013f
C25 z      vss    0.017f
C27 c      vss    0.054f
C28 b      vss    0.049f
C29 a      vss    0.047f
.ends
