.subckt nd4_x2 a b c d vdd vss z
*   SPICE3 file   created from nd4_x2.ext -      technology: scmos
m00 z      a      vdd    vdd p w=39u  l=2.3636u ad=195p     pd=49u      as=273p     ps=72.5u
m01 vdd    b      z      vdd p w=39u  l=2.3636u ad=273p     pd=72.5u    as=195p     ps=49u
m02 z      c      vdd    vdd p w=39u  l=2.3636u ad=195p     pd=49u      as=273p     ps=72.5u
m03 vdd    d      z      vdd p w=39u  l=2.3636u ad=273p     pd=72.5u    as=195p     ps=49u
m04 w1     a      vss    vss n w=23u  l=2.3636u ad=69p      pd=29u      as=195.5p   ps=63u
m05 w2     b      w1     vss n w=23u  l=2.3636u ad=69p      pd=29u      as=69p      ps=29u
m06 w3     c      w2     vss n w=23u  l=2.3636u ad=69p      pd=29u      as=69p      ps=29u
m07 z      d      w3     vss n w=23u  l=2.3636u ad=115p     pd=33u      as=69p      ps=29u
m08 w4     d      z      vss n w=23u  l=2.3636u ad=69p      pd=29u      as=115p     ps=33u
m09 w5     c      w4     vss n w=23u  l=2.3636u ad=69p      pd=29u      as=69p      ps=29u
m10 w6     b      w5     vss n w=23u  l=2.3636u ad=69p      pd=29u      as=69p      ps=29u
m11 vss    a      w6     vss n w=23u  l=2.3636u ad=195.5p   pd=63u      as=69p      ps=29u
C0  vss    z      0.324f
C1  w5     a      0.006f
C2  vss    d      0.032f
C3  z      vdd    0.358f
C4  w3     a      0.006f
C5  w6     vss    0.010f
C6  vdd    d      0.029f
C7  vss    b      0.015f
C8  w1     a      0.006f
C9  z      c      0.104f
C10 w4     vss    0.010f
C11 vdd    b      0.174f
C12 z      a      0.394f
C13 d      c      0.377f
C14 w3     z      0.013f
C15 w2     vss    0.010f
C16 d      a      0.154f
C17 c      b      0.344f
C18 w6     a      0.006f
C19 w1     z      0.013f
C20 b      a      0.235f
C21 w4     a      0.006f
C22 z      d      0.022f
C23 vss    c      0.042f
C24 w2     a      0.006f
C25 w5     vss    0.010f
C26 vss    a      0.145f
C27 z      b      0.278f
C28 vdd    c      0.021f
C29 w3     vss    0.010f
C30 vdd    a      0.009f
C31 d      b      0.178f
C32 w2     z      0.013f
C33 w1     vss    0.010f
C34 c      a      0.291f
C36 z      vss    0.012f
C38 d      vss    0.045f
C39 c      vss    0.051f
C40 b      vss    0.051f
C41 a      vss    0.055f
.ends
