magic
tech scmos
timestamp 1179387776
<< checkpaint >>
rect -22 -22 94 94
<< ab >>
rect 0 0 72 72
<< pwell >>
rect -4 -4 76 32
<< nwell >>
rect -4 32 76 76
<< polysilicon >>
rect 32 68 63 70
rect 9 56 11 61
rect 19 59 25 60
rect 19 55 20 59
rect 24 55 25 59
rect 32 56 34 68
rect 61 63 63 68
rect 19 54 25 55
rect 29 54 34 56
rect 39 59 45 60
rect 39 55 40 59
rect 44 55 45 59
rect 39 54 45 55
rect 19 51 21 54
rect 29 51 31 54
rect 39 51 41 54
rect 49 51 51 56
rect 9 35 11 38
rect 19 36 21 39
rect 9 34 15 35
rect 9 30 10 34
rect 14 30 15 34
rect 19 33 23 36
rect 29 35 31 39
rect 39 36 41 39
rect 49 36 51 39
rect 9 29 15 30
rect 9 26 11 29
rect 21 26 23 33
rect 35 34 41 36
rect 48 35 54 36
rect 61 35 63 51
rect 35 31 37 34
rect 31 29 37 31
rect 48 31 49 35
rect 53 31 54 35
rect 48 30 54 31
rect 58 34 64 35
rect 58 30 59 34
rect 63 30 64 34
rect 31 26 33 29
rect 41 26 43 30
rect 51 26 53 30
rect 58 29 64 30
rect 61 26 63 29
rect 9 12 11 17
rect 21 15 23 20
rect 31 15 33 20
rect 41 4 43 20
rect 51 15 53 20
rect 61 4 63 20
rect 41 2 63 4
<< ndiffusion >>
rect 2 25 9 26
rect 2 21 3 25
rect 7 21 9 25
rect 2 20 9 21
rect 4 17 9 20
rect 11 20 21 26
rect 23 25 31 26
rect 23 21 25 25
rect 29 21 31 25
rect 23 20 31 21
rect 33 25 41 26
rect 33 21 35 25
rect 39 21 41 25
rect 33 20 41 21
rect 43 25 51 26
rect 43 21 45 25
rect 49 21 51 25
rect 43 20 51 21
rect 53 20 61 26
rect 63 25 70 26
rect 63 21 65 25
rect 69 21 70 25
rect 63 20 70 21
rect 11 17 19 20
rect 13 8 19 17
rect 13 4 14 8
rect 18 4 19 8
rect 13 3 19 4
rect 55 13 59 20
rect 53 11 59 13
rect 53 7 54 11
rect 58 7 59 11
rect 53 6 59 7
<< pdiffusion >>
rect 13 68 19 69
rect 13 64 14 68
rect 18 64 19 68
rect 13 62 19 64
rect 13 56 17 62
rect 4 44 9 56
rect 2 43 9 44
rect 2 39 3 43
rect 7 39 9 43
rect 2 38 9 39
rect 11 51 17 56
rect 53 65 59 66
rect 53 61 54 65
rect 58 63 59 65
rect 58 61 61 63
rect 53 51 61 61
rect 63 59 68 63
rect 63 58 70 59
rect 63 54 65 58
rect 69 54 70 58
rect 63 53 70 54
rect 63 51 68 53
rect 11 39 19 51
rect 21 44 29 51
rect 21 40 23 44
rect 27 40 29 44
rect 21 39 29 40
rect 31 44 39 51
rect 31 40 33 44
rect 37 40 39 44
rect 31 39 39 40
rect 41 44 49 51
rect 41 40 43 44
rect 47 40 49 44
rect 41 39 49 40
rect 51 39 59 51
rect 11 38 17 39
<< metal1 >>
rect -2 68 74 72
rect -2 64 4 68
rect 8 64 14 68
rect 18 64 24 68
rect 28 65 74 68
rect 28 64 54 65
rect 53 61 54 64
rect 58 64 74 65
rect 58 61 59 64
rect 9 55 20 59
rect 24 55 25 59
rect 9 54 25 55
rect 39 55 40 59
rect 44 58 45 59
rect 44 55 65 58
rect 39 54 65 55
rect 69 54 70 58
rect 9 46 15 54
rect 25 47 55 51
rect 25 45 29 47
rect 23 44 29 45
rect 2 39 3 43
rect 7 42 8 43
rect 7 39 15 42
rect 27 40 29 44
rect 32 40 33 44
rect 37 40 38 44
rect 23 39 29 40
rect 2 38 15 39
rect 2 26 6 38
rect 9 30 10 34
rect 14 30 19 34
rect 2 25 7 26
rect 2 21 3 25
rect 2 20 7 21
rect 15 17 19 30
rect 25 25 29 39
rect 25 20 29 21
rect 34 26 38 40
rect 42 40 43 44
rect 47 40 48 44
rect 34 25 39 26
rect 34 21 35 25
rect 42 25 46 40
rect 51 36 55 47
rect 49 35 55 36
rect 53 31 55 35
rect 49 30 55 31
rect 58 34 63 35
rect 58 30 59 34
rect 58 29 63 30
rect 42 21 45 25
rect 49 21 50 25
rect 34 20 39 21
rect 34 17 38 20
rect 58 18 62 29
rect 66 26 70 54
rect 65 25 70 26
rect 69 21 70 25
rect 65 20 70 21
rect 15 13 38 17
rect 49 14 62 18
rect 53 8 54 11
rect -2 4 4 8
rect 8 4 14 8
rect 18 4 33 8
rect 37 7 54 8
rect 58 8 59 11
rect 58 7 74 8
rect 37 4 74 7
rect -2 0 74 4
<< ntransistor >>
rect 9 17 11 26
rect 21 20 23 26
rect 31 20 33 26
rect 41 20 43 26
rect 51 20 53 26
rect 61 20 63 26
<< ptransistor >>
rect 9 38 11 56
rect 61 51 63 63
rect 19 39 21 51
rect 29 39 31 51
rect 39 39 41 51
rect 49 39 51 51
<< polycontact >>
rect 20 55 24 59
rect 40 55 44 59
rect 10 30 14 34
rect 49 31 53 35
rect 59 30 63 34
<< ndcontact >>
rect 3 21 7 25
rect 25 21 29 25
rect 35 21 39 25
rect 45 21 49 25
rect 65 21 69 25
rect 14 4 18 8
rect 54 7 58 11
<< pdcontact >>
rect 14 64 18 68
rect 3 39 7 43
rect 54 61 58 65
rect 65 54 69 58
rect 23 40 27 44
rect 33 40 37 44
rect 43 40 47 44
<< psubstratepcontact >>
rect 4 4 8 8
rect 33 4 37 8
<< nsubstratencontact >>
rect 4 64 8 68
rect 24 64 28 68
<< psubstratepdiff >>
rect 3 8 9 9
rect 3 4 4 8
rect 8 4 9 8
rect 3 3 9 4
rect 32 8 38 9
rect 32 4 33 8
rect 37 4 38 8
rect 32 3 38 4
<< nsubstratendiff >>
rect 3 68 9 69
rect 3 64 4 68
rect 8 64 9 68
rect 3 63 9 64
rect 23 68 29 69
rect 23 64 24 68
rect 28 64 29 68
rect 23 63 29 64
<< labels >>
rlabel polycontact 12 32 12 32 6 zn
rlabel polycontact 42 57 42 57 6 bn
rlabel polycontact 51 33 51 33 6 an
rlabel metal1 4 28 4 28 6 z
rlabel metal1 12 40 12 40 6 z
rlabel metal1 12 52 12 52 6 a
rlabel metal1 14 32 14 32 6 zn
rlabel metal1 27 35 27 35 6 an
rlabel metal1 20 56 20 56 6 a
rlabel metal1 36 4 36 4 6 vss
rlabel metal1 52 16 52 16 6 b
rlabel metal1 53 40 53 40 6 an
rlabel metal1 44 32 44 32 6 ai
rlabel metal1 36 28 36 28 6 zn
rlabel metal1 36 68 36 68 6 vdd
rlabel metal1 60 28 60 28 6 b
rlabel metal1 54 56 54 56 6 bn
rlabel metal1 68 39 68 39 6 bn
<< end >>
