magic
tech scmos
timestamp 1179385262
<< checkpaint >>
rect -22 -25 62 105
<< ab >>
rect 0 0 40 80
<< pwell >>
rect -4 -7 44 36
<< nwell >>
rect -4 36 44 87
<< polysilicon >>
rect 29 66 31 71
rect 9 58 11 63
rect 19 58 21 63
rect 29 47 31 50
rect 29 46 35 47
rect 29 42 30 46
rect 34 42 35 46
rect 9 39 11 42
rect 9 38 15 39
rect 9 34 10 38
rect 14 34 15 38
rect 9 33 15 34
rect 19 35 21 42
rect 29 41 35 42
rect 19 34 25 35
rect 12 25 14 33
rect 19 30 20 34
rect 24 30 25 34
rect 19 29 25 30
rect 22 26 24 29
rect 29 26 31 41
rect 12 15 14 19
rect 22 15 24 19
rect 29 15 31 19
<< ndiffusion >>
rect 17 25 22 26
rect 3 19 12 25
rect 14 24 22 25
rect 14 20 16 24
rect 20 20 22 24
rect 14 19 22 20
rect 24 19 29 26
rect 31 19 38 26
rect 3 12 10 19
rect 33 13 38 19
rect 3 8 5 12
rect 9 8 10 12
rect 3 7 10 8
rect 32 12 38 13
rect 32 8 33 12
rect 37 8 38 12
rect 32 7 38 8
<< pdiffusion >>
rect 21 72 27 73
rect 21 68 22 72
rect 26 68 27 72
rect 21 66 27 68
rect 21 65 29 66
rect 23 58 29 65
rect 4 55 9 58
rect 2 54 9 55
rect 2 50 3 54
rect 7 50 9 54
rect 2 47 9 50
rect 2 43 3 47
rect 7 43 9 47
rect 2 42 9 43
rect 11 57 19 58
rect 11 53 13 57
rect 17 53 19 57
rect 11 42 19 53
rect 21 50 29 58
rect 31 63 36 66
rect 31 62 38 63
rect 31 58 33 62
rect 37 58 38 62
rect 31 55 38 58
rect 31 51 33 55
rect 37 51 38 55
rect 31 50 38 51
rect 21 42 27 50
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect -2 72 42 78
rect -2 68 22 72
rect 26 68 42 72
rect 13 62 37 63
rect 13 59 33 62
rect 13 57 17 59
rect 2 54 7 55
rect 2 50 3 54
rect 33 55 37 58
rect 13 52 17 53
rect 2 47 7 50
rect 26 47 30 55
rect 33 50 37 51
rect 2 43 3 47
rect 2 42 7 43
rect 2 23 6 42
rect 10 41 22 47
rect 26 46 38 47
rect 26 42 30 46
rect 34 42 38 46
rect 26 41 38 42
rect 10 38 14 41
rect 10 33 14 34
rect 19 30 20 34
rect 24 33 25 34
rect 24 30 30 33
rect 19 29 30 30
rect 16 24 20 25
rect 2 20 16 23
rect 26 23 30 29
rect 20 20 22 23
rect 2 17 22 20
rect 26 17 38 23
rect -2 8 5 12
rect 9 8 33 12
rect 37 8 42 12
rect -2 2 42 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
<< ntransistor >>
rect 12 19 14 25
rect 22 19 24 26
rect 29 19 31 26
<< ptransistor >>
rect 9 42 11 58
rect 19 42 21 58
rect 29 50 31 66
<< polycontact >>
rect 30 42 34 46
rect 10 34 14 38
rect 20 30 24 34
<< ndcontact >>
rect 16 20 20 24
rect 5 8 9 12
rect 33 8 37 12
<< pdcontact >>
rect 22 68 26 72
rect 3 50 7 54
rect 3 43 7 47
rect 13 53 17 57
rect 33 58 37 62
rect 33 51 37 55
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
<< psubstratepdiff >>
rect 0 2 40 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 40 2
rect 0 -3 40 -2
<< nsubstratendiff >>
rect 0 82 40 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 40 82
rect 0 77 40 78
<< labels >>
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 20 12 20 6 z
rlabel metal1 12 40 12 40 6 b
rlabel metal1 15 57 15 57 6 n1
rlabel metal1 20 6 20 6 6 vss
rlabel metal1 20 20 20 20 6 z
rlabel metal1 28 24 28 24 6 a2
rlabel metal1 20 44 20 44 6 b
rlabel metal1 28 48 28 48 6 a1
rlabel metal1 20 74 20 74 6 vdd
rlabel metal1 36 20 36 20 6 a2
rlabel metal1 36 44 36 44 6 a1
rlabel metal1 35 56 35 56 6 n1
<< end >>
