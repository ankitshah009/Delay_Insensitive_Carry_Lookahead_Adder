magic
tech scmos
timestamp 1179386540
<< checkpaint >>
rect -22 -25 62 105
<< ab >>
rect 0 0 40 80
<< pwell >>
rect -4 -7 44 36
<< nwell >>
rect -4 36 44 87
<< polysilicon >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 9 39 11 50
rect 19 47 21 50
rect 19 46 25 47
rect 19 42 20 46
rect 24 42 25 46
rect 19 41 25 42
rect 9 38 15 39
rect 9 34 10 38
rect 14 34 15 38
rect 9 33 15 34
rect 12 30 14 33
rect 19 30 21 41
rect 29 39 31 50
rect 29 38 35 39
rect 29 35 30 38
rect 26 34 30 35
rect 34 34 35 38
rect 26 33 35 34
rect 26 30 28 33
rect 12 6 14 10
rect 19 6 21 10
rect 26 6 28 10
<< ndiffusion >>
rect 7 22 12 30
rect 5 21 12 22
rect 5 17 6 21
rect 10 17 12 21
rect 5 16 12 17
rect 7 10 12 16
rect 14 10 19 30
rect 21 10 26 30
rect 28 14 36 30
rect 28 10 31 14
rect 35 10 36 14
rect 30 8 36 10
<< pdiffusion >>
rect 4 63 9 70
rect 2 62 9 63
rect 2 58 3 62
rect 7 58 9 62
rect 2 55 9 58
rect 2 51 3 55
rect 7 51 9 55
rect 2 50 9 51
rect 11 69 19 70
rect 11 65 13 69
rect 17 65 19 69
rect 11 62 19 65
rect 11 58 13 62
rect 17 58 19 62
rect 11 50 19 58
rect 21 62 29 70
rect 21 58 23 62
rect 27 58 29 62
rect 21 55 29 58
rect 21 51 23 55
rect 27 51 29 55
rect 21 50 29 51
rect 31 69 38 70
rect 31 65 33 69
rect 37 65 38 69
rect 31 62 38 65
rect 31 58 33 62
rect 37 58 38 62
rect 31 50 38 58
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect -2 69 42 78
rect -2 68 13 69
rect 12 65 13 68
rect 17 68 33 69
rect 17 65 18 68
rect 2 62 7 63
rect 2 58 3 62
rect 12 62 18 65
rect 32 65 33 68
rect 37 68 42 69
rect 37 65 38 68
rect 12 58 13 62
rect 17 58 18 62
rect 23 62 27 63
rect 32 62 38 65
rect 32 58 33 62
rect 37 58 38 62
rect 2 55 7 58
rect 2 51 3 55
rect 23 55 27 58
rect 7 51 23 54
rect 2 50 27 51
rect 2 17 6 50
rect 34 46 38 55
rect 19 42 20 46
rect 24 42 38 46
rect 10 38 14 39
rect 25 34 30 38
rect 10 30 14 34
rect 10 25 23 30
rect 10 17 11 21
rect 34 17 38 38
rect 30 12 31 14
rect -2 10 31 12
rect 35 12 36 14
rect 35 10 42 12
rect -2 2 42 10
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
<< ntransistor >>
rect 12 10 14 30
rect 19 10 21 30
rect 26 10 28 30
<< ptransistor >>
rect 9 50 11 70
rect 19 50 21 70
rect 29 50 31 70
<< polycontact >>
rect 20 42 24 46
rect 10 34 14 38
rect 30 34 34 38
<< ndcontact >>
rect 6 17 10 21
rect 31 10 35 14
<< pdcontact >>
rect 3 58 7 62
rect 3 51 7 55
rect 13 65 17 69
rect 13 58 17 62
rect 23 58 27 62
rect 23 51 27 55
rect 33 65 37 69
rect 33 58 37 62
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
<< psubstratepdiff >>
rect 0 2 40 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 40 2
rect 0 -3 40 -2
<< nsubstratendiff >>
rect 0 82 40 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 40 82
rect 0 77 40 78
<< labels >>
rlabel metal1 4 40 4 40 6 z
rlabel metal1 12 32 12 32 6 c
rlabel metal1 12 52 12 52 6 z
rlabel metal1 20 6 20 6 6 vss
rlabel metal1 20 28 20 28 6 c
rlabel metal1 28 36 28 36 6 a
rlabel metal1 28 44 28 44 6 b
rlabel metal1 20 52 20 52 6 z
rlabel metal1 20 74 20 74 6 vdd
rlabel metal1 36 24 36 24 6 a
rlabel metal1 36 52 36 52 6 b
<< end >>
