magic
tech scmos
timestamp 1179387280
<< checkpaint >>
rect -22 -25 110 105
<< ab >>
rect 0 0 88 80
<< pwell >>
rect -4 -7 92 36
<< nwell >>
rect -4 36 92 87
<< polysilicon >>
rect 21 68 23 73
rect 28 68 30 73
rect 35 68 37 73
rect 42 68 44 73
rect 52 68 54 73
rect 59 68 61 73
rect 66 68 68 73
rect 73 68 75 73
rect 9 60 11 65
rect 21 45 23 50
rect 18 44 24 45
rect 9 34 11 42
rect 18 40 19 44
rect 23 40 24 44
rect 18 39 24 40
rect 9 33 15 34
rect 9 29 10 33
rect 14 29 15 33
rect 9 28 15 29
rect 9 25 11 28
rect 21 22 23 39
rect 28 35 30 50
rect 35 41 37 50
rect 42 47 44 50
rect 52 47 54 50
rect 42 46 55 47
rect 42 45 50 46
rect 49 42 50 45
rect 54 42 55 46
rect 49 41 55 42
rect 35 39 45 41
rect 28 34 39 35
rect 28 33 34 34
rect 31 30 34 33
rect 38 30 39 34
rect 31 29 39 30
rect 43 31 45 39
rect 43 30 49 31
rect 31 22 33 29
rect 43 26 44 30
rect 48 26 49 30
rect 43 25 49 26
rect 43 22 45 25
rect 53 22 55 41
rect 59 31 61 50
rect 66 41 68 50
rect 73 47 75 50
rect 73 46 81 47
rect 73 45 76 46
rect 75 42 76 45
rect 80 42 81 46
rect 75 41 81 42
rect 65 40 71 41
rect 65 36 66 40
rect 70 36 71 40
rect 65 35 71 36
rect 59 30 65 31
rect 59 26 60 30
rect 64 26 65 30
rect 59 25 65 26
rect 9 11 11 16
rect 21 11 23 16
rect 31 11 33 16
rect 43 11 45 16
rect 53 11 55 16
<< ndiffusion >>
rect 4 22 9 25
rect 2 21 9 22
rect 2 17 3 21
rect 7 17 9 21
rect 2 16 9 17
rect 11 22 19 25
rect 11 16 21 22
rect 23 21 31 22
rect 23 17 25 21
rect 29 17 31 21
rect 23 16 31 17
rect 33 16 43 22
rect 45 21 53 22
rect 45 17 47 21
rect 51 17 53 21
rect 45 16 53 17
rect 55 16 63 22
rect 13 12 19 16
rect 13 8 14 12
rect 18 8 19 12
rect 35 12 41 16
rect 13 7 19 8
rect 35 8 36 12
rect 40 8 41 12
rect 57 12 63 16
rect 35 7 41 8
rect 57 8 58 12
rect 62 8 63 12
rect 57 7 63 8
<< pdiffusion >>
rect 13 69 19 70
rect 13 65 14 69
rect 18 68 19 69
rect 18 65 21 68
rect 13 60 21 65
rect 4 55 9 60
rect 2 54 9 55
rect 2 50 3 54
rect 7 50 9 54
rect 2 47 9 50
rect 2 43 3 47
rect 7 43 9 47
rect 2 42 9 43
rect 11 50 21 60
rect 23 50 28 68
rect 30 50 35 68
rect 37 50 42 68
rect 44 62 52 68
rect 44 58 46 62
rect 50 58 52 62
rect 44 50 52 58
rect 54 50 59 68
rect 61 50 66 68
rect 68 50 73 68
rect 75 67 82 68
rect 75 63 77 67
rect 81 63 82 67
rect 75 50 82 63
rect 11 42 16 50
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect -2 69 90 78
rect -2 68 14 69
rect 13 65 14 68
rect 18 68 90 69
rect 18 65 19 68
rect 77 67 81 68
rect 2 55 6 63
rect 10 58 46 62
rect 50 58 51 62
rect 2 54 7 55
rect 2 50 3 54
rect 2 47 7 50
rect 2 43 3 47
rect 2 42 7 43
rect 2 22 6 42
rect 10 33 14 58
rect 58 54 62 63
rect 77 62 81 63
rect 18 50 81 54
rect 18 44 23 50
rect 75 46 81 50
rect 18 40 19 44
rect 18 39 23 40
rect 26 42 50 46
rect 54 42 55 46
rect 26 33 30 42
rect 65 40 71 46
rect 75 42 76 46
rect 80 42 81 46
rect 65 38 66 40
rect 34 36 66 38
rect 70 36 71 40
rect 34 34 71 36
rect 14 29 23 32
rect 10 28 23 29
rect 2 21 16 22
rect 2 17 3 21
rect 7 17 16 21
rect 19 21 23 28
rect 34 25 38 30
rect 43 26 44 30
rect 48 26 60 30
rect 64 26 65 30
rect 19 17 25 21
rect 29 17 47 21
rect 51 17 52 21
rect 58 17 62 26
rect -2 8 14 12
rect 18 8 36 12
rect 40 8 58 12
rect 62 8 90 12
rect -2 2 90 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
<< ntransistor >>
rect 9 16 11 25
rect 21 16 23 22
rect 31 16 33 22
rect 43 16 45 22
rect 53 16 55 22
<< ptransistor >>
rect 9 42 11 60
rect 21 50 23 68
rect 28 50 30 68
rect 35 50 37 68
rect 42 50 44 68
rect 52 50 54 68
rect 59 50 61 68
rect 66 50 68 68
rect 73 50 75 68
<< polycontact >>
rect 19 40 23 44
rect 10 29 14 33
rect 50 42 54 46
rect 34 30 38 34
rect 44 26 48 30
rect 76 42 80 46
rect 66 36 70 40
rect 60 26 64 30
<< ndcontact >>
rect 3 17 7 21
rect 25 17 29 21
rect 47 17 51 21
rect 14 8 18 12
rect 36 8 40 12
rect 58 8 62 12
<< pdcontact >>
rect 14 65 18 69
rect 3 50 7 54
rect 3 43 7 47
rect 46 58 50 62
rect 77 63 81 67
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
<< psubstratepdiff >>
rect 0 2 88 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 88 2
rect 0 -3 88 -2
<< nsubstratendiff >>
rect 0 82 88 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 88 82
rect 0 77 88 78
<< labels >>
rlabel polycontact 12 31 12 31 6 zn
rlabel metal1 12 20 12 20 6 z
rlabel metal1 4 40 4 40 6 z
rlabel metal1 12 45 12 45 6 zn
rlabel metal1 20 44 20 44 6 a
rlabel metal1 28 36 28 36 6 d
rlabel metal1 28 52 28 52 6 a
rlabel metal1 44 6 44 6 6 vss
rlabel metal1 36 28 36 28 6 b
rlabel metal1 35 19 35 19 6 zn
rlabel metal1 36 44 36 44 6 d
rlabel metal1 44 36 44 36 6 b
rlabel metal1 44 44 44 44 6 d
rlabel metal1 44 52 44 52 6 a
rlabel metal1 36 52 36 52 6 a
rlabel metal1 30 60 30 60 6 zn
rlabel metal1 44 74 44 74 6 vdd
rlabel metal1 52 28 52 28 6 c
rlabel metal1 60 24 60 24 6 c
rlabel metal1 52 36 52 36 6 b
rlabel polycontact 52 44 52 44 6 d
rlabel metal1 60 36 60 36 6 b
rlabel metal1 68 40 68 40 6 b
rlabel metal1 68 52 68 52 6 a
rlabel metal1 52 52 52 52 6 a
rlabel metal1 60 56 60 56 6 a
rlabel metal1 76 52 76 52 6 a
<< end >>
