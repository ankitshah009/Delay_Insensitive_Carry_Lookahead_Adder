magic
tech scmos
timestamp 1179386000
<< checkpaint >>
rect -22 -25 46 105
<< ab >>
rect 0 0 24 80
<< pwell >>
rect -4 -7 28 36
<< nwell >>
rect -4 36 28 87
<< polysilicon >>
rect 9 70 11 74
rect 9 39 11 42
rect 9 38 22 39
rect 9 37 17 38
rect 9 30 11 37
rect 16 34 17 37
rect 21 34 22 38
rect 16 33 22 34
rect 9 15 11 19
<< ndiffusion >>
rect 2 29 9 30
rect 2 25 3 29
rect 7 25 9 29
rect 2 24 9 25
rect 4 19 9 24
rect 11 19 20 30
rect 13 12 20 19
rect 13 8 14 12
rect 18 8 20 12
rect 13 7 20 8
<< pdiffusion >>
rect 13 72 20 73
rect 13 70 14 72
rect 4 55 9 70
rect 2 54 9 55
rect 2 50 3 54
rect 7 50 9 54
rect 2 47 9 50
rect 2 43 3 47
rect 7 43 9 47
rect 2 42 9 43
rect 11 68 14 70
rect 18 68 20 72
rect 11 42 20 68
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect -2 72 26 78
rect -2 68 14 72
rect 18 68 26 72
rect 2 57 22 63
rect 2 50 3 54
rect 7 50 8 54
rect 2 47 8 50
rect 2 43 3 47
rect 7 43 8 47
rect 2 30 6 43
rect 18 39 22 57
rect 16 38 22 39
rect 16 34 17 38
rect 21 34 22 38
rect 16 33 22 34
rect 2 29 7 30
rect 2 25 3 29
rect 2 23 7 25
rect 2 17 22 23
rect -2 8 14 12
rect 18 8 26 12
rect -2 2 26 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
<< ntransistor >>
rect 9 19 11 30
<< ptransistor >>
rect 9 42 11 70
<< polycontact >>
rect 17 34 21 38
<< ndcontact >>
rect 3 25 7 29
rect 14 8 18 12
<< pdcontact >>
rect 3 50 7 54
rect 3 43 7 47
rect 14 68 18 72
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
<< psubstratepdiff >>
rect 0 2 24 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 24 2
rect 0 -3 24 -2
<< nsubstratendiff >>
rect 0 82 24 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 24 82
rect 0 77 24 78
<< labels >>
rlabel metal1 4 32 4 32 6 z
rlabel metal1 4 60 4 60 6 a
rlabel metal1 12 6 12 6 6 vss
rlabel metal1 12 20 12 20 6 z
rlabel metal1 12 60 12 60 6 a
rlabel metal1 12 74 12 74 6 vdd
rlabel metal1 20 20 20 20 6 z
rlabel metal1 20 48 20 48 6 a
<< end >>
