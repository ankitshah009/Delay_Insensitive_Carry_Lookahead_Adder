magic
tech scmos
timestamp 1185094800
<< checkpaint >>
rect -22 -22 102 122
<< ab >>
rect 0 0 80 100
<< pwell >>
rect -4 -4 84 48
<< nwell >>
rect -4 48 84 104
<< polysilicon >>
rect 25 94 27 98
rect 37 94 39 98
rect 45 94 47 98
rect 57 94 59 98
rect 65 94 67 98
rect 25 52 27 55
rect 25 51 31 52
rect 25 48 26 51
rect 12 47 26 48
rect 30 47 31 51
rect 12 46 31 47
rect 12 36 14 46
rect 37 43 39 55
rect 45 52 47 55
rect 45 51 53 52
rect 45 47 48 51
rect 52 47 53 51
rect 45 46 53 47
rect 35 42 41 43
rect 35 40 36 42
rect 33 38 36 40
rect 40 38 41 42
rect 33 37 41 38
rect 33 34 35 37
rect 45 34 47 46
rect 57 43 59 55
rect 65 52 67 55
rect 65 51 73 52
rect 65 49 68 51
rect 67 47 68 49
rect 72 47 73 51
rect 67 46 73 47
rect 57 42 63 43
rect 57 38 58 42
rect 62 38 63 42
rect 57 37 63 38
rect 57 34 59 37
rect 67 34 69 46
rect 12 12 14 17
rect 33 12 35 17
rect 45 12 47 17
rect 57 12 59 17
rect 67 12 69 17
<< ndiffusion >>
rect 3 32 12 36
rect 3 28 5 32
rect 9 28 12 32
rect 3 22 12 28
rect 3 18 5 22
rect 9 18 12 22
rect 3 17 12 18
rect 14 35 22 36
rect 14 31 17 35
rect 21 31 22 35
rect 14 30 22 31
rect 14 17 19 30
rect 28 23 33 34
rect 25 22 33 23
rect 25 18 26 22
rect 30 18 33 22
rect 25 17 33 18
rect 35 32 45 34
rect 35 28 38 32
rect 42 28 45 32
rect 35 17 45 28
rect 47 22 57 34
rect 47 18 50 22
rect 54 18 57 22
rect 47 17 57 18
rect 59 17 67 34
rect 69 31 74 34
rect 69 30 77 31
rect 69 26 72 30
rect 76 26 77 30
rect 69 22 77 26
rect 69 18 72 22
rect 76 18 77 22
rect 69 17 77 18
rect 61 10 65 17
rect 61 9 67 10
rect 61 5 62 9
rect 66 5 67 9
rect 61 4 67 5
<< pdiffusion >>
rect 20 69 25 94
rect 17 68 25 69
rect 17 64 18 68
rect 22 64 25 68
rect 17 60 25 64
rect 17 56 18 60
rect 22 56 25 60
rect 17 55 25 56
rect 27 92 37 94
rect 27 88 30 92
rect 34 88 37 92
rect 27 82 37 88
rect 27 78 30 82
rect 34 78 37 82
rect 27 55 37 78
rect 39 55 45 94
rect 47 82 57 94
rect 47 78 50 82
rect 54 78 57 82
rect 47 74 57 78
rect 47 70 50 74
rect 54 70 57 74
rect 47 55 57 70
rect 59 55 65 94
rect 67 92 76 94
rect 67 88 70 92
rect 74 88 76 92
rect 67 82 76 88
rect 67 78 70 82
rect 74 78 76 82
rect 67 55 76 78
<< metal1 >>
rect -2 96 82 100
rect -2 92 8 96
rect 12 92 82 96
rect -2 88 30 92
rect 34 88 70 92
rect 74 88 82 92
rect 18 68 22 83
rect 30 82 34 88
rect 30 77 34 78
rect 50 82 54 83
rect 50 74 54 78
rect 70 82 74 88
rect 70 77 74 78
rect 18 60 22 64
rect 18 42 22 56
rect 28 70 50 72
rect 28 68 54 70
rect 28 52 32 68
rect 58 67 72 73
rect 26 51 32 52
rect 30 47 32 51
rect 26 46 32 47
rect 7 38 22 42
rect 17 35 22 38
rect 5 32 9 33
rect 5 22 9 28
rect 21 31 22 35
rect 17 27 22 31
rect 28 32 32 46
rect 38 58 53 63
rect 38 43 42 58
rect 36 42 42 43
rect 40 38 42 42
rect 36 37 42 38
rect 48 51 52 53
rect 48 32 52 47
rect 57 42 62 63
rect 68 51 72 67
rect 68 46 72 47
rect 57 38 58 42
rect 62 38 73 42
rect 28 28 38 32
rect 42 28 43 32
rect 48 27 63 32
rect 71 26 72 30
rect 76 26 77 30
rect 71 22 77 26
rect 25 18 26 22
rect 30 18 50 22
rect 54 18 72 22
rect 76 18 77 22
rect 5 12 9 18
rect -2 9 82 12
rect -2 8 62 9
rect -2 4 8 8
rect 12 4 18 8
rect 22 5 62 8
rect 66 5 82 9
rect 22 4 82 5
rect -2 0 82 4
<< ntransistor >>
rect 12 17 14 36
rect 33 17 35 34
rect 45 17 47 34
rect 57 17 59 34
rect 67 17 69 34
<< ptransistor >>
rect 25 55 27 94
rect 37 55 39 94
rect 45 55 47 94
rect 57 55 59 94
rect 65 55 67 94
<< polycontact >>
rect 26 47 30 51
rect 48 47 52 51
rect 36 38 40 42
rect 68 47 72 51
rect 58 38 62 42
<< ndcontact >>
rect 5 28 9 32
rect 5 18 9 22
rect 17 31 21 35
rect 26 18 30 22
rect 38 28 42 32
rect 50 18 54 22
rect 72 26 76 30
rect 72 18 76 22
rect 62 5 66 9
<< pdcontact >>
rect 18 64 22 68
rect 18 56 22 60
rect 30 88 34 92
rect 30 78 34 82
rect 50 78 54 82
rect 50 70 54 74
rect 70 88 74 92
rect 70 78 74 82
<< psubstratepcontact >>
rect 8 4 12 8
rect 18 4 22 8
<< nsubstratencontact >>
rect 8 92 12 96
<< psubstratepdiff >>
rect 7 8 23 9
rect 7 4 8 8
rect 12 4 18 8
rect 22 4 23 8
rect 7 3 23 4
<< nsubstratendiff >>
rect 7 96 13 97
rect 7 92 8 96
rect 12 92 13 96
rect 7 91 13 92
<< labels >>
rlabel polycontact 28 49 28 49 6 zn
rlabel metal1 10 40 10 40 6 z
rlabel metal1 20 55 20 55 6 z
rlabel metal1 40 6 40 6 6 vss
rlabel metal1 35 30 35 30 6 zn
rlabel polycontact 29 49 29 49 6 zn
rlabel metal1 40 50 40 50 6 b1
rlabel metal1 40 94 40 94 6 vdd
rlabel metal1 60 30 60 30 6 b2
rlabel metal1 50 40 50 40 6 b2
rlabel metal1 60 50 60 50 6 a2
rlabel metal1 50 60 50 60 6 b1
rlabel metal1 60 70 60 70 6 a1
rlabel metal1 52 75 52 75 6 zn
rlabel metal1 74 24 74 24 6 n3
rlabel ndcontact 51 20 51 20 6 n3
rlabel metal1 70 40 70 40 6 a2
rlabel metal1 70 60 70 60 6 a1
<< end >>
