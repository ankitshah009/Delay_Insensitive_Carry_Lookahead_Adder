magic
tech scmos
timestamp 1180640021
<< checkpaint >>
rect -24 -26 174 126
<< ab >>
rect 0 0 150 100
<< pwell >>
rect -4 -6 154 49
<< nwell >>
rect -4 49 154 106
<< polysilicon >>
rect 123 93 125 98
rect 135 93 137 98
rect 11 87 13 92
rect 23 87 25 92
rect 35 87 37 92
rect 47 87 49 92
rect 59 87 61 92
rect 67 87 69 92
rect 79 87 81 92
rect 87 87 89 92
rect 99 87 101 92
rect 111 87 113 92
rect 11 53 13 56
rect 7 52 13 53
rect 7 48 8 52
rect 12 48 13 52
rect 7 47 13 48
rect 11 33 13 47
rect 23 53 25 56
rect 35 53 37 56
rect 23 52 37 53
rect 23 48 28 52
rect 32 48 37 52
rect 47 53 49 56
rect 59 53 61 56
rect 47 52 63 53
rect 47 51 58 52
rect 23 47 37 48
rect 57 48 58 51
rect 62 48 63 52
rect 57 47 63 48
rect 23 33 25 47
rect 35 33 37 47
rect 47 42 53 43
rect 47 38 48 42
rect 52 38 53 42
rect 47 37 53 38
rect 47 33 49 37
rect 59 33 61 47
rect 67 43 69 56
rect 79 43 81 56
rect 67 42 81 43
rect 67 38 72 42
rect 76 38 81 42
rect 67 37 81 38
rect 67 33 69 37
rect 79 33 81 37
rect 87 53 89 56
rect 99 53 101 56
rect 111 53 113 56
rect 87 52 93 53
rect 87 48 88 52
rect 92 48 93 52
rect 87 47 93 48
rect 97 52 113 53
rect 97 48 98 52
rect 102 51 113 52
rect 102 48 103 51
rect 97 47 103 48
rect 123 47 125 56
rect 135 47 137 56
rect 87 33 89 47
rect 118 46 137 47
rect 118 42 119 46
rect 123 45 137 46
rect 123 42 125 45
rect 118 41 125 42
rect 123 37 125 41
rect 135 37 137 45
rect 23 14 25 19
rect 35 14 37 19
rect 59 14 61 19
rect 67 14 69 19
rect 79 14 81 19
rect 87 14 89 19
rect 123 14 125 19
rect 135 14 137 19
rect 11 2 13 6
rect 47 2 49 6
<< ndiffusion >>
rect 3 32 11 33
rect 3 28 4 32
rect 8 28 11 32
rect 3 22 11 28
rect 3 18 4 22
rect 8 18 11 22
rect 3 12 11 18
rect 3 8 4 12
rect 8 8 11 12
rect 3 6 11 8
rect 13 32 23 33
rect 13 28 16 32
rect 20 28 23 32
rect 13 24 23 28
rect 13 20 16 24
rect 20 20 23 24
rect 13 19 23 20
rect 25 32 35 33
rect 25 28 28 32
rect 32 28 35 32
rect 25 19 35 28
rect 37 24 47 33
rect 37 20 40 24
rect 44 20 47 24
rect 37 19 47 20
rect 13 6 18 19
rect 42 6 47 19
rect 49 22 59 33
rect 49 18 52 22
rect 56 19 59 22
rect 61 19 67 33
rect 69 32 79 33
rect 69 28 72 32
rect 76 28 79 32
rect 69 24 79 28
rect 69 20 72 24
rect 76 20 79 24
rect 69 19 79 20
rect 81 19 87 33
rect 89 24 98 33
rect 89 20 92 24
rect 96 20 98 24
rect 89 19 98 20
rect 114 32 123 37
rect 114 28 116 32
rect 120 28 123 32
rect 114 24 123 28
rect 114 20 116 24
rect 120 20 123 24
rect 114 19 123 20
rect 125 36 135 37
rect 125 32 128 36
rect 132 32 135 36
rect 125 28 135 32
rect 125 24 128 28
rect 132 24 135 28
rect 125 19 135 24
rect 137 32 146 37
rect 137 28 140 32
rect 144 28 146 32
rect 137 24 146 28
rect 137 20 140 24
rect 144 20 146 24
rect 137 19 146 20
rect 56 18 57 19
rect 49 12 57 18
rect 49 8 52 12
rect 56 8 57 12
rect 49 6 57 8
<< pdiffusion >>
rect 51 92 57 93
rect 91 92 97 93
rect 115 92 123 93
rect 51 88 52 92
rect 56 88 57 92
rect 51 87 57 88
rect 91 88 92 92
rect 96 88 97 92
rect 91 87 97 88
rect 115 88 116 92
rect 120 88 123 92
rect 115 87 123 88
rect 3 82 11 87
rect 3 78 4 82
rect 8 78 11 82
rect 3 56 11 78
rect 13 82 23 87
rect 13 78 16 82
rect 20 78 23 82
rect 13 56 23 78
rect 25 62 35 87
rect 25 58 28 62
rect 32 58 35 62
rect 25 56 35 58
rect 37 82 47 87
rect 37 78 40 82
rect 44 78 47 82
rect 37 56 47 78
rect 49 56 59 87
rect 61 56 67 87
rect 69 62 79 87
rect 69 58 72 62
rect 76 58 79 62
rect 69 56 79 58
rect 81 56 87 87
rect 89 56 99 87
rect 101 80 111 87
rect 101 76 104 80
rect 108 76 111 80
rect 101 72 111 76
rect 101 68 104 72
rect 108 68 111 72
rect 101 56 111 68
rect 113 82 123 87
rect 113 78 116 82
rect 120 78 123 82
rect 113 72 123 78
rect 113 68 116 72
rect 120 68 123 72
rect 113 56 123 68
rect 125 72 135 93
rect 125 68 128 72
rect 132 68 135 72
rect 125 62 135 68
rect 125 58 128 62
rect 132 58 135 62
rect 125 56 135 58
rect 137 92 146 93
rect 137 88 140 92
rect 144 88 146 92
rect 137 82 146 88
rect 137 78 140 82
rect 144 78 146 82
rect 137 72 146 78
rect 137 68 140 72
rect 144 68 146 72
rect 137 56 146 68
<< metal1 >>
rect -2 92 152 100
rect -2 88 52 92
rect 56 88 92 92
rect 96 88 116 92
rect 120 88 140 92
rect 144 88 152 92
rect 4 82 8 88
rect 116 82 120 88
rect 15 78 16 82
rect 20 78 40 82
rect 44 80 108 82
rect 44 78 104 80
rect 4 77 8 78
rect 104 72 108 76
rect 8 68 93 72
rect 8 52 12 68
rect 8 47 12 48
rect 18 52 22 63
rect 27 58 28 62
rect 32 58 72 62
rect 76 58 77 62
rect 18 48 28 52
rect 32 48 33 52
rect 18 37 22 48
rect 4 32 8 33
rect 38 32 42 58
rect 87 52 93 68
rect 104 67 108 68
rect 116 72 120 78
rect 140 82 144 88
rect 116 67 120 68
rect 128 72 132 73
rect 128 62 132 68
rect 140 72 144 78
rect 140 67 144 68
rect 57 48 58 52
rect 62 48 88 52
rect 92 48 93 52
rect 97 52 103 62
rect 97 48 98 52
rect 102 48 103 52
rect 97 42 103 48
rect 128 52 132 58
rect 128 48 143 52
rect 47 38 48 42
rect 52 38 72 42
rect 76 38 103 42
rect 108 42 119 46
rect 123 42 124 46
rect 108 32 112 42
rect 128 36 132 48
rect 4 22 8 28
rect 15 28 16 32
rect 20 28 21 32
rect 27 28 28 32
rect 32 28 72 32
rect 76 28 112 32
rect 116 32 120 33
rect 15 24 21 28
rect 72 24 76 28
rect 116 24 120 28
rect 15 20 16 24
rect 20 20 40 24
rect 44 20 45 24
rect 52 22 56 23
rect 4 12 8 18
rect 72 19 76 20
rect 91 20 92 24
rect 96 20 97 24
rect 52 12 56 18
rect 91 12 97 20
rect 128 28 132 32
rect 128 23 132 24
rect 140 32 144 33
rect 140 24 144 28
rect 116 12 120 20
rect 140 12 144 20
rect -2 8 4 12
rect 8 8 52 12
rect 56 8 152 12
rect -2 0 152 8
<< ntransistor >>
rect 11 6 13 33
rect 23 19 25 33
rect 35 19 37 33
rect 47 6 49 33
rect 59 19 61 33
rect 67 19 69 33
rect 79 19 81 33
rect 87 19 89 33
rect 123 19 125 37
rect 135 19 137 37
<< ptransistor >>
rect 11 56 13 87
rect 23 56 25 87
rect 35 56 37 87
rect 47 56 49 87
rect 59 56 61 87
rect 67 56 69 87
rect 79 56 81 87
rect 87 56 89 87
rect 99 56 101 87
rect 111 56 113 87
rect 123 56 125 93
rect 135 56 137 93
<< polycontact >>
rect 8 48 12 52
rect 28 48 32 52
rect 58 48 62 52
rect 48 38 52 42
rect 72 38 76 42
rect 88 48 92 52
rect 98 48 102 52
rect 119 42 123 46
<< ndcontact >>
rect 4 28 8 32
rect 4 18 8 22
rect 4 8 8 12
rect 16 28 20 32
rect 16 20 20 24
rect 28 28 32 32
rect 40 20 44 24
rect 52 18 56 22
rect 72 28 76 32
rect 72 20 76 24
rect 92 20 96 24
rect 116 28 120 32
rect 116 20 120 24
rect 128 32 132 36
rect 128 24 132 28
rect 140 28 144 32
rect 140 20 144 24
rect 52 8 56 12
<< pdcontact >>
rect 52 88 56 92
rect 92 88 96 92
rect 116 88 120 92
rect 4 78 8 82
rect 16 78 20 82
rect 28 58 32 62
rect 40 78 44 82
rect 72 58 76 62
rect 104 76 108 80
rect 104 68 108 72
rect 116 78 120 82
rect 116 68 120 72
rect 128 68 132 72
rect 128 58 132 62
rect 140 88 144 92
rect 140 78 144 82
rect 140 68 144 72
<< psubstratepcontact >>
rect 108 4 112 8
rect 118 4 122 8
<< psubstratepdiff >>
rect 107 8 123 9
rect 107 4 108 8
rect 112 4 118 8
rect 122 4 123 8
rect 107 3 123 4
<< labels >>
rlabel polycontact 121 44 121 44 6 zn
rlabel metal1 18 26 18 26 6 n4
rlabel metal1 20 50 20 50 6 c
rlabel metal1 20 50 20 50 6 c
rlabel metal1 10 60 10 60 6 a
rlabel metal1 10 60 10 60 6 a
rlabel metal1 20 70 20 70 6 a
rlabel metal1 20 70 20 70 6 a
rlabel metal1 30 22 30 22 6 n4
rlabel polycontact 50 40 50 40 6 b
rlabel polycontact 50 40 50 40 6 b
rlabel polycontact 30 50 30 50 6 c
rlabel polycontact 30 50 30 50 6 c
rlabel metal1 30 70 30 70 6 a
rlabel metal1 30 70 30 70 6 a
rlabel metal1 40 70 40 70 6 a
rlabel metal1 50 70 50 70 6 a
rlabel metal1 40 70 40 70 6 a
rlabel metal1 50 70 50 70 6 a
rlabel metal1 75 6 75 6 6 vss
rlabel metal1 75 6 75 6 6 vss
rlabel metal1 74 25 74 25 6 zn
rlabel metal1 70 40 70 40 6 b
rlabel metal1 80 40 80 40 6 b
rlabel metal1 70 40 70 40 6 b
rlabel metal1 80 40 80 40 6 b
rlabel metal1 60 40 60 40 6 b
rlabel metal1 60 40 60 40 6 b
rlabel polycontact 60 50 60 50 6 a
rlabel polycontact 60 50 60 50 6 a
rlabel metal1 80 50 80 50 6 a
rlabel metal1 70 50 70 50 6 a
rlabel metal1 70 50 70 50 6 a
rlabel metal1 80 50 80 50 6 a
rlabel metal1 52 60 52 60 6 zn
rlabel metal1 60 70 60 70 6 a
rlabel metal1 60 70 60 70 6 a
rlabel metal1 80 70 80 70 6 a
rlabel metal1 70 70 70 70 6 a
rlabel metal1 70 70 70 70 6 a
rlabel metal1 80 70 80 70 6 a
rlabel metal1 75 94 75 94 6 vdd
rlabel metal1 75 94 75 94 6 vdd
rlabel metal1 69 30 69 30 6 zn
rlabel metal1 90 40 90 40 6 b
rlabel metal1 90 40 90 40 6 b
rlabel polycontact 100 50 100 50 6 b
rlabel polycontact 100 50 100 50 6 b
rlabel metal1 90 60 90 60 6 a
rlabel metal1 90 60 90 60 6 a
rlabel metal1 106 74 106 74 6 n2
rlabel metal1 61 80 61 80 6 n2
rlabel metal1 116 44 116 44 6 zn
rlabel metal1 130 50 130 50 6 z
rlabel metal1 140 50 140 50 6 z
rlabel metal1 130 50 130 50 6 z
rlabel metal1 140 50 140 50 6 z
<< end >>
