magic
tech scmos
timestamp 1179387411
<< checkpaint >>
rect -22 -25 102 105
<< ab >>
rect 0 0 80 80
<< pwell >>
rect -4 -7 84 36
<< nwell >>
rect -4 36 84 87
<< polysilicon >>
rect 9 70 11 74
rect 27 70 29 74
rect 37 70 39 74
rect 44 70 46 74
rect 57 70 59 74
rect 67 70 69 74
rect 9 39 11 42
rect 27 39 29 42
rect 9 38 29 39
rect 9 34 10 38
rect 14 37 29 38
rect 14 34 15 37
rect 37 35 39 42
rect 44 39 46 42
rect 57 39 59 42
rect 9 33 15 34
rect 33 34 39 35
rect 11 26 13 33
rect 33 31 34 34
rect 21 30 34 31
rect 38 30 39 34
rect 43 38 49 39
rect 43 34 44 38
rect 48 35 49 38
rect 57 38 63 39
rect 48 34 52 35
rect 43 33 52 34
rect 57 34 58 38
rect 62 34 63 38
rect 57 33 63 34
rect 67 36 69 42
rect 67 35 73 36
rect 21 29 39 30
rect 21 26 23 29
rect 50 27 52 33
rect 60 27 62 33
rect 67 31 68 35
rect 72 31 73 35
rect 67 30 73 31
rect 67 27 69 30
rect 11 8 13 13
rect 21 8 23 13
rect 50 6 52 10
rect 60 6 62 10
rect 67 6 69 10
<< ndiffusion >>
rect 4 18 11 26
rect 4 14 5 18
rect 9 14 11 18
rect 4 13 11 14
rect 13 25 21 26
rect 13 21 15 25
rect 19 21 21 25
rect 13 13 21 21
rect 23 25 31 26
rect 23 21 26 25
rect 30 21 31 25
rect 45 23 50 27
rect 23 20 31 21
rect 42 22 50 23
rect 23 13 28 20
rect 42 18 43 22
rect 47 18 50 22
rect 42 17 50 18
rect 45 10 50 17
rect 52 26 60 27
rect 52 22 54 26
rect 58 22 60 26
rect 52 10 60 22
rect 62 10 67 27
rect 69 15 76 27
rect 69 11 71 15
rect 75 11 76 15
rect 69 10 76 11
<< pdiffusion >>
rect 2 69 9 70
rect 2 65 3 69
rect 7 65 9 69
rect 2 62 9 65
rect 2 58 3 62
rect 7 58 9 62
rect 2 42 9 58
rect 11 48 16 70
rect 22 63 27 70
rect 20 62 27 63
rect 20 58 21 62
rect 25 58 27 62
rect 20 57 27 58
rect 11 47 18 48
rect 11 43 13 47
rect 17 43 18 47
rect 11 42 18 43
rect 22 42 27 57
rect 29 47 37 70
rect 29 43 31 47
rect 35 43 37 47
rect 29 42 37 43
rect 39 42 44 70
rect 46 69 57 70
rect 46 65 49 69
rect 53 65 57 69
rect 46 42 57 65
rect 59 62 67 70
rect 59 58 61 62
rect 65 58 67 62
rect 59 55 67 58
rect 59 51 61 55
rect 65 51 67 55
rect 59 42 67 51
rect 69 69 77 70
rect 69 65 71 69
rect 75 65 77 69
rect 69 62 77 65
rect 69 58 71 62
rect 75 58 77 62
rect 69 42 77 58
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect -2 69 82 78
rect -2 68 3 69
rect 2 65 3 68
rect 7 68 49 69
rect 7 65 8 68
rect 48 65 49 68
rect 53 68 71 69
rect 53 65 54 68
rect 70 65 71 68
rect 75 68 82 69
rect 75 65 76 68
rect 2 62 8 65
rect 61 62 66 63
rect 2 58 3 62
rect 7 58 8 62
rect 20 58 21 62
rect 25 58 55 62
rect 51 55 55 58
rect 65 58 66 62
rect 70 62 76 65
rect 70 58 71 62
rect 75 58 76 62
rect 61 55 66 58
rect 18 50 46 54
rect 18 47 22 50
rect 2 39 6 47
rect 12 43 13 47
rect 17 43 22 47
rect 2 38 14 39
rect 2 34 10 38
rect 2 33 14 34
rect 2 25 6 33
rect 18 25 22 43
rect 14 21 15 25
rect 19 21 22 25
rect 26 43 31 47
rect 35 43 36 47
rect 26 25 30 43
rect 42 39 46 50
rect 51 51 61 55
rect 65 51 66 55
rect 42 38 48 39
rect 34 34 38 35
rect 42 34 44 38
rect 42 33 48 34
rect 51 30 55 51
rect 58 41 78 47
rect 58 38 62 41
rect 58 33 62 34
rect 68 35 72 36
rect 34 26 55 30
rect 66 29 78 31
rect 51 22 54 26
rect 58 22 59 26
rect 65 25 78 29
rect 30 21 43 22
rect 5 18 9 19
rect 26 18 43 21
rect 47 18 48 22
rect 65 18 71 25
rect 5 12 9 14
rect 70 12 71 15
rect -2 11 71 12
rect 75 12 76 15
rect 75 11 82 12
rect -2 2 82 11
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
<< ntransistor >>
rect 11 13 13 26
rect 21 13 23 26
rect 50 10 52 27
rect 60 10 62 27
rect 67 10 69 27
<< ptransistor >>
rect 9 42 11 70
rect 27 42 29 70
rect 37 42 39 70
rect 44 42 46 70
rect 57 42 59 70
rect 67 42 69 70
<< polycontact >>
rect 10 34 14 38
rect 34 30 38 34
rect 44 34 48 38
rect 58 34 62 38
rect 68 31 72 35
<< ndcontact >>
rect 5 14 9 18
rect 15 21 19 25
rect 26 21 30 25
rect 43 18 47 22
rect 54 22 58 26
rect 71 11 75 15
<< pdcontact >>
rect 3 65 7 69
rect 3 58 7 62
rect 21 58 25 62
rect 13 43 17 47
rect 31 43 35 47
rect 49 65 53 69
rect 61 58 65 62
rect 61 51 65 55
rect 71 65 75 69
rect 71 58 75 62
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
<< psubstratepdiff >>
rect 0 2 80 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 80 2
rect 0 -3 80 -2
<< nsubstratendiff >>
rect 0 82 80 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 80 82
rect 0 77 80 78
<< labels >>
rlabel polycontact 36 32 36 32 6 an
rlabel ptransistor 45 53 45 53 6 bn
rlabel metal1 4 36 4 36 6 b
rlabel polycontact 12 36 12 36 6 b
rlabel metal1 17 45 17 45 6 bn
rlabel metal1 28 36 28 36 6 z
rlabel metal1 20 37 20 37 6 bn
rlabel metal1 40 6 40 6 6 vss
rlabel ndcontact 44 20 44 20 6 z
rlabel metal1 36 20 36 20 6 z
rlabel metal1 36 30 36 30 6 an
rlabel metal1 40 74 40 74 6 vdd
rlabel polycontact 45 36 45 36 6 bn
rlabel metal1 60 40 60 40 6 a2
rlabel metal1 53 42 53 42 6 an
rlabel metal1 37 60 37 60 6 an
rlabel metal1 68 24 68 24 6 a1
rlabel metal1 76 28 76 28 6 a1
rlabel metal1 68 44 68 44 6 a2
rlabel metal1 76 44 76 44 6 a2
rlabel metal1 63 57 63 57 6 an
<< end >>
