magic
tech scmos
timestamp 1179386995
<< checkpaint >>
rect -22 -25 86 105
<< ab >>
rect 0 0 64 80
<< pwell >>
rect -4 -7 68 36
<< nwell >>
rect -4 36 68 87
<< polysilicon >>
rect 12 70 14 74
rect 22 70 24 74
rect 29 70 31 74
rect 12 49 14 55
rect 9 48 15 49
rect 9 44 10 48
rect 14 44 15 48
rect 9 43 15 44
rect 9 23 11 43
rect 39 68 41 72
rect 39 47 41 50
rect 39 46 55 47
rect 39 45 50 46
rect 49 42 50 45
rect 54 42 55 46
rect 22 39 24 42
rect 17 38 24 39
rect 17 34 18 38
rect 22 34 24 38
rect 17 33 24 34
rect 29 39 31 42
rect 49 41 55 42
rect 29 38 35 39
rect 29 34 30 38
rect 34 34 35 38
rect 29 33 35 34
rect 19 23 21 33
rect 29 23 31 33
rect 49 30 51 41
rect 49 16 51 21
rect 9 6 11 10
rect 19 6 21 10
rect 29 6 31 10
<< ndiffusion >>
rect 42 29 49 30
rect 42 25 43 29
rect 47 25 49 29
rect 42 24 49 25
rect 2 22 9 23
rect 2 18 3 22
rect 7 18 9 22
rect 2 17 9 18
rect 4 10 9 17
rect 11 22 19 23
rect 11 18 13 22
rect 17 18 19 22
rect 11 10 19 18
rect 21 15 29 23
rect 21 11 23 15
rect 27 11 29 15
rect 21 10 29 11
rect 31 22 38 23
rect 31 18 33 22
rect 37 18 38 22
rect 44 21 49 24
rect 51 26 58 30
rect 51 22 53 26
rect 57 22 58 26
rect 51 21 58 22
rect 31 17 38 18
rect 31 10 36 17
<< pdiffusion >>
rect 4 69 12 70
rect 4 65 6 69
rect 10 65 12 69
rect 4 55 12 65
rect 14 62 22 70
rect 14 58 16 62
rect 20 58 22 62
rect 14 55 22 58
rect 17 42 22 55
rect 24 42 29 70
rect 31 68 37 70
rect 31 67 39 68
rect 31 63 33 67
rect 37 63 39 67
rect 31 60 39 63
rect 31 56 33 60
rect 37 56 39 60
rect 31 50 39 56
rect 41 63 46 68
rect 41 62 48 63
rect 41 58 43 62
rect 47 58 48 62
rect 41 55 48 58
rect 41 51 43 55
rect 47 51 48 55
rect 41 50 48 51
rect 31 42 37 50
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect -2 69 66 78
rect -2 68 6 69
rect 5 65 6 68
rect 10 68 66 69
rect 10 65 11 68
rect 33 67 37 68
rect 2 58 16 62
rect 20 58 23 62
rect 33 60 37 63
rect 2 22 6 58
rect 33 55 37 56
rect 43 62 47 63
rect 43 55 47 58
rect 10 48 14 49
rect 43 46 47 51
rect 58 47 62 55
rect 10 30 14 44
rect 18 42 47 46
rect 18 38 22 42
rect 25 34 30 38
rect 34 34 39 38
rect 18 33 22 34
rect 10 26 23 30
rect 33 26 39 34
rect 43 29 47 42
rect 50 46 62 47
rect 54 42 62 46
rect 50 41 62 42
rect 43 24 47 25
rect 53 26 57 27
rect 2 18 3 22
rect 7 18 8 22
rect 12 18 13 22
rect 17 18 33 22
rect 37 18 38 22
rect 2 17 8 18
rect 22 12 23 15
rect -2 11 23 12
rect 27 12 28 15
rect 53 12 57 22
rect 27 11 66 12
rect -2 2 66 11
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
<< ntransistor >>
rect 9 10 11 23
rect 19 10 21 23
rect 29 10 31 23
rect 49 21 51 30
<< ptransistor >>
rect 12 55 14 70
rect 22 42 24 70
rect 29 42 31 70
rect 39 50 41 68
<< polycontact >>
rect 10 44 14 48
rect 50 42 54 46
rect 18 34 22 38
rect 30 34 34 38
<< ndcontact >>
rect 43 25 47 29
rect 3 18 7 22
rect 13 18 17 22
rect 23 11 27 15
rect 33 18 37 22
rect 53 22 57 26
<< pdcontact >>
rect 6 65 10 69
rect 16 58 20 62
rect 33 63 37 67
rect 33 56 37 60
rect 43 58 47 62
rect 43 51 47 55
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
<< psubstratepdiff >>
rect 0 2 64 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 64 2
rect 0 -3 64 -2
<< nsubstratendiff >>
rect 0 82 64 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 64 82
rect 0 77 64 78
<< labels >>
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 40 12 40 6 b
rlabel metal1 12 60 12 60 6 z
rlabel metal1 20 28 20 28 6 b
rlabel metal1 28 36 28 36 6 a1
rlabel metal1 20 60 20 60 6 z
rlabel metal1 32 6 32 6 6 vss
rlabel metal1 25 20 25 20 6 n1
rlabel metal1 36 32 36 32 6 a1
rlabel metal1 32 74 32 74 6 vdd
rlabel polycontact 52 44 52 44 6 a2
rlabel metal1 60 48 60 48 6 a2
<< end >>
