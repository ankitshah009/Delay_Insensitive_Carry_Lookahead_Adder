magic
tech scmos
timestamp 1182081791
<< checkpaint >>
rect -25 -26 57 114
<< ab >>
rect 0 0 32 88
<< pwell >>
rect -7 -8 39 40
<< nwell >>
rect -7 40 39 96
<< polysilicon >>
rect 5 80 14 86
rect 18 80 27 86
rect 9 77 11 80
rect 21 77 23 80
rect 9 48 11 51
rect 21 48 23 51
rect 2 47 11 48
rect 2 43 6 47
rect 10 43 11 47
rect 2 42 11 43
rect 15 47 30 48
rect 15 43 22 47
rect 26 43 30 47
rect 15 42 30 43
rect 2 37 17 38
rect 2 33 6 37
rect 10 33 17 37
rect 2 32 17 33
rect 21 37 30 38
rect 21 33 22 37
rect 26 33 30 37
rect 21 32 30 33
rect 9 29 11 32
rect 21 29 23 32
rect 9 8 11 11
rect 21 8 23 11
rect 5 2 14 8
rect 18 2 27 8
<< ndiffusion >>
rect 2 24 9 29
rect 2 20 3 24
rect 7 20 9 24
rect 2 17 9 20
rect 2 13 3 17
rect 7 13 9 17
rect 2 11 9 13
rect 11 11 21 29
rect 23 25 30 29
rect 23 21 25 25
rect 29 21 30 25
rect 23 18 30 21
rect 23 14 25 18
rect 29 14 30 18
rect 23 11 30 14
<< pdiffusion >>
rect 2 75 9 77
rect 2 71 3 75
rect 7 71 9 75
rect 2 68 9 71
rect 2 64 3 68
rect 7 64 9 68
rect 2 51 9 64
rect 11 66 21 77
rect 11 62 14 66
rect 18 62 21 66
rect 11 58 21 62
rect 11 54 14 58
rect 18 54 21 58
rect 11 51 21 54
rect 23 75 30 77
rect 23 71 25 75
rect 29 71 30 75
rect 23 68 30 71
rect 23 64 25 68
rect 29 64 30 68
rect 23 51 30 64
<< metal1 >>
rect -2 86 2 90
rect 30 86 34 90
rect 2 82 7 85
rect -2 81 7 82
rect 3 75 7 81
rect 3 68 7 71
rect 25 82 30 85
rect 25 81 34 82
rect 25 75 29 81
rect 25 68 29 71
rect 3 63 7 64
rect 14 66 18 67
rect 25 63 29 64
rect 14 58 18 62
rect 6 47 10 51
rect 6 37 10 43
rect 6 29 10 33
rect 14 26 18 54
rect 22 47 26 59
rect 22 37 26 43
rect 22 32 26 33
rect 14 25 29 26
rect 3 24 7 25
rect 14 21 25 25
rect 3 17 7 20
rect 22 18 29 21
rect 22 14 25 18
rect 22 13 29 14
rect 3 7 7 13
rect -2 6 7 7
rect 2 3 7 6
rect 30 6 34 7
rect -2 -2 2 2
rect 30 -2 34 2
<< metal2 >>
rect -2 86 34 90
rect 2 82 30 86
rect -2 80 34 82
rect -2 6 34 8
rect 2 2 30 6
rect -2 -2 34 2
<< ntransistor >>
rect 9 11 11 29
rect 21 11 23 29
<< ptransistor >>
rect 9 51 11 77
rect 21 51 23 77
<< polycontact >>
rect 6 43 10 47
rect 22 43 26 47
rect 6 33 10 37
rect 22 33 26 37
<< ndcontact >>
rect 3 20 7 24
rect 3 13 7 17
rect 25 21 29 25
rect 25 14 29 18
<< pdcontact >>
rect 3 71 7 75
rect 3 64 7 68
rect 14 62 18 66
rect 14 54 18 58
rect 25 71 29 75
rect 25 64 29 68
<< m2contact >>
rect -2 82 2 86
rect 30 82 34 86
rect -2 2 2 6
rect 30 2 34 6
<< psubstratepcontact >>
rect -2 2 2 6
rect 30 2 34 6
<< nsubstratencontact >>
rect -2 82 2 86
rect 30 82 34 86
<< psubstratepdiff >>
rect -3 6 3 7
rect -3 2 -2 6
rect 2 2 3 6
rect 29 6 35 7
rect 29 2 30 6
rect 34 2 35 6
rect -3 0 3 2
rect 29 0 35 2
<< nsubstratendiff >>
rect -3 86 3 88
rect 29 86 35 88
rect -3 82 -2 86
rect 2 82 3 86
rect -3 81 3 82
rect 29 82 30 86
rect 34 82 35 86
rect 29 81 35 82
<< labels >>
rlabel metal1 8 40 8 40 6 a
rlabel metal1 16 44 16 44 6 z
rlabel metal1 24 20 24 20 6 z
rlabel metal1 24 48 24 48 6 b
rlabel metal2 16 4 16 4 6 vss
rlabel metal2 16 84 16 84 6 vdd
<< end >>
