magic
tech scmos
timestamp 1179387611
<< checkpaint >>
rect -22 -22 158 94
<< ab >>
rect 0 0 136 72
<< pwell >>
rect -4 -4 140 32
<< nwell >>
rect -4 32 140 76
<< polysilicon >>
rect 9 66 11 70
rect 19 66 21 70
rect 29 66 31 70
rect 39 66 41 70
rect 49 66 51 70
rect 59 66 61 70
rect 66 66 68 70
rect 78 68 104 70
rect 78 59 80 68
rect 85 62 97 64
rect 85 59 87 62
rect 95 59 97 62
rect 102 59 104 68
rect 115 66 117 70
rect 125 57 127 61
rect 9 35 11 38
rect 19 35 21 38
rect 29 35 31 38
rect 39 35 41 38
rect 49 35 51 38
rect 59 35 61 38
rect 9 33 21 35
rect 25 34 51 35
rect 9 32 15 33
rect 9 28 10 32
rect 14 28 15 32
rect 25 30 26 34
rect 30 33 51 34
rect 55 34 61 35
rect 30 30 31 33
rect 25 29 31 30
rect 55 30 56 34
rect 60 30 61 34
rect 66 35 68 38
rect 78 35 80 38
rect 66 33 80 35
rect 85 35 87 38
rect 85 34 91 35
rect 95 34 97 38
rect 102 35 104 38
rect 115 35 117 38
rect 125 35 127 38
rect 101 34 107 35
rect 55 29 61 30
rect 85 30 86 34
rect 90 30 91 34
rect 101 30 102 34
rect 106 30 107 34
rect 85 29 91 30
rect 9 27 15 28
rect 19 27 31 29
rect 12 24 14 27
rect 19 24 21 27
rect 29 24 31 27
rect 36 24 38 29
rect 55 26 57 29
rect 12 4 14 12
rect 19 8 21 12
rect 29 8 31 12
rect 36 4 38 12
rect 12 2 38 4
rect 75 25 77 29
rect 85 25 87 29
rect 95 28 107 30
rect 95 25 97 28
rect 105 25 107 28
rect 115 34 127 35
rect 115 30 122 34
rect 126 30 127 34
rect 115 29 127 30
rect 115 26 117 29
rect 125 26 127 29
rect 55 6 57 11
rect 125 12 127 16
rect 85 8 87 12
rect 95 8 97 12
rect 105 8 107 12
rect 75 4 77 7
rect 115 4 117 12
rect 75 2 117 4
<< ndiffusion >>
rect 40 24 55 26
rect 3 12 12 24
rect 14 12 19 24
rect 21 18 29 24
rect 21 14 23 18
rect 27 14 29 18
rect 21 12 29 14
rect 31 12 36 24
rect 38 12 55 24
rect 3 8 10 12
rect 3 4 5 8
rect 9 4 10 8
rect 3 3 10 4
rect 40 11 55 12
rect 57 25 64 26
rect 109 25 115 26
rect 57 21 59 25
rect 63 21 64 25
rect 57 20 64 21
rect 57 11 62 20
rect 70 19 75 25
rect 68 18 75 19
rect 68 14 69 18
rect 73 14 75 18
rect 68 13 75 14
rect 40 8 53 11
rect 40 4 41 8
rect 45 4 48 8
rect 52 4 53 8
rect 70 7 75 13
rect 77 24 85 25
rect 77 20 79 24
rect 83 20 85 24
rect 77 17 85 20
rect 77 13 79 17
rect 83 13 85 17
rect 77 12 85 13
rect 87 17 95 25
rect 87 13 89 17
rect 93 13 95 17
rect 87 12 95 13
rect 97 24 105 25
rect 97 20 99 24
rect 103 20 105 24
rect 97 17 105 20
rect 97 13 99 17
rect 103 13 105 17
rect 97 12 105 13
rect 107 17 115 25
rect 107 13 109 17
rect 113 13 115 17
rect 107 12 115 13
rect 117 25 125 26
rect 117 21 119 25
rect 123 21 125 25
rect 117 16 125 21
rect 127 21 134 26
rect 127 17 129 21
rect 133 17 134 21
rect 127 16 134 17
rect 117 12 122 16
rect 77 7 82 12
rect 40 3 53 4
<< pdiffusion >>
rect 70 68 76 69
rect 70 66 71 68
rect 4 59 9 66
rect 2 58 9 59
rect 2 54 3 58
rect 7 54 9 58
rect 2 51 9 54
rect 2 47 3 51
rect 7 47 9 51
rect 2 46 9 47
rect 4 38 9 46
rect 11 51 19 66
rect 11 47 13 51
rect 17 47 19 51
rect 11 43 19 47
rect 11 39 13 43
rect 17 39 19 43
rect 11 38 19 39
rect 21 58 29 66
rect 21 54 23 58
rect 27 54 29 58
rect 21 38 29 54
rect 31 43 39 66
rect 31 39 33 43
rect 37 39 39 43
rect 31 38 39 39
rect 41 58 49 66
rect 41 54 43 58
rect 47 54 49 58
rect 41 38 49 54
rect 51 43 59 66
rect 51 39 53 43
rect 57 39 59 43
rect 51 38 59 39
rect 61 38 66 66
rect 68 64 71 66
rect 75 64 76 68
rect 68 59 76 64
rect 106 68 113 69
rect 106 64 108 68
rect 112 66 113 68
rect 112 64 115 66
rect 106 59 115 64
rect 68 38 78 59
rect 80 38 85 59
rect 87 50 95 59
rect 87 46 89 50
rect 93 46 95 50
rect 87 43 95 46
rect 87 39 89 43
rect 93 39 95 43
rect 87 38 95 39
rect 97 38 102 59
rect 104 38 115 59
rect 117 57 122 66
rect 117 51 125 57
rect 117 47 119 51
rect 123 47 125 51
rect 117 44 125 47
rect 117 40 119 44
rect 123 40 125 44
rect 117 38 125 40
rect 127 56 134 57
rect 127 52 129 56
rect 133 52 134 56
rect 127 38 134 52
<< metal1 >>
rect -2 68 138 72
rect -2 64 71 68
rect 75 64 108 68
rect 112 64 128 68
rect 132 64 138 68
rect 2 54 3 58
rect 7 54 23 58
rect 27 54 43 58
rect 47 54 48 58
rect 54 55 123 59
rect 2 51 7 54
rect 54 51 58 55
rect 119 51 123 55
rect 129 56 133 64
rect 129 51 133 52
rect 2 47 3 51
rect 12 47 13 51
rect 17 47 58 51
rect 64 50 93 51
rect 64 47 89 50
rect 2 46 7 47
rect 2 18 6 46
rect 24 43 28 47
rect 64 43 68 47
rect 89 43 93 46
rect 119 44 123 47
rect 12 39 13 43
rect 17 39 28 43
rect 32 39 33 43
rect 37 39 53 43
rect 57 39 68 43
rect 24 34 28 39
rect 10 32 14 33
rect 24 30 26 34
rect 30 30 31 34
rect 10 26 14 28
rect 34 26 38 39
rect 74 34 78 43
rect 89 38 93 39
rect 106 35 110 43
rect 98 34 110 35
rect 49 30 56 34
rect 60 30 86 34
rect 90 30 91 34
rect 98 30 102 34
rect 106 30 110 34
rect 98 29 110 30
rect 10 25 103 26
rect 10 22 59 25
rect 58 21 59 22
rect 63 24 103 25
rect 63 22 79 24
rect 63 21 64 22
rect 83 22 99 24
rect 2 14 23 18
rect 27 14 69 18
rect 73 14 74 18
rect 79 17 83 20
rect 106 21 110 29
rect 114 40 119 43
rect 114 39 123 40
rect 114 25 118 39
rect 130 35 134 43
rect 122 34 134 35
rect 126 30 134 34
rect 122 29 134 30
rect 114 21 119 25
rect 123 21 124 25
rect 129 21 133 22
rect 99 17 103 20
rect 79 12 83 13
rect 88 13 89 17
rect 93 13 94 17
rect 88 8 94 13
rect 99 12 103 13
rect 108 13 109 17
rect 113 13 114 17
rect 108 8 114 13
rect 129 8 133 17
rect -2 4 5 8
rect 9 4 41 8
rect 45 4 48 8
rect 52 4 128 8
rect 132 4 138 8
rect -2 0 138 4
<< ntransistor >>
rect 12 12 14 24
rect 19 12 21 24
rect 29 12 31 24
rect 36 12 38 24
rect 55 11 57 26
rect 75 7 77 25
rect 85 12 87 25
rect 95 12 97 25
rect 105 12 107 25
rect 115 12 117 26
rect 125 16 127 26
<< ptransistor >>
rect 9 38 11 66
rect 19 38 21 66
rect 29 38 31 66
rect 39 38 41 66
rect 49 38 51 66
rect 59 38 61 66
rect 66 38 68 66
rect 78 38 80 59
rect 85 38 87 59
rect 95 38 97 59
rect 102 38 104 59
rect 115 38 117 66
rect 125 38 127 57
<< polycontact >>
rect 10 28 14 32
rect 26 30 30 34
rect 56 30 60 34
rect 86 30 90 34
rect 102 30 106 34
rect 122 30 126 34
<< ndcontact >>
rect 23 14 27 18
rect 5 4 9 8
rect 59 21 63 25
rect 69 14 73 18
rect 41 4 45 8
rect 48 4 52 8
rect 79 20 83 24
rect 79 13 83 17
rect 89 13 93 17
rect 99 20 103 24
rect 99 13 103 17
rect 109 13 113 17
rect 119 21 123 25
rect 129 17 133 21
<< pdcontact >>
rect 3 54 7 58
rect 3 47 7 51
rect 13 47 17 51
rect 13 39 17 43
rect 23 54 27 58
rect 33 39 37 43
rect 43 54 47 58
rect 53 39 57 43
rect 71 64 75 68
rect 108 64 112 68
rect 89 46 93 50
rect 89 39 93 43
rect 119 47 123 51
rect 119 40 123 44
rect 129 52 133 56
<< psubstratepcontact >>
rect 128 4 132 8
<< nsubstratencontact >>
rect 128 64 132 68
<< psubstratepdiff >>
rect 127 8 133 9
rect 127 4 128 8
rect 132 4 133 8
rect 127 3 133 4
<< nsubstratendiff >>
rect 127 68 133 69
rect 127 64 128 68
rect 132 64 133 68
rect 127 63 133 64
<< labels >>
rlabel ntransistor 13 18 13 18 6 an
rlabel polycontact 28 31 28 31 6 bn
rlabel metal1 12 16 12 16 6 z
rlabel metal1 20 16 20 16 6 z
rlabel metal1 12 27 12 27 6 an
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 56 12 56 6 z
rlabel metal1 20 56 20 56 6 z
rlabel metal1 36 16 36 16 6 z
rlabel metal1 44 16 44 16 6 z
rlabel metal1 28 16 28 16 6 z
rlabel polycontact 27 32 27 32 6 bn
rlabel metal1 20 41 20 41 6 bn
rlabel metal1 36 56 36 56 6 z
rlabel pdcontact 44 56 44 56 6 z
rlabel metal1 28 56 28 56 6 z
rlabel metal1 68 4 68 4 6 vss
rlabel metal1 60 16 60 16 6 z
rlabel metal1 68 16 68 16 6 z
rlabel metal1 52 16 52 16 6 z
rlabel metal1 60 32 60 32 6 a2
rlabel metal1 68 32 68 32 6 a2
rlabel metal1 52 32 52 32 6 a2
rlabel metal1 76 36 76 36 6 a2
rlabel metal1 50 41 50 41 6 an
rlabel metal1 35 49 35 49 6 bn
rlabel metal1 68 68 68 68 6 vdd
rlabel metal1 101 19 101 19 6 an
rlabel metal1 81 19 81 19 6 an
rlabel metal1 56 24 56 24 6 an
rlabel metal1 100 32 100 32 6 a1
rlabel metal1 108 32 108 32 6 a1
rlabel metal1 84 32 84 32 6 a2
rlabel metal1 91 44 91 44 6 an
rlabel metal1 119 23 119 23 6 bn
rlabel polycontact 124 32 124 32 6 b
rlabel metal1 132 36 132 36 6 b
rlabel pdcontact 121 49 121 49 6 bn
<< end >>
