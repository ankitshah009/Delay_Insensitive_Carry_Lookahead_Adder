magic
tech scmos
timestamp 1180600747
<< checkpaint >>
rect -22 -22 92 122
<< ab >>
rect 0 0 70 100
<< pwell >>
rect -4 -4 74 48
<< nwell >>
rect -4 48 74 104
<< polysilicon >>
rect 35 94 37 98
rect 47 94 49 98
rect 57 94 59 98
rect 11 84 13 88
rect 23 85 25 89
rect 11 43 13 55
rect 23 53 25 56
rect 35 53 37 56
rect 21 51 25 53
rect 33 51 37 53
rect 21 43 23 51
rect 33 43 35 51
rect 7 42 13 43
rect 7 38 8 42
rect 12 38 13 42
rect 7 37 13 38
rect 17 42 23 43
rect 17 38 18 42
rect 22 38 23 42
rect 17 37 23 38
rect 27 42 35 43
rect 27 38 28 42
rect 32 38 35 42
rect 47 43 49 55
rect 57 43 59 55
rect 47 42 53 43
rect 47 39 48 42
rect 27 37 35 38
rect 11 34 13 37
rect 21 34 23 37
rect 33 34 35 37
rect 45 38 48 39
rect 52 38 53 42
rect 45 37 53 38
rect 57 42 63 43
rect 57 38 58 42
rect 62 38 63 42
rect 57 37 63 38
rect 45 34 47 37
rect 57 34 59 37
rect 11 12 13 16
rect 21 13 23 17
rect 33 13 35 17
rect 45 13 47 17
rect 57 12 59 16
<< ndiffusion >>
rect 3 16 11 34
rect 13 17 21 34
rect 23 22 33 34
rect 23 18 26 22
rect 30 18 33 22
rect 23 17 33 18
rect 35 22 45 34
rect 35 18 38 22
rect 42 18 45 22
rect 35 17 45 18
rect 47 17 57 34
rect 13 16 18 17
rect 3 12 9 16
rect 49 16 57 17
rect 59 22 67 34
rect 59 18 62 22
rect 66 18 67 22
rect 59 16 67 18
rect 49 12 55 16
rect 3 8 4 12
rect 8 8 9 12
rect 3 7 9 8
rect 49 8 50 12
rect 54 8 55 12
rect 49 7 55 8
<< pdiffusion >>
rect 15 92 21 93
rect 15 88 16 92
rect 20 88 21 92
rect 15 85 21 88
rect 30 85 35 94
rect 15 84 23 85
rect 3 82 11 84
rect 3 78 4 82
rect 8 78 11 82
rect 3 55 11 78
rect 13 56 23 84
rect 25 82 35 85
rect 25 78 28 82
rect 32 78 35 82
rect 25 56 35 78
rect 37 72 47 94
rect 37 68 40 72
rect 44 68 47 72
rect 37 56 47 68
rect 13 55 18 56
rect 42 55 47 56
rect 49 55 57 94
rect 59 82 67 94
rect 59 78 62 82
rect 66 78 67 82
rect 59 55 67 78
<< metal1 >>
rect -2 92 72 100
rect -2 88 16 92
rect 20 88 72 92
rect 3 78 4 82
rect 8 78 28 82
rect 32 78 62 82
rect 66 78 67 82
rect 8 42 12 73
rect 8 17 12 38
rect 18 42 22 73
rect 18 27 22 38
rect 28 42 32 73
rect 28 37 32 38
rect 38 72 42 73
rect 38 68 40 72
rect 44 68 45 72
rect 28 32 32 33
rect 38 32 42 68
rect 28 28 42 32
rect 28 22 32 28
rect 38 27 42 28
rect 48 42 52 63
rect 48 27 52 38
rect 58 42 62 73
rect 58 27 62 38
rect 25 18 26 22
rect 30 18 32 22
rect 37 18 38 22
rect 42 18 62 22
rect 66 18 67 22
rect 28 17 32 18
rect -2 8 4 12
rect 8 10 50 12
rect 8 8 22 10
rect -2 6 22 8
rect 26 6 30 10
rect 34 6 38 10
rect 42 8 50 10
rect 54 8 72 12
rect 42 6 72 8
rect -2 0 72 6
<< ntransistor >>
rect 11 16 13 34
rect 21 17 23 34
rect 33 17 35 34
rect 45 17 47 34
rect 57 16 59 34
<< ptransistor >>
rect 11 55 13 84
rect 23 56 25 85
rect 35 56 37 94
rect 47 55 49 94
rect 57 55 59 94
<< polycontact >>
rect 8 38 12 42
rect 18 38 22 42
rect 28 38 32 42
rect 48 38 52 42
rect 58 38 62 42
<< ndcontact >>
rect 26 18 30 22
rect 38 18 42 22
rect 62 18 66 22
rect 4 8 8 12
rect 50 8 54 12
<< pdcontact >>
rect 16 88 20 92
rect 4 78 8 82
rect 28 78 32 82
rect 40 68 44 72
rect 62 78 66 82
<< psubstratepcontact >>
rect 22 6 26 10
rect 30 6 34 10
rect 38 6 42 10
<< psubstratepdiff >>
rect 21 10 43 11
rect 21 6 22 10
rect 26 6 30 10
rect 34 6 38 10
rect 42 6 43 10
rect 21 5 43 6
<< labels >>
rlabel metal1 10 45 10 45 6 i0
rlabel metal1 30 25 30 25 6 nq
rlabel metal1 20 50 20 50 6 i1
rlabel metal1 30 55 30 55 6 i4
rlabel metal1 35 6 35 6 6 vss
rlabel metal1 50 45 50 45 6 i2
rlabel metal1 40 50 40 50 6 nq
rlabel metal1 35 94 35 94 6 vdd
rlabel metal1 60 50 60 50 6 i3
<< end >>
