magic
tech scmos
timestamp 1179386267
<< checkpaint >>
rect -22 -22 118 94
<< ab >>
rect 0 0 96 72
<< pwell >>
rect -4 -4 100 32
<< nwell >>
rect -4 32 100 76
<< polysilicon >>
rect 9 62 11 67
rect 19 62 21 67
rect 29 62 31 67
rect 39 62 41 67
rect 49 62 51 67
rect 59 62 61 67
rect 69 62 71 67
rect 79 54 81 59
rect 9 35 11 38
rect 19 35 21 38
rect 29 35 31 38
rect 39 35 41 38
rect 49 35 51 38
rect 59 35 61 38
rect 69 35 71 38
rect 79 35 81 38
rect 9 34 15 35
rect 9 30 10 34
rect 14 30 15 34
rect 9 29 15 30
rect 19 34 33 35
rect 19 30 27 34
rect 31 30 33 34
rect 19 29 33 30
rect 12 26 14 29
rect 19 26 21 29
rect 31 26 33 29
rect 38 34 51 35
rect 38 30 39 34
rect 43 30 46 34
rect 50 30 51 34
rect 38 29 51 30
rect 55 34 62 35
rect 55 30 57 34
rect 61 30 62 34
rect 55 29 62 30
rect 66 34 81 35
rect 66 30 76 34
rect 80 30 81 34
rect 66 29 81 30
rect 38 26 40 29
rect 48 26 50 29
rect 55 26 57 29
rect 66 26 68 29
rect 12 2 14 6
rect 19 2 21 6
rect 31 2 33 6
rect 38 2 40 6
rect 48 2 50 6
rect 55 2 57 6
rect 66 2 68 6
<< ndiffusion >>
rect 5 25 12 26
rect 5 21 6 25
rect 10 21 12 25
rect 5 18 12 21
rect 5 14 6 18
rect 10 14 12 18
rect 5 13 12 14
rect 7 6 12 13
rect 14 6 19 26
rect 21 11 31 26
rect 21 7 24 11
rect 28 7 31 11
rect 21 6 31 7
rect 33 6 38 26
rect 40 25 48 26
rect 40 21 42 25
rect 46 21 48 25
rect 40 18 48 21
rect 40 14 42 18
rect 46 14 48 18
rect 40 6 48 14
rect 50 6 55 26
rect 57 18 66 26
rect 57 14 60 18
rect 64 14 66 18
rect 57 11 66 14
rect 57 7 60 11
rect 64 7 66 11
rect 57 6 66 7
rect 68 25 75 26
rect 68 21 70 25
rect 74 21 75 25
rect 68 18 75 21
rect 68 14 70 18
rect 74 14 75 18
rect 68 13 75 14
rect 68 6 73 13
<< pdiffusion >>
rect 2 61 9 62
rect 2 57 3 61
rect 7 57 9 61
rect 2 38 9 57
rect 11 58 19 62
rect 11 54 13 58
rect 17 54 19 58
rect 11 50 19 54
rect 11 46 13 50
rect 17 46 19 50
rect 11 38 19 46
rect 21 61 29 62
rect 21 57 23 61
rect 27 57 29 61
rect 21 38 29 57
rect 31 58 39 62
rect 31 54 33 58
rect 37 54 39 58
rect 31 50 39 54
rect 31 46 33 50
rect 37 46 39 50
rect 31 38 39 46
rect 41 61 49 62
rect 41 57 43 61
rect 47 57 49 61
rect 41 38 49 57
rect 51 58 59 62
rect 51 54 53 58
rect 57 54 59 58
rect 51 51 59 54
rect 51 47 53 51
rect 57 47 59 51
rect 51 38 59 47
rect 61 61 69 62
rect 61 57 63 61
rect 67 57 69 61
rect 61 53 69 57
rect 61 49 63 53
rect 67 49 69 53
rect 61 38 69 49
rect 71 54 76 62
rect 71 50 79 54
rect 71 46 73 50
rect 77 46 79 50
rect 71 43 79 46
rect 71 39 73 43
rect 77 39 79 43
rect 71 38 79 39
rect 81 53 89 54
rect 81 49 83 53
rect 87 49 89 53
rect 81 45 89 49
rect 81 41 83 45
rect 87 41 89 45
rect 81 38 89 41
<< metal1 >>
rect -2 68 98 72
rect -2 64 82 68
rect 86 64 98 68
rect 3 61 7 64
rect 23 61 27 64
rect 3 56 7 57
rect 13 58 17 59
rect 43 61 47 64
rect 23 56 27 57
rect 33 58 38 59
rect 13 51 17 54
rect 2 50 17 51
rect 37 54 38 58
rect 63 61 67 64
rect 43 56 47 57
rect 53 58 57 59
rect 33 50 38 54
rect 53 51 57 54
rect 2 46 13 50
rect 17 46 33 50
rect 37 47 53 50
rect 63 53 67 57
rect 83 53 87 64
rect 63 48 67 49
rect 73 50 77 51
rect 37 46 57 47
rect 2 21 6 46
rect 73 43 77 46
rect 17 35 23 42
rect 10 34 23 35
rect 14 30 23 34
rect 10 29 23 30
rect 27 39 73 42
rect 83 45 87 49
rect 83 40 87 41
rect 27 38 77 39
rect 27 34 31 38
rect 57 34 61 38
rect 27 29 31 30
rect 17 26 23 29
rect 35 26 39 34
rect 43 30 46 34
rect 50 30 51 34
rect 57 26 61 30
rect 74 34 86 35
rect 74 30 76 34
rect 80 30 86 34
rect 74 29 86 30
rect 10 21 11 25
rect 17 22 39 26
rect 42 25 47 26
rect 5 18 11 21
rect 46 21 47 25
rect 57 25 74 26
rect 57 22 70 25
rect 42 18 47 21
rect 70 18 74 21
rect 5 14 6 18
rect 10 14 42 18
rect 46 14 47 18
rect 59 14 60 18
rect 64 14 65 18
rect 59 11 65 14
rect 70 13 74 14
rect 82 13 86 29
rect 23 8 24 11
rect -2 7 24 8
rect 28 8 29 11
rect 59 8 60 11
rect 28 7 60 8
rect 64 8 65 11
rect 64 7 82 8
rect -2 4 82 7
rect 86 4 98 8
rect -2 0 98 4
<< ntransistor >>
rect 12 6 14 26
rect 19 6 21 26
rect 31 6 33 26
rect 38 6 40 26
rect 48 6 50 26
rect 55 6 57 26
rect 66 6 68 26
<< ptransistor >>
rect 9 38 11 62
rect 19 38 21 62
rect 29 38 31 62
rect 39 38 41 62
rect 49 38 51 62
rect 59 38 61 62
rect 69 38 71 62
rect 79 38 81 54
<< polycontact >>
rect 10 30 14 34
rect 27 30 31 34
rect 39 30 43 34
rect 46 30 50 34
rect 57 30 61 34
rect 76 30 80 34
<< ndcontact >>
rect 6 21 10 25
rect 6 14 10 18
rect 24 7 28 11
rect 42 21 46 25
rect 42 14 46 18
rect 60 14 64 18
rect 60 7 64 11
rect 70 21 74 25
rect 70 14 74 18
<< pdcontact >>
rect 3 57 7 61
rect 13 54 17 58
rect 13 46 17 50
rect 23 57 27 61
rect 33 54 37 58
rect 33 46 37 50
rect 43 57 47 61
rect 53 54 57 58
rect 53 47 57 51
rect 63 57 67 61
rect 63 49 67 53
rect 73 46 77 50
rect 73 39 77 43
rect 83 49 87 53
rect 83 41 87 45
<< psubstratepcontact >>
rect 82 4 86 8
<< nsubstratencontact >>
rect 82 64 86 68
<< psubstratepdiff >>
rect 80 8 88 24
rect 80 4 82 8
rect 86 4 88 8
rect 80 3 88 4
<< nsubstratendiff >>
rect 80 68 88 69
rect 80 64 82 68
rect 86 64 88 68
rect 80 61 88 64
<< labels >>
rlabel polycontact 58 32 58 32 6 an
rlabel metal1 12 16 12 16 6 z
rlabel polycontact 12 32 12 32 6 b
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 48 12 48 6 z
rlabel metal1 28 16 28 16 6 z
rlabel metal1 20 16 20 16 6 z
rlabel metal1 28 24 28 24 6 b
rlabel metal1 29 35 29 35 6 an
rlabel metal1 20 32 20 32 6 b
rlabel metal1 20 48 20 48 6 z
rlabel metal1 28 48 28 48 6 z
rlabel metal1 48 4 48 4 6 vss
rlabel ndcontact 44 16 44 16 6 z
rlabel metal1 36 16 36 16 6 z
rlabel metal1 36 24 36 24 6 b
rlabel metal1 44 32 44 32 6 b
rlabel metal1 36 52 36 52 6 z
rlabel metal1 44 48 44 48 6 z
rlabel metal1 52 48 52 48 6 z
rlabel metal1 48 68 48 68 6 vdd
rlabel metal1 72 19 72 19 6 an
rlabel metal1 76 32 76 32 6 a
rlabel polycontact 59 32 59 32 6 an
rlabel metal1 75 44 75 44 6 an
rlabel metal1 84 24 84 24 6 a
<< end >>
