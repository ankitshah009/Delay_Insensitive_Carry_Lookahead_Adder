.subckt nr2v0x05 a b vdd vss z
*   SPICE3 file   created from nr2v0x05.ext -      technology: scmos
m00 w1     b      z      vdd p w=20u  l=2.3636u ad=50p      pd=25u      as=112p     ps=54u
m01 vdd    a      w1     vdd p w=20u  l=2.3636u ad=180p     pd=58u      as=50p      ps=25u
m02 z      b      vss    vss n w=6u   l=2.3636u ad=24p      pd=14u      as=48p      ps=28u
m03 vss    a      z      vss n w=6u   l=2.3636u ad=48p      pd=28u      as=24p      ps=14u
C0  a      b      0.130f
C1  vdd    z      0.083f
C2  vss    a      0.044f
C3  vdd    b      0.031f
C4  z      b      0.132f
C5  vss    vdd    0.007f
C6  vdd    w1     0.005f
C7  vss    z      0.138f
C8  vdd    a      0.023f
C9  vss    b      0.011f
C10 z      a      0.054f
C11 w1     b      0.006f
C14 z      vss    0.018f
C15 a      vss    0.026f
C16 b      vss    0.021f
.ends
