magic
tech scmos
timestamp 1179386392
<< checkpaint >>
rect -22 -25 54 105
<< ab >>
rect 0 0 32 80
<< pwell >>
rect -4 -7 36 36
<< nwell >>
rect -4 36 36 87
<< polysilicon >>
rect 10 61 12 66
rect 20 61 22 65
rect 10 40 12 43
rect 9 39 15 40
rect 9 35 10 39
rect 14 35 15 39
rect 20 36 22 43
rect 9 34 15 35
rect 19 35 30 36
rect 12 27 14 34
rect 19 31 25 35
rect 29 31 30 35
rect 19 30 30 31
rect 19 27 21 30
rect 12 15 14 19
rect 19 14 21 19
<< ndiffusion >>
rect 5 26 12 27
rect 5 22 6 26
rect 10 22 12 26
rect 5 21 12 22
rect 7 19 12 21
rect 14 19 19 27
rect 21 20 30 27
rect 21 19 25 20
rect 23 16 25 19
rect 29 16 30 20
rect 23 15 30 16
<< pdiffusion >>
rect 2 62 8 63
rect 2 58 3 62
rect 7 61 8 62
rect 7 58 10 61
rect 2 43 10 58
rect 12 60 20 61
rect 12 56 14 60
rect 18 56 20 60
rect 12 53 20 56
rect 12 49 14 53
rect 18 49 20 53
rect 12 43 20 49
rect 22 60 30 61
rect 22 56 25 60
rect 29 56 30 60
rect 22 53 30 56
rect 22 49 25 53
rect 29 49 30 53
rect 22 43 30 49
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect -2 68 34 78
rect 2 62 8 68
rect 2 58 3 62
rect 7 58 8 62
rect 24 60 30 68
rect 13 56 14 60
rect 18 56 19 60
rect 13 54 19 56
rect 2 53 19 54
rect 2 49 14 53
rect 18 49 19 53
rect 24 56 25 60
rect 29 56 30 60
rect 24 53 30 56
rect 24 49 25 53
rect 29 49 30 53
rect 2 22 6 49
rect 17 43 23 46
rect 10 39 23 43
rect 10 33 14 35
rect 24 31 25 35
rect 29 31 30 35
rect 10 22 11 26
rect 18 25 30 31
rect 18 17 22 25
rect 25 20 29 21
rect 25 12 29 16
rect -2 2 34 12
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
<< ntransistor >>
rect 12 19 14 27
rect 19 19 21 27
<< ptransistor >>
rect 10 43 12 61
rect 20 43 22 61
<< polycontact >>
rect 10 35 14 39
rect 25 31 29 35
<< ndcontact >>
rect 6 22 10 26
rect 25 16 29 20
<< pdcontact >>
rect 3 58 7 62
rect 14 56 18 60
rect 14 49 18 53
rect 25 56 29 60
rect 25 49 29 53
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
<< psubstratepdiff >>
rect 0 2 32 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 32 2
rect 0 -3 32 -2
<< nsubstratendiff >>
rect 0 82 32 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 32 82
rect 0 77 32 78
<< labels >>
rlabel metal1 4 36 4 36 6 z
rlabel polycontact 12 36 12 36 6 b
rlabel metal1 12 52 12 52 6 z
rlabel metal1 16 6 16 6 6 vss
rlabel metal1 20 24 20 24 6 a
rlabel metal1 20 44 20 44 6 b
rlabel metal1 16 74 16 74 6 vdd
rlabel metal1 28 28 28 28 6 a
<< end >>
