magic
tech scmos
timestamp 1179385773
<< checkpaint >>
rect -22 -22 86 94
<< ab >>
rect 0 0 64 72
<< pwell >>
rect -4 -4 68 32
<< nwell >>
rect -4 32 68 76
<< polysilicon >>
rect 20 68 26 69
rect 20 64 21 68
rect 25 64 26 68
rect 20 63 26 64
rect 9 53 11 61
rect 9 43 11 46
rect 9 42 18 43
rect 9 41 13 42
rect 12 38 13 41
rect 17 38 18 42
rect 12 29 18 38
rect 22 41 26 63
rect 36 62 38 67
rect 43 62 45 67
rect 36 51 38 54
rect 43 51 45 54
rect 32 50 38 51
rect 32 46 33 50
rect 37 46 38 50
rect 32 45 38 46
rect 42 50 48 51
rect 42 46 43 50
rect 47 46 48 50
rect 42 45 48 46
rect 22 37 37 41
rect 9 27 18 29
rect 23 32 29 33
rect 23 28 24 32
rect 28 28 29 32
rect 23 27 29 28
rect 33 31 37 37
rect 33 27 49 31
rect 9 24 11 27
rect 16 24 18 27
rect 26 24 28 27
rect 33 24 35 27
rect 40 24 42 27
rect 47 24 49 27
rect 9 2 11 18
rect 16 2 18 18
rect 26 13 28 18
rect 33 13 35 18
rect 40 13 42 18
rect 47 13 49 18
<< ndiffusion >>
rect 2 23 9 24
rect 2 19 3 23
rect 7 19 9 23
rect 2 18 9 19
rect 11 18 16 24
rect 18 23 26 24
rect 18 19 20 23
rect 24 19 26 23
rect 18 18 26 19
rect 28 18 33 24
rect 35 18 40 24
rect 42 18 47 24
rect 49 23 56 24
rect 49 19 51 23
rect 55 19 56 23
rect 49 18 56 19
<< pdiffusion >>
rect 2 51 9 53
rect 2 47 3 51
rect 7 47 9 51
rect 2 46 9 47
rect 11 51 18 53
rect 11 47 13 51
rect 17 47 18 51
rect 11 46 18 47
rect 28 68 34 69
rect 28 64 29 68
rect 33 64 34 68
rect 28 62 34 64
rect 28 54 36 62
rect 38 54 43 62
rect 45 59 56 62
rect 45 55 51 59
rect 55 55 56 59
rect 45 54 56 55
<< metal1 >>
rect -2 68 66 72
rect -2 64 4 68
rect 8 64 12 68
rect 16 64 21 68
rect 25 64 29 68
rect 33 64 66 68
rect 2 51 8 59
rect 2 47 3 51
rect 7 47 8 51
rect 2 34 8 47
rect 12 51 18 64
rect 12 47 13 51
rect 17 47 18 51
rect 12 46 18 47
rect 22 55 51 59
rect 55 55 56 59
rect 22 42 28 55
rect 12 38 13 42
rect 17 38 28 42
rect 33 50 39 51
rect 37 46 39 50
rect 33 34 39 46
rect 2 28 19 34
rect 23 32 39 34
rect 23 28 24 32
rect 28 28 39 32
rect 43 50 47 51
rect 2 23 8 28
rect 2 19 3 23
rect 7 19 8 23
rect 2 13 8 19
rect 19 23 25 24
rect 19 19 20 23
rect 24 19 25 23
rect 19 8 25 19
rect 43 8 47 46
rect 50 23 56 55
rect 50 19 51 23
rect 55 19 56 23
rect 50 13 56 19
rect -2 4 42 8
rect 46 4 50 8
rect 54 4 66 8
rect -2 0 66 4
<< ntransistor >>
rect 9 18 11 24
rect 16 18 18 24
rect 26 18 28 24
rect 33 18 35 24
rect 40 18 42 24
rect 47 18 49 24
<< ptransistor >>
rect 9 46 11 53
rect 36 54 38 62
rect 43 54 45 62
<< polycontact >>
rect 21 64 25 68
rect 13 38 17 42
rect 33 46 37 50
rect 43 46 47 50
rect 24 28 28 32
<< ndcontact >>
rect 3 19 7 23
rect 20 19 24 23
rect 51 19 55 23
<< pdcontact >>
rect 3 47 7 51
rect 13 47 17 51
rect 29 64 33 68
rect 51 55 55 59
<< psubstratepcontact >>
rect 42 4 46 8
rect 50 4 54 8
<< nsubstratencontact >>
rect 4 64 8 68
rect 12 64 16 68
<< psubstratepdiff >>
rect 41 8 55 9
rect 41 4 42 8
rect 46 4 50 8
rect 54 4 55 8
rect 41 3 55 4
<< nsubstratendiff >>
rect 3 68 17 69
rect 3 64 4 68
rect 8 64 12 68
rect 16 64 17 68
rect 3 63 17 64
<< labels >>
rlabel polysilicon 15 35 15 35 6 an
rlabel metal1 12 32 12 32 6 z
rlabel metal1 4 36 4 36 6 z
rlabel metal1 28 32 28 32 6 a
rlabel metal1 20 40 20 40 6 an
rlabel metal1 32 4 32 4 6 vss
rlabel metal1 36 40 36 40 6 a
rlabel metal1 32 68 32 68 6 vdd
rlabel metal1 53 36 53 36 6 an
<< end >>
