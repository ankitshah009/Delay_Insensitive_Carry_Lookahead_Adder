magic
tech scmos
timestamp 1179387255
<< checkpaint >>
rect -22 -25 78 105
<< ab >>
rect 0 0 56 80
<< pwell >>
rect -4 -7 60 36
<< nwell >>
rect -4 36 60 87
<< polysilicon >>
rect 9 70 11 74
rect 22 70 24 74
rect 29 70 31 74
rect 36 70 38 74
rect 9 39 11 42
rect 22 39 24 42
rect 9 38 15 39
rect 9 34 10 38
rect 14 34 15 38
rect 9 33 15 34
rect 19 38 25 39
rect 19 34 20 38
rect 24 34 25 38
rect 19 33 25 34
rect 9 29 11 33
rect 19 23 21 33
rect 29 32 31 42
rect 36 39 38 42
rect 36 38 49 39
rect 36 37 44 38
rect 41 34 44 37
rect 48 34 49 38
rect 41 33 49 34
rect 29 31 37 32
rect 29 27 32 31
rect 36 27 37 31
rect 29 26 37 27
rect 29 23 31 26
rect 41 23 43 33
rect 9 10 11 15
rect 19 10 21 15
rect 29 10 31 15
rect 41 10 43 15
<< ndiffusion >>
rect 2 28 9 29
rect 2 24 3 28
rect 7 24 9 28
rect 2 23 9 24
rect 4 15 9 23
rect 11 23 16 29
rect 11 20 19 23
rect 11 16 13 20
rect 17 16 19 20
rect 11 15 19 16
rect 21 22 29 23
rect 21 18 23 22
rect 27 18 29 22
rect 21 15 29 18
rect 31 15 41 23
rect 43 22 50 23
rect 43 18 45 22
rect 49 18 50 22
rect 43 17 50 18
rect 43 15 48 17
rect 33 12 39 15
rect 33 8 34 12
rect 38 8 39 12
rect 33 7 39 8
<< pdiffusion >>
rect 13 72 20 73
rect 13 70 14 72
rect 4 64 9 70
rect 2 63 9 64
rect 2 59 3 63
rect 7 59 9 63
rect 2 56 9 59
rect 2 52 3 56
rect 7 52 9 56
rect 2 51 9 52
rect 4 42 9 51
rect 11 68 14 70
rect 18 70 20 72
rect 18 68 22 70
rect 11 42 22 68
rect 24 42 29 70
rect 31 42 36 70
rect 38 63 43 70
rect 38 62 45 63
rect 38 58 40 62
rect 44 58 45 62
rect 38 57 45 58
rect 38 42 43 57
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect -2 72 58 78
rect -2 68 14 72
rect 18 68 58 72
rect 2 59 3 63
rect 7 59 14 63
rect 2 57 14 59
rect 18 58 40 62
rect 44 58 45 62
rect 2 56 7 57
rect 2 52 3 56
rect 2 51 7 52
rect 2 29 6 51
rect 18 47 22 58
rect 34 49 46 55
rect 10 43 22 47
rect 10 38 14 43
rect 26 38 30 47
rect 17 34 20 38
rect 24 34 30 38
rect 10 29 14 34
rect 34 31 38 39
rect 42 38 46 49
rect 42 34 44 38
rect 48 34 49 38
rect 2 28 7 29
rect 2 24 3 28
rect 10 25 26 29
rect 31 27 32 31
rect 36 30 38 31
rect 36 27 47 30
rect 31 26 47 27
rect 2 23 7 24
rect 2 17 6 23
rect 22 22 26 25
rect 13 20 17 21
rect 22 18 23 22
rect 27 18 45 22
rect 49 18 50 22
rect 13 12 17 16
rect -2 8 34 12
rect 38 8 58 12
rect -2 2 58 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
<< ntransistor >>
rect 9 15 11 29
rect 19 15 21 23
rect 29 15 31 23
rect 41 15 43 23
<< ptransistor >>
rect 9 42 11 70
rect 22 42 24 70
rect 29 42 31 70
rect 36 42 38 70
<< polycontact >>
rect 10 34 14 38
rect 20 34 24 38
rect 44 34 48 38
rect 32 27 36 31
<< ndcontact >>
rect 3 24 7 28
rect 13 16 17 20
rect 23 18 27 22
rect 45 18 49 22
rect 34 8 38 12
<< pdcontact >>
rect 3 59 7 63
rect 3 52 7 56
rect 14 68 18 72
rect 40 58 44 62
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
<< psubstratepdiff >>
rect 0 2 56 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 56 2
rect 0 -3 56 -2
<< nsubstratendiff >>
rect 0 82 56 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 56 82
rect 0 77 56 78
<< labels >>
rlabel polycontact 12 36 12 36 6 zn
rlabel metal1 4 40 4 40 6 z
rlabel metal1 20 36 20 36 6 a
rlabel polycontact 12 36 12 36 6 zn
rlabel metal1 12 60 12 60 6 z
rlabel metal1 28 6 28 6 6 vss
rlabel metal1 36 32 36 32 6 b
rlabel metal1 28 44 28 44 6 a
rlabel metal1 36 52 36 52 6 c
rlabel metal1 28 74 28 74 6 vdd
rlabel metal1 36 20 36 20 6 zn
rlabel metal1 44 28 44 28 6 b
rlabel metal1 44 48 44 48 6 c
rlabel metal1 31 60 31 60 6 zn
<< end >>
