magic
tech scmos
timestamp 1179385830
<< checkpaint >>
rect -22 -25 54 105
<< ab >>
rect 0 0 32 80
<< pwell >>
rect -4 -7 36 36
<< nwell >>
rect -4 36 36 87
<< polysilicon >>
rect 10 69 12 73
rect 20 61 22 65
rect 10 40 12 45
rect 20 40 22 45
rect 10 39 30 40
rect 10 38 25 39
rect 10 30 12 38
rect 20 35 25 38
rect 29 35 30 39
rect 20 34 30 35
rect 20 30 22 34
rect 10 15 12 20
rect 20 15 22 20
<< ndiffusion >>
rect 2 22 10 30
rect 2 18 3 22
rect 7 20 10 22
rect 12 29 20 30
rect 12 25 14 29
rect 18 25 20 29
rect 12 20 20 25
rect 22 25 30 30
rect 22 21 25 25
rect 29 21 30 25
rect 22 20 30 21
rect 7 18 8 20
rect 2 17 8 18
<< pdiffusion >>
rect 2 68 10 69
rect 2 64 4 68
rect 8 64 10 68
rect 2 61 10 64
rect 2 57 4 61
rect 8 57 10 61
rect 2 45 10 57
rect 12 61 17 69
rect 12 54 20 61
rect 12 50 14 54
rect 18 50 20 54
rect 12 45 20 50
rect 22 60 30 61
rect 22 56 24 60
rect 28 56 30 60
rect 22 53 30 56
rect 22 49 24 53
rect 28 49 30 53
rect 22 45 30 49
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect -2 68 34 78
rect 3 64 4 68
rect 8 64 9 68
rect 3 61 9 64
rect 3 57 4 61
rect 8 57 9 61
rect 23 60 29 68
rect 23 56 24 60
rect 28 56 29 60
rect 2 50 14 54
rect 18 50 19 54
rect 23 53 29 56
rect 2 31 6 50
rect 23 49 24 53
rect 28 49 29 53
rect 17 42 30 46
rect 24 39 30 42
rect 24 35 25 39
rect 29 35 30 39
rect 26 33 30 35
rect 2 29 22 31
rect 2 25 14 29
rect 18 25 22 29
rect 25 25 29 26
rect 2 18 3 22
rect 7 18 8 22
rect 2 12 8 18
rect 25 12 29 21
rect -2 2 34 12
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
<< ntransistor >>
rect 10 20 12 30
rect 20 20 22 30
<< ptransistor >>
rect 10 45 12 69
rect 20 45 22 61
<< polycontact >>
rect 25 35 29 39
<< ndcontact >>
rect 3 18 7 22
rect 14 25 18 29
rect 25 21 29 25
<< pdcontact >>
rect 4 64 8 68
rect 4 57 8 61
rect 14 50 18 54
rect 24 56 28 60
rect 24 49 28 53
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
<< psubstratepdiff >>
rect 0 2 32 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 32 2
rect 0 -3 32 -2
<< nsubstratendiff >>
rect 0 82 32 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 32 82
rect 0 77 32 78
<< labels >>
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 28 12 28 6 z
rlabel metal1 12 52 12 52 6 z
rlabel metal1 16 6 16 6 6 vss
rlabel metal1 20 28 20 28 6 z
rlabel metal1 20 44 20 44 6 a
rlabel metal1 16 74 16 74 6 vdd
rlabel polycontact 28 36 28 36 6 a
<< end >>
