magic
tech scmos
timestamp 1179387745
<< checkpaint >>
rect -22 -25 94 105
<< ab >>
rect 0 0 72 80
<< pwell >>
rect -4 -7 76 36
<< nwell >>
rect -4 36 76 87
<< polysilicon >>
rect 25 70 27 74
rect 32 70 34 74
rect 42 70 44 74
rect 52 70 54 74
rect 2 62 8 63
rect 2 58 3 62
rect 7 59 8 62
rect 7 58 11 59
rect 2 57 11 58
rect 9 54 11 57
rect 61 54 63 58
rect 9 40 11 43
rect 25 40 27 43
rect 9 38 27 40
rect 32 39 34 43
rect 42 39 44 43
rect 52 40 54 43
rect 61 40 63 43
rect 32 38 38 39
rect 9 30 11 38
rect 19 30 21 38
rect 32 34 33 38
rect 37 34 38 38
rect 26 30 28 34
rect 32 33 38 34
rect 42 38 48 39
rect 52 38 63 40
rect 42 34 43 38
rect 47 34 48 38
rect 42 33 48 34
rect 36 30 38 33
rect 43 30 45 33
rect 54 30 56 38
rect 9 19 11 24
rect 54 18 56 24
rect 64 21 70 22
rect 64 18 65 21
rect 19 13 21 18
rect 26 10 28 18
rect 36 14 38 18
rect 43 14 45 18
rect 54 17 65 18
rect 69 17 70 21
rect 54 16 70 17
rect 54 10 56 16
rect 26 8 56 10
<< ndiffusion >>
rect 2 29 9 30
rect 2 25 3 29
rect 7 25 9 29
rect 2 24 9 25
rect 11 29 19 30
rect 11 25 13 29
rect 17 25 19 29
rect 11 24 19 25
rect 13 18 19 24
rect 21 18 26 30
rect 28 23 36 30
rect 28 19 30 23
rect 34 19 36 23
rect 28 18 36 19
rect 38 18 43 30
rect 45 24 54 30
rect 56 29 63 30
rect 56 25 58 29
rect 62 25 63 29
rect 56 24 63 25
rect 45 23 52 24
rect 45 19 47 23
rect 51 19 52 23
rect 45 18 52 19
<< pdiffusion >>
rect 13 65 25 70
rect 13 61 19 65
rect 23 61 25 65
rect 13 54 25 61
rect 4 49 9 54
rect 2 48 9 49
rect 2 44 3 48
rect 7 44 9 48
rect 2 43 9 44
rect 11 43 25 54
rect 27 43 32 70
rect 34 48 42 70
rect 34 44 36 48
rect 40 44 42 48
rect 34 43 42 44
rect 44 43 52 70
rect 54 65 61 70
rect 54 61 56 65
rect 60 61 61 65
rect 54 60 61 61
rect 54 54 59 60
rect 54 43 61 54
rect 63 49 68 54
rect 63 48 70 49
rect 63 44 65 48
rect 69 44 70 48
rect 63 43 70 44
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect -2 68 74 78
rect 19 65 23 68
rect 2 62 7 63
rect 2 58 3 62
rect 19 60 23 61
rect 56 65 60 68
rect 56 60 60 61
rect 2 54 14 58
rect 10 49 14 54
rect 18 52 49 56
rect 3 48 7 49
rect 18 45 22 52
rect 35 46 36 48
rect 7 44 22 45
rect 3 41 22 44
rect 26 44 36 46
rect 40 44 41 48
rect 26 42 41 44
rect 3 29 7 41
rect 3 24 7 25
rect 13 29 17 30
rect 13 12 17 25
rect 26 19 30 42
rect 33 38 38 39
rect 45 38 49 52
rect 37 34 38 38
rect 42 34 43 38
rect 47 34 49 38
rect 59 44 65 48
rect 69 44 70 48
rect 33 33 38 34
rect 34 31 38 33
rect 59 31 63 44
rect 34 29 63 31
rect 34 27 58 29
rect 57 25 58 27
rect 62 25 63 29
rect 34 19 35 23
rect 46 19 47 23
rect 51 19 52 23
rect 66 22 70 31
rect 46 12 52 19
rect 57 21 70 22
rect 57 17 65 21
rect 69 17 70 21
rect -2 2 74 12
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
<< ntransistor >>
rect 9 24 11 30
rect 19 18 21 30
rect 26 18 28 30
rect 36 18 38 30
rect 43 18 45 30
rect 54 24 56 30
<< ptransistor >>
rect 9 43 11 54
rect 25 43 27 70
rect 32 43 34 70
rect 42 43 44 70
rect 52 43 54 70
rect 61 43 63 54
<< polycontact >>
rect 3 58 7 62
rect 33 34 37 38
rect 43 34 47 38
rect 65 17 69 21
<< ndcontact >>
rect 3 25 7 29
rect 13 25 17 29
rect 30 19 34 23
rect 58 25 62 29
rect 47 19 51 23
<< pdcontact >>
rect 19 61 23 65
rect 3 44 7 48
rect 36 44 40 48
rect 56 61 60 65
rect 65 44 69 48
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
<< psubstratepdiff >>
rect 0 2 72 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 72 2
rect 0 -3 72 -2
<< nsubstratendiff >>
rect 0 82 72 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 72 82
rect 0 77 72 78
<< labels >>
rlabel polycontact 35 36 35 36 6 bn
rlabel polycontact 45 36 45 36 6 an
rlabel metal1 5 36 5 36 6 an
rlabel polycontact 4 60 4 60 6 a
rlabel metal1 12 52 12 52 6 a
rlabel metal1 36 6 36 6 6 vss
rlabel metal1 36 33 36 33 6 bn
rlabel metal1 28 32 28 32 6 z
rlabel metal1 36 44 36 44 6 z
rlabel metal1 36 74 36 74 6 vdd
rlabel metal1 47 45 47 45 6 an
rlabel metal1 60 20 60 20 6 b
rlabel metal1 68 24 68 24 6 b
rlabel metal1 64 46 64 46 6 bn
rlabel metal1 61 36 61 36 6 bn
<< end >>
