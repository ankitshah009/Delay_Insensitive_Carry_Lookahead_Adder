magic
tech scmos
timestamp 1179386656
<< checkpaint >>
rect -22 -25 102 105
<< ab >>
rect 0 0 80 80
<< pwell >>
rect -4 -7 84 36
<< nwell >>
rect -4 36 84 87
<< polysilicon >>
rect 9 69 11 74
rect 19 69 21 74
rect 32 69 34 74
rect 42 69 44 74
rect 64 54 70 55
rect 64 50 65 54
rect 69 50 70 54
rect 64 49 70 50
rect 54 46 60 47
rect 9 35 11 44
rect 19 41 21 44
rect 32 41 34 44
rect 19 40 25 41
rect 19 36 20 40
rect 24 36 25 40
rect 32 40 38 41
rect 32 37 33 40
rect 19 35 25 36
rect 29 36 33 37
rect 37 36 38 40
rect 29 35 38 36
rect 42 39 44 44
rect 54 42 55 46
rect 59 42 60 46
rect 54 41 60 42
rect 42 38 49 39
rect 9 34 15 35
rect 9 30 10 34
rect 14 31 15 34
rect 14 30 17 31
rect 9 29 17 30
rect 15 26 17 29
rect 22 26 24 35
rect 29 26 31 35
rect 42 34 44 38
rect 48 34 49 38
rect 42 33 49 34
rect 42 31 48 33
rect 54 32 56 41
rect 64 37 66 49
rect 36 29 48 31
rect 36 26 38 29
rect 46 26 48 29
rect 53 29 56 32
rect 60 35 66 37
rect 53 26 55 29
rect 60 26 62 35
rect 72 34 78 35
rect 72 31 73 34
rect 67 30 73 31
rect 77 30 78 34
rect 67 29 78 30
rect 67 26 69 29
rect 15 6 17 11
rect 22 6 24 11
rect 29 6 31 11
rect 36 6 38 11
rect 46 6 48 11
rect 53 6 55 11
rect 60 6 62 11
rect 67 6 69 11
<< ndiffusion >>
rect 6 12 15 26
rect 6 8 8 12
rect 12 11 15 12
rect 17 11 22 26
rect 24 11 29 26
rect 31 11 36 26
rect 38 22 46 26
rect 38 18 40 22
rect 44 18 46 22
rect 38 11 46 18
rect 48 11 53 26
rect 55 11 60 26
rect 62 11 67 26
rect 69 16 77 26
rect 69 12 71 16
rect 75 12 77 16
rect 69 11 77 12
rect 12 8 13 11
rect 6 7 13 8
<< pdiffusion >>
rect 24 69 30 71
rect 2 68 9 69
rect 2 64 3 68
rect 7 64 9 68
rect 2 61 9 64
rect 2 57 3 61
rect 7 57 9 61
rect 2 44 9 57
rect 11 62 19 69
rect 11 58 13 62
rect 17 58 19 62
rect 11 54 19 58
rect 11 50 13 54
rect 17 50 19 54
rect 11 44 19 50
rect 21 65 25 69
rect 29 65 32 69
rect 21 44 32 65
rect 34 62 42 69
rect 34 58 36 62
rect 40 58 42 62
rect 34 44 42 58
rect 44 68 52 69
rect 44 64 46 68
rect 50 64 52 68
rect 44 61 52 64
rect 44 57 46 61
rect 50 57 52 61
rect 44 44 52 57
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect -2 69 82 78
rect -2 68 25 69
rect 2 64 3 68
rect 7 64 8 68
rect 24 65 25 68
rect 29 68 82 69
rect 29 65 30 68
rect 2 61 8 64
rect 45 64 46 68
rect 50 64 51 68
rect 2 57 3 61
rect 7 57 8 61
rect 12 58 13 62
rect 17 58 36 62
rect 40 58 41 62
rect 45 61 51 64
rect 12 54 18 58
rect 45 57 46 61
rect 50 57 51 61
rect 58 54 62 63
rect 2 50 13 54
rect 17 50 18 54
rect 24 50 65 54
rect 69 50 71 54
rect 2 22 6 50
rect 24 46 28 50
rect 17 42 28 46
rect 33 42 55 46
rect 59 42 60 46
rect 64 42 71 46
rect 20 40 24 42
rect 20 35 24 36
rect 33 40 39 42
rect 37 36 39 40
rect 64 38 68 42
rect 10 34 14 35
rect 33 34 39 36
rect 43 34 44 38
rect 48 34 68 38
rect 72 34 78 35
rect 72 30 73 34
rect 77 30 78 34
rect 10 26 78 30
rect 58 25 78 26
rect 2 18 40 22
rect 44 18 47 22
rect 58 17 62 25
rect 71 16 75 17
rect -2 8 8 12
rect 12 8 82 12
rect -2 2 82 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
<< ntransistor >>
rect 15 11 17 26
rect 22 11 24 26
rect 29 11 31 26
rect 36 11 38 26
rect 46 11 48 26
rect 53 11 55 26
rect 60 11 62 26
rect 67 11 69 26
<< ptransistor >>
rect 9 44 11 69
rect 19 44 21 69
rect 32 44 34 69
rect 42 44 44 69
<< polycontact >>
rect 65 50 69 54
rect 20 36 24 40
rect 33 36 37 40
rect 55 42 59 46
rect 10 30 14 34
rect 44 34 48 38
rect 73 30 77 34
<< ndcontact >>
rect 8 8 12 12
rect 40 18 44 22
rect 71 12 75 16
<< pdcontact >>
rect 3 64 7 68
rect 3 57 7 61
rect 13 58 17 62
rect 13 50 17 54
rect 25 65 29 69
rect 36 58 40 62
rect 46 64 50 68
rect 46 57 50 61
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
<< psubstratepdiff >>
rect 0 2 80 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 80 2
rect 0 -3 80 -2
<< nsubstratendiff >>
rect 0 82 80 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 80 82
rect 0 77 80 78
<< labels >>
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 20 12 20 6 z
rlabel metal1 20 20 20 20 6 z
rlabel metal1 20 28 20 28 6 a
rlabel metal1 28 20 28 20 6 z
rlabel metal1 28 28 28 28 6 a
rlabel metal1 20 44 20 44 6 b
rlabel metal1 28 52 28 52 6 b
rlabel metal1 12 52 12 52 6 z
rlabel metal1 20 60 20 60 6 z
rlabel metal1 28 60 28 60 6 z
rlabel metal1 40 6 40 6 6 vss
rlabel metal1 36 20 36 20 6 z
rlabel metal1 36 28 36 28 6 a
rlabel metal1 44 20 44 20 6 z
rlabel metal1 44 28 44 28 6 a
rlabel metal1 36 40 36 40 6 c
rlabel metal1 44 44 44 44 6 c
rlabel metal1 36 52 36 52 6 b
rlabel metal1 44 52 44 52 6 b
rlabel metal1 36 60 36 60 6 z
rlabel metal1 40 74 40 74 6 vdd
rlabel metal1 52 28 52 28 6 a
rlabel metal1 60 24 60 24 6 a
rlabel metal1 52 36 52 36 6 d
rlabel metal1 52 44 52 44 6 c
rlabel metal1 60 36 60 36 6 d
rlabel metal1 52 52 52 52 6 b
rlabel metal1 60 56 60 56 6 b
rlabel metal1 68 28 68 28 6 a
rlabel metal1 76 28 76 28 6 a
rlabel metal1 68 44 68 44 6 d
rlabel polycontact 68 52 68 52 6 b
<< end >>
