magic
tech scmos
timestamp 1171447624
<< checkpaint >>
rect -22 -26 118 114
<< ab >>
rect 0 0 96 88
<< pwell >>
rect -4 -8 100 40
<< nwell >>
rect -4 40 100 96
<< polysilicon >>
rect 2 77 11 83
rect 9 74 11 77
rect 21 77 30 83
rect 34 77 43 83
rect 21 74 23 77
rect 41 74 43 77
rect 53 77 62 83
rect 66 77 75 83
rect 53 74 55 77
rect 73 74 75 77
rect 85 82 94 83
rect 85 78 86 82
rect 90 78 94 82
rect 85 77 94 78
rect 85 74 87 77
rect 9 43 11 46
rect 21 43 23 46
rect 41 43 43 46
rect 53 43 55 46
rect 73 43 75 46
rect 85 43 87 46
rect 2 42 14 43
rect 2 38 6 42
rect 10 38 14 42
rect 2 37 14 38
rect 18 42 30 43
rect 18 38 22 42
rect 26 38 30 42
rect 18 37 30 38
rect 34 42 46 43
rect 34 38 38 42
rect 42 38 46 42
rect 34 37 46 38
rect 50 42 62 43
rect 50 38 54 42
rect 58 38 62 42
rect 50 37 62 38
rect 66 42 78 43
rect 66 38 70 42
rect 74 38 78 42
rect 66 37 78 38
rect 82 37 94 43
rect 9 34 11 37
rect 21 34 23 37
rect 41 34 43 37
rect 53 34 55 37
rect 73 34 75 37
rect 85 34 87 37
rect 9 11 11 14
rect 2 5 11 11
rect 21 11 23 14
rect 41 11 43 14
rect 21 5 30 11
rect 34 5 43 11
rect 53 11 55 14
rect 73 11 75 14
rect 53 5 62 11
rect 66 5 75 11
rect 85 11 87 14
rect 85 5 94 11
<< ndiffusion >>
rect 2 28 9 34
rect 2 24 3 28
rect 7 24 9 28
rect 2 21 9 24
rect 2 17 3 21
rect 7 17 9 21
rect 2 14 9 17
rect 11 15 21 34
rect 11 14 14 15
rect 13 11 14 14
rect 18 14 21 15
rect 23 30 30 34
rect 23 26 25 30
rect 29 26 30 30
rect 23 14 30 26
rect 34 29 41 34
rect 34 25 35 29
rect 39 25 41 29
rect 34 22 41 25
rect 34 18 35 22
rect 39 18 41 22
rect 34 14 41 18
rect 43 33 53 34
rect 43 29 46 33
rect 50 29 53 33
rect 43 14 53 29
rect 55 19 62 34
rect 55 15 57 19
rect 61 15 62 19
rect 55 14 62 15
rect 66 33 73 34
rect 66 29 67 33
rect 71 29 73 33
rect 66 26 73 29
rect 66 22 67 26
rect 71 22 73 26
rect 66 14 73 22
rect 75 26 85 34
rect 75 22 78 26
rect 82 22 85 26
rect 75 18 85 22
rect 75 14 78 18
rect 82 14 85 18
rect 87 14 94 34
rect 18 11 19 14
rect 13 6 19 11
rect 13 3 14 6
rect 18 3 19 6
rect 13 2 19 3
rect 45 2 51 14
rect 77 2 83 14
<< pdiffusion >>
rect 13 85 19 86
rect 13 82 14 85
rect 18 82 19 85
rect 13 77 19 82
rect 13 74 14 77
rect 2 69 9 74
rect 2 65 3 69
rect 7 65 9 69
rect 2 62 9 65
rect 2 58 3 62
rect 7 58 9 62
rect 2 46 9 58
rect 11 73 14 74
rect 18 74 19 77
rect 45 74 51 86
rect 77 74 83 86
rect 18 73 21 74
rect 11 46 21 73
rect 23 62 30 74
rect 23 58 25 62
rect 29 58 30 62
rect 23 46 30 58
rect 34 73 41 74
rect 34 69 35 73
rect 39 69 41 73
rect 34 46 41 69
rect 43 51 53 74
rect 43 47 46 51
rect 50 47 53 51
rect 43 46 53 47
rect 55 73 62 74
rect 55 69 57 73
rect 61 69 62 73
rect 55 66 62 69
rect 55 62 57 66
rect 61 62 62 66
rect 55 46 62 62
rect 66 66 73 74
rect 66 62 67 66
rect 71 62 73 66
rect 66 59 73 62
rect 66 55 67 59
rect 71 55 73 59
rect 66 46 73 55
rect 75 70 78 74
rect 82 70 85 74
rect 75 67 85 70
rect 75 63 78 67
rect 82 63 85 67
rect 75 46 85 63
rect 87 46 94 74
<< metal1 >>
rect -2 86 2 90
rect 10 86 22 90
rect 30 86 34 90
rect 42 86 54 90
rect 62 86 66 90
rect 74 86 86 90
rect 94 86 98 90
rect 14 85 18 86
rect 14 77 18 78
rect 78 82 82 86
rect 78 74 82 78
rect 86 82 90 86
rect 86 77 90 78
rect 14 72 18 73
rect 22 69 35 73
rect 39 69 40 73
rect 56 69 57 73
rect 61 69 62 73
rect 2 65 3 69
rect 7 65 26 69
rect 56 66 62 69
rect 78 67 82 70
rect 2 62 8 65
rect 2 58 3 62
rect 7 58 8 62
rect 6 42 10 55
rect 6 33 10 38
rect 14 29 18 65
rect 30 62 57 66
rect 61 62 62 66
rect 67 66 71 67
rect 78 62 82 63
rect 24 58 25 62
rect 29 58 34 62
rect 67 59 71 62
rect 22 42 26 55
rect 22 33 26 38
rect 30 30 34 58
rect 38 55 67 59
rect 71 55 82 59
rect 38 42 42 55
rect 38 37 42 38
rect 46 51 50 52
rect 46 33 50 47
rect 3 28 18 29
rect 7 25 18 28
rect 24 26 25 30
rect 29 29 39 30
rect 29 26 35 29
rect 3 21 7 24
rect 14 23 18 25
rect 14 19 26 23
rect 3 16 7 17
rect 14 15 18 16
rect 14 10 18 11
rect 22 13 26 19
rect 35 22 39 25
rect 35 17 39 18
rect 46 17 50 29
rect 54 42 74 47
rect 54 25 58 38
rect 70 37 74 38
rect 78 34 82 55
rect 67 33 82 34
rect 71 30 82 33
rect 67 26 71 29
rect 67 21 71 22
rect 78 26 82 27
rect 57 19 61 20
rect 57 13 61 15
rect 22 9 61 13
rect 78 18 82 22
rect 78 10 82 14
rect 14 2 18 3
rect 78 2 82 6
rect -2 -2 2 2
rect 10 -2 22 2
rect 30 -2 34 2
rect 42 -2 54 2
rect 62 -2 66 2
rect 74 -2 86 2
rect 94 -2 98 2
<< metal2 >>
rect -2 86 6 90
rect 10 86 22 90
rect 26 86 38 90
rect 42 86 54 90
rect 58 86 70 90
rect 74 86 86 90
rect 90 86 98 90
rect -2 82 98 86
rect -2 78 14 82
rect 18 78 78 82
rect 82 78 98 82
rect -2 76 98 78
rect -2 10 98 12
rect -2 6 14 10
rect 18 6 78 10
rect 82 6 98 10
rect -2 2 98 6
rect -2 -2 6 2
rect 10 -2 22 2
rect 26 -2 38 2
rect 42 -2 54 2
rect 58 -2 70 2
rect 74 -2 86 2
rect 90 -2 98 2
<< ntransistor >>
rect 9 14 11 34
rect 21 14 23 34
rect 41 14 43 34
rect 53 14 55 34
rect 73 14 75 34
rect 85 14 87 34
<< ptransistor >>
rect 9 46 11 74
rect 21 46 23 74
rect 41 46 43 74
rect 53 46 55 74
rect 73 46 75 74
rect 85 46 87 74
<< polycontact >>
rect 86 78 90 82
rect 6 38 10 42
rect 22 38 26 42
rect 38 38 42 42
rect 54 38 58 42
rect 70 38 74 42
<< ndcontact >>
rect 3 24 7 28
rect 3 17 7 21
rect 14 11 18 15
rect 25 26 29 30
rect 35 25 39 29
rect 35 18 39 22
rect 46 29 50 33
rect 57 15 61 19
rect 67 29 71 33
rect 67 22 71 26
rect 78 22 82 26
rect 78 14 82 18
rect 14 3 18 6
<< pdcontact >>
rect 14 82 18 85
rect 3 65 7 69
rect 3 58 7 62
rect 14 73 18 77
rect 25 58 29 62
rect 35 69 39 73
rect 46 47 50 51
rect 57 69 61 73
rect 57 62 61 66
rect 67 62 71 66
rect 67 55 71 59
rect 78 70 82 74
rect 78 63 82 67
<< m2contact >>
rect 6 86 10 90
rect 22 86 26 90
rect 38 86 42 90
rect 54 86 58 90
rect 70 86 74 90
rect 86 86 90 90
rect 14 78 18 82
rect 78 78 82 82
rect 14 6 18 10
rect 78 6 82 10
rect 6 -2 10 2
rect 22 -2 26 2
rect 38 -2 42 2
rect 54 -2 58 2
rect 70 -2 74 2
rect 86 -2 90 2
<< psubstratepcontact >>
rect 2 -2 6 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 90 -2 94 2
<< nsubstratencontact >>
rect 2 86 6 90
rect 26 86 30 90
rect 34 86 38 90
rect 58 86 62 90
rect 66 86 70 90
rect 90 86 94 90
<< psubstratepdiff >>
rect 0 2 7 3
rect 25 2 39 3
rect 57 2 71 3
rect 89 2 96 3
rect 0 -2 2 2
rect 6 -2 7 2
rect 0 -3 7 -2
rect 25 -2 26 2
rect 30 -2 34 2
rect 38 -2 39 2
rect 25 -3 39 -2
rect 57 -2 58 2
rect 62 -2 66 2
rect 70 -2 71 2
rect 57 -3 71 -2
rect 89 -2 90 2
rect 94 -2 96 2
rect 89 -3 96 -2
<< nsubstratendiff >>
rect 0 90 7 91
rect 0 86 2 90
rect 6 86 7 90
rect 25 90 39 91
rect 25 86 26 90
rect 30 86 34 90
rect 38 86 39 90
rect 57 90 71 91
rect 57 86 58 90
rect 62 86 66 90
rect 70 86 71 90
rect 89 90 96 91
rect 89 86 90 90
rect 94 86 96 90
rect 0 85 7 86
rect 25 85 39 86
rect 57 85 71 86
rect 89 85 96 86
<< labels >>
rlabel metal1 8 44 8 44 6 a1
rlabel metal1 24 44 24 44 6 a0
rlabel ndcontact 48 32 48 32 6 z
rlabel metal1 56 36 56 36 6 s
rlabel metal1 64 44 64 44 6 s
rlabel metal1 72 44 72 44 6 s
rlabel metal2 48 6 48 6 6 vss
rlabel metal2 48 82 48 82 6 vdd
<< end >>
