magic
tech scmos
timestamp 1179386261
<< checkpaint >>
rect -22 -25 86 105
<< ab >>
rect 0 0 64 80
<< pwell >>
rect -4 -7 68 36
<< nwell >>
rect -4 36 68 87
<< polysilicon >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 39 70 41 74
rect 49 70 51 74
rect 9 39 11 46
rect 19 39 21 46
rect 29 39 31 46
rect 39 39 41 46
rect 49 40 51 43
rect 9 38 15 39
rect 9 34 10 38
rect 14 34 15 38
rect 9 33 15 34
rect 19 38 31 39
rect 19 34 26 38
rect 30 34 31 38
rect 19 33 31 34
rect 35 38 41 39
rect 35 34 36 38
rect 40 34 41 38
rect 45 39 51 40
rect 45 35 46 39
rect 50 35 51 39
rect 45 34 51 35
rect 35 33 41 34
rect 12 30 14 33
rect 19 30 21 33
rect 29 30 31 33
rect 36 30 38 33
rect 47 30 49 34
rect 47 11 49 16
rect 12 6 14 10
rect 19 6 21 10
rect 29 6 31 10
rect 36 6 38 10
<< ndiffusion >>
rect 4 15 12 30
rect 4 11 6 15
rect 10 11 12 15
rect 4 10 12 11
rect 14 10 19 30
rect 21 22 29 30
rect 21 18 23 22
rect 27 18 29 22
rect 21 10 29 18
rect 31 10 36 30
rect 38 22 47 30
rect 38 18 40 22
rect 44 18 47 22
rect 38 16 47 18
rect 49 29 56 30
rect 49 25 51 29
rect 55 25 56 29
rect 49 22 56 25
rect 49 18 51 22
rect 55 18 56 22
rect 49 16 56 18
rect 38 15 45 16
rect 38 11 40 15
rect 44 11 45 15
rect 38 10 45 11
<< pdiffusion >>
rect 2 69 9 70
rect 2 65 3 69
rect 7 65 9 69
rect 2 62 9 65
rect 2 58 3 62
rect 7 58 9 62
rect 2 46 9 58
rect 11 61 19 70
rect 11 57 13 61
rect 17 57 19 61
rect 11 54 19 57
rect 11 50 13 54
rect 17 50 19 54
rect 11 46 19 50
rect 21 69 29 70
rect 21 65 23 69
rect 27 65 29 69
rect 21 62 29 65
rect 21 58 23 62
rect 27 58 29 62
rect 21 46 29 58
rect 31 61 39 70
rect 31 57 33 61
rect 37 57 39 61
rect 31 54 39 57
rect 31 50 33 54
rect 37 50 39 54
rect 31 46 39 50
rect 41 69 49 70
rect 41 65 43 69
rect 47 65 49 69
rect 41 62 49 65
rect 41 58 43 62
rect 47 58 49 62
rect 41 46 49 58
rect 43 43 49 46
rect 51 56 56 70
rect 51 55 58 56
rect 51 51 53 55
rect 57 51 58 55
rect 51 48 58 51
rect 51 44 53 48
rect 57 44 58 48
rect 51 43 58 44
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect -2 69 66 78
rect -2 68 3 69
rect 2 65 3 68
rect 7 68 23 69
rect 7 65 8 68
rect 2 62 8 65
rect 22 65 23 68
rect 27 68 43 69
rect 27 65 28 68
rect 22 62 28 65
rect 42 65 43 68
rect 47 68 66 69
rect 47 65 48 68
rect 2 58 3 62
rect 7 58 8 62
rect 13 61 17 62
rect 22 58 23 62
rect 27 58 28 62
rect 33 61 38 63
rect 13 54 17 57
rect 37 57 38 61
rect 42 62 48 65
rect 42 58 43 62
rect 47 58 48 62
rect 33 54 38 57
rect 53 55 57 56
rect 2 50 13 54
rect 17 50 33 54
rect 37 50 38 54
rect 2 22 6 50
rect 42 46 46 55
rect 53 48 57 51
rect 10 38 14 39
rect 17 38 23 46
rect 33 42 50 46
rect 46 39 50 42
rect 17 34 26 38
rect 30 34 31 38
rect 35 34 36 38
rect 40 34 41 38
rect 46 34 50 35
rect 10 30 14 34
rect 35 30 41 34
rect 53 30 57 44
rect 10 29 57 30
rect 10 26 51 29
rect 55 26 57 29
rect 51 22 55 25
rect 2 18 23 22
rect 27 18 31 22
rect 39 18 40 22
rect 44 18 45 22
rect 39 15 45 18
rect 51 17 55 18
rect 5 12 6 15
rect -2 11 6 12
rect 10 12 11 15
rect 39 12 40 15
rect 10 11 40 12
rect 44 12 45 15
rect 44 11 66 12
rect -2 2 66 11
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
<< ntransistor >>
rect 12 10 14 30
rect 19 10 21 30
rect 29 10 31 30
rect 36 10 38 30
rect 47 16 49 30
<< ptransistor >>
rect 9 46 11 70
rect 19 46 21 70
rect 29 46 31 70
rect 39 46 41 70
rect 49 43 51 70
<< polycontact >>
rect 10 34 14 38
rect 26 34 30 38
rect 36 34 40 38
rect 46 35 50 39
<< ndcontact >>
rect 6 11 10 15
rect 23 18 27 22
rect 40 18 44 22
rect 51 25 55 29
rect 51 18 55 22
rect 40 11 44 15
<< pdcontact >>
rect 3 65 7 69
rect 3 58 7 62
rect 13 57 17 61
rect 13 50 17 54
rect 23 65 27 69
rect 23 58 27 62
rect 33 57 37 61
rect 33 50 37 54
rect 43 65 47 69
rect 43 58 47 62
rect 53 51 57 55
rect 53 44 57 48
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
<< psubstratepdiff >>
rect 0 2 64 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 64 2
rect 0 -3 64 -2
<< nsubstratendiff >>
rect 0 82 64 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 64 82
rect 0 77 64 78
<< labels >>
rlabel polycontact 12 36 12 36 6 an
rlabel polycontact 38 36 38 36 6 an
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 20 12 20 6 z
rlabel metal1 20 20 20 20 6 z
rlabel metal1 12 32 12 32 6 an
rlabel metal1 20 40 20 40 6 b
rlabel metal1 20 52 20 52 6 z
rlabel metal1 12 52 12 52 6 z
rlabel metal1 32 6 32 6 6 vss
rlabel metal1 28 20 28 20 6 z
rlabel polycontact 28 36 28 36 6 b
rlabel metal1 36 44 36 44 6 a
rlabel metal1 28 52 28 52 6 z
rlabel pdcontact 36 60 36 60 6 z
rlabel metal1 32 74 32 74 6 vdd
rlabel metal1 38 32 38 32 6 an
rlabel metal1 44 48 44 48 6 a
rlabel metal1 53 23 53 23 6 an
rlabel metal1 55 41 55 41 6 an
<< end >>
