magic
tech scmos
timestamp 1185039137
<< checkpaint >>
rect -22 -24 72 124
<< ab >>
rect 0 0 50 100
<< pwell >>
rect -2 -4 52 49
<< nwell >>
rect -2 49 52 104
<< polysilicon >>
rect 11 85 13 88
rect 23 85 25 88
rect 35 85 37 88
rect 11 63 13 65
rect 11 62 19 63
rect 11 58 14 62
rect 18 58 19 62
rect 11 57 19 58
rect 3 52 9 53
rect 3 48 4 52
rect 8 51 9 52
rect 23 51 25 65
rect 8 49 25 51
rect 8 48 9 49
rect 3 47 9 48
rect 11 42 19 43
rect 11 38 14 42
rect 18 38 19 42
rect 11 37 19 38
rect 11 35 13 37
rect 23 35 25 49
rect 35 43 37 65
rect 35 42 43 43
rect 35 39 38 42
rect 31 38 38 39
rect 42 38 43 42
rect 31 37 43 38
rect 31 35 33 37
rect 11 22 13 25
rect 23 12 25 15
rect 31 12 33 15
<< ndiffusion >>
rect 3 32 11 35
rect 3 28 4 32
rect 8 28 11 32
rect 3 25 11 28
rect 13 25 23 35
rect 15 15 23 25
rect 25 15 31 35
rect 33 22 41 35
rect 33 18 36 22
rect 40 18 41 22
rect 33 15 41 18
rect 15 12 21 15
rect 15 8 16 12
rect 20 8 21 12
rect 15 7 21 8
<< pdiffusion >>
rect 15 92 21 93
rect 15 88 16 92
rect 20 88 21 92
rect 39 92 45 93
rect 39 88 40 92
rect 44 88 45 92
rect 15 85 21 88
rect 39 85 45 88
rect 3 82 11 85
rect 3 78 4 82
rect 8 78 11 82
rect 3 72 11 78
rect 3 68 4 72
rect 8 68 11 72
rect 3 65 11 68
rect 13 65 23 85
rect 25 82 35 85
rect 25 78 28 82
rect 32 78 35 82
rect 25 72 35 78
rect 25 68 28 72
rect 32 68 35 72
rect 25 65 35 68
rect 37 65 45 85
<< metal1 >>
rect -2 92 52 101
rect -2 88 16 92
rect 20 88 40 92
rect 44 88 52 92
rect -2 87 52 88
rect 3 82 9 83
rect 27 82 33 83
rect 3 78 4 82
rect 8 78 9 82
rect 3 77 9 78
rect 4 73 8 77
rect 3 72 9 73
rect 3 68 4 72
rect 8 68 9 72
rect 3 67 9 68
rect 4 53 8 67
rect 17 63 23 82
rect 13 62 23 63
rect 13 58 14 62
rect 18 58 23 62
rect 13 57 23 58
rect 3 52 9 53
rect 3 48 4 52
rect 8 48 9 52
rect 3 47 9 48
rect 4 33 8 47
rect 17 43 23 57
rect 13 42 23 43
rect 13 38 14 42
rect 18 38 23 42
rect 13 37 23 38
rect 3 32 9 33
rect 3 28 4 32
rect 8 28 9 32
rect 3 27 9 28
rect 17 18 23 37
rect 27 78 28 82
rect 32 78 33 82
rect 27 72 33 78
rect 27 68 28 72
rect 32 68 33 72
rect 27 23 33 68
rect 37 42 43 82
rect 37 38 38 42
rect 42 38 43 42
rect 37 28 43 38
rect 27 22 41 23
rect 27 18 36 22
rect 40 18 41 22
rect 27 17 41 18
rect -2 12 52 13
rect -2 8 16 12
rect 20 8 52 12
rect -2 4 4 8
rect 8 4 28 8
rect 32 4 42 8
rect 46 4 52 8
rect -2 -1 52 4
<< ntransistor >>
rect 11 25 13 35
rect 23 15 25 35
rect 31 15 33 35
<< ptransistor >>
rect 11 65 13 85
rect 23 65 25 85
rect 35 65 37 85
<< polycontact >>
rect 14 58 18 62
rect 4 48 8 52
rect 14 38 18 42
rect 38 38 42 42
<< ndcontact >>
rect 4 28 8 32
rect 36 18 40 22
rect 16 8 20 12
<< pdcontact >>
rect 16 88 20 92
rect 40 88 44 92
rect 4 78 8 82
rect 4 68 8 72
rect 28 78 32 82
rect 28 68 32 72
<< psubstratepcontact >>
rect 4 4 8 8
rect 28 4 32 8
rect 42 4 46 8
<< psubstratepdiff >>
rect 3 8 9 15
rect 3 4 4 8
rect 8 4 9 8
rect 27 8 47 9
rect 3 3 9 4
rect 27 4 28 8
rect 32 4 42 8
rect 46 4 47 8
rect 27 3 47 4
<< labels >>
rlabel metal1 20 50 20 50 6 i1
rlabel metal1 20 50 20 50 6 i1
rlabel metal1 25 6 25 6 6 vss
rlabel metal1 25 6 25 6 6 vss
rlabel metal1 30 50 30 50 6 q
rlabel metal1 30 50 30 50 6 q
rlabel metal1 25 94 25 94 6 vdd
rlabel metal1 25 94 25 94 6 vdd
rlabel metal1 40 55 40 55 6 i0
rlabel metal1 40 55 40 55 6 i0
<< end >>
