magic
tech scmos
timestamp 1179385827
<< checkpaint >>
rect -22 -22 54 94
<< ab >>
rect 0 0 32 72
<< pwell >>
rect -4 -4 36 32
<< nwell >>
rect -4 32 36 76
<< polysilicon >>
rect 10 65 12 69
rect 20 57 22 61
rect 10 36 12 41
rect 20 36 22 41
rect 10 35 30 36
rect 10 34 25 35
rect 10 26 12 34
rect 20 31 25 34
rect 29 31 30 35
rect 20 30 30 31
rect 20 26 22 30
rect 10 11 12 16
rect 20 11 22 16
<< ndiffusion >>
rect 2 18 10 26
rect 2 14 3 18
rect 7 16 10 18
rect 12 25 20 26
rect 12 21 14 25
rect 18 21 20 25
rect 12 16 20 21
rect 22 21 30 26
rect 22 17 25 21
rect 29 17 30 21
rect 22 16 30 17
rect 7 14 8 16
rect 2 13 8 14
<< pdiffusion >>
rect 2 64 10 65
rect 2 60 4 64
rect 8 60 10 64
rect 2 57 10 60
rect 2 53 4 57
rect 8 53 10 57
rect 2 41 10 53
rect 12 57 17 65
rect 12 50 20 57
rect 12 46 14 50
rect 18 46 20 50
rect 12 41 20 46
rect 22 56 30 57
rect 22 52 24 56
rect 28 52 30 56
rect 22 49 30 52
rect 22 45 24 49
rect 28 45 30 49
rect 22 41 30 45
<< metal1 >>
rect -2 68 34 72
rect -2 64 23 68
rect 27 64 34 68
rect 3 60 4 64
rect 8 60 9 64
rect 3 57 9 60
rect 3 53 4 57
rect 8 53 9 57
rect 23 56 29 64
rect 23 52 24 56
rect 28 52 29 56
rect 2 46 14 50
rect 18 46 19 50
rect 23 49 29 52
rect 2 27 6 46
rect 23 45 24 49
rect 28 45 29 49
rect 17 38 30 42
rect 24 35 30 38
rect 24 31 25 35
rect 29 31 30 35
rect 26 29 30 31
rect 2 25 22 27
rect 2 21 14 25
rect 18 21 22 25
rect 25 21 29 22
rect 2 14 3 18
rect 7 14 8 18
rect 2 8 8 14
rect 25 8 29 17
rect -2 4 4 8
rect 8 4 24 8
rect 28 4 34 8
rect -2 0 34 4
<< ntransistor >>
rect 10 16 12 26
rect 20 16 22 26
<< ptransistor >>
rect 10 41 12 65
rect 20 41 22 57
<< polycontact >>
rect 25 31 29 35
<< ndcontact >>
rect 3 14 7 18
rect 14 21 18 25
rect 25 17 29 21
<< pdcontact >>
rect 4 60 8 64
rect 4 53 8 57
rect 14 46 18 50
rect 24 52 28 56
rect 24 45 28 49
<< psubstratepcontact >>
rect 4 4 8 8
rect 24 4 28 8
<< nsubstratencontact >>
rect 23 64 27 68
<< psubstratepdiff >>
rect 3 8 29 9
rect 3 4 4 8
rect 8 4 24 8
rect 28 4 29 8
rect 3 3 29 4
<< nsubstratendiff >>
rect 22 68 28 69
rect 22 64 23 68
rect 27 64 28 68
rect 22 63 28 64
<< labels >>
rlabel metal1 4 32 4 32 6 z
rlabel metal1 12 24 12 24 6 z
rlabel metal1 12 48 12 48 6 z
rlabel metal1 16 4 16 4 6 vss
rlabel metal1 20 24 20 24 6 z
rlabel metal1 20 40 20 40 6 a
rlabel metal1 16 68 16 68 6 vdd
rlabel polycontact 28 32 28 32 6 a
<< end >>
