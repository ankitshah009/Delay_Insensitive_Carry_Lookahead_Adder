.subckt oai21v0x1 a1 a2 b vdd vss z
*   SPICE3 file   created from oai21v0x1.ext -      technology: scmos
m00 z      b      vdd    vdd p w=14u  l=2.3636u ad=60.439p  pd=23.9024u as=102.78p  ps=38.2439u
m01 w1     a2     z      vdd p w=27u  l=2.3636u ad=67.5p    pd=32u      as=116.561p ps=46.0976u
m02 vdd    a1     w1     vdd p w=27u  l=2.3636u ad=198.22p  pd=73.7561u as=67.5p    ps=32u
m03 n1     b      z      vss n w=12u  l=2.3636u ad=56p      pd=26u      as=72p      ps=38u
m04 vss    a2     n1     vss n w=12u  l=2.3636u ad=48p      pd=20u      as=56p      ps=26u
m05 n1     a1     vss    vss n w=12u  l=2.3636u ad=56p      pd=26u      as=48p      ps=20u
C0  a1     b      0.056f
C1  z      vdd    0.176f
C2  vss    n1     0.198f
C3  a2     vdd    0.033f
C4  vss    z      0.042f
C5  n1     a1     0.069f
C6  vss    a2     0.019f
C7  z      a1     0.016f
C8  w1     a2     0.017f
C9  n1     b      0.083f
C10 z      b      0.212f
C11 a1     a2     0.170f
C12 w1     vdd    0.005f
C13 a2     b      0.208f
C14 a1     vdd    0.020f
C15 b      vdd    0.018f
C16 vss    a1     0.026f
C17 n1     z      0.048f
C18 n1     a2     0.029f
C19 vss    b      0.032f
C20 n1     vdd    0.005f
C21 z      a2     0.072f
C23 z      vss    0.018f
C24 a1     vss    0.027f
C25 a2     vss    0.021f
C26 b      vss    0.033f
.ends
