.subckt nmx3_x4 cmd0 cmd1 i0 i1 i2 nq vdd vss
*   SPICE3 file   created from nmx3_x4.ext -      technology: scmos
m00 w1     i2     w2     vdd p w=19u  l=2.3636u ad=95p      pd=29.7838u as=114.339p ps=38u
m01 w3     cmd1   w1     vdd p w=18u  l=2.3636u ad=124.364p pd=41.2364u as=90p      ps=28.2162u
m02 w4     cmd1   vdd    vdd p w=14u  l=2.3636u ad=112p     pd=44u      as=92.5556p ps=28.1728u
m03 w5     w4     w3     vdd p w=19u  l=2.3636u ad=57p      pd=25u      as=131.273p ps=43.5273u
m04 w2     i1     w5     vdd p w=19u  l=2.3636u ad=114.339p pd=38u      as=57p      ps=25u
m05 vdd    w6     w2     vdd p w=18u  l=2.3636u ad=119p     pd=36.2222u as=108.321p ps=36u
m06 w7     cmd0   vdd    vdd p w=18u  l=2.3636u ad=54p      pd=24u      as=119p     ps=36.2222u
m07 w3     i0     w7     vdd p w=18u  l=2.3636u ad=124.364p pd=41.2364u as=54p      ps=24u
m08 w4     cmd1   vss    vss n w=8u   l=2.3636u ad=64p      pd=32u      as=59.6444p ps=21.5111u
m09 vdd    cmd0   w6     vdd p w=14u  l=2.3636u ad=92.5556p pd=28.1728u as=112p     ps=44u
m10 nq     w8     vdd    vdd p w=39u  l=2.3636u ad=195p     pd=49u      as=257.833p ps=78.4815u
m11 vdd    w8     nq     vdd p w=39u  l=2.3636u ad=257.833p pd=78.4815u as=195p     ps=49u
m12 w8     w3     vdd    vdd p w=20u  l=2.3636u ad=160p     pd=56u      as=132.222p ps=40.2469u
m13 w9     i2     w10    vss n w=12u  l=2.3636u ad=60p      pd=22u      as=82p      ps=31.3333u
m14 w3     w4     w9     vss n w=12u  l=2.3636u ad=100p     pd=37.3333u as=60p      ps=22u
m15 w11    cmd1   w3     vss n w=12u  l=2.3636u ad=36p      pd=18u      as=100p     ps=37.3333u
m16 w10    i1     w11    vss n w=12u  l=2.3636u ad=82p      pd=31.3333u as=36p      ps=18u
m17 vss    cmd0   w6     vss n w=8u   l=2.3636u ad=59.6444p pd=21.5111u as=64p      ps=32u
m18 vss    cmd0   w10    vss n w=12u  l=2.3636u ad=89.4667p pd=32.2667u as=82p      ps=31.3333u
m19 w12    w6     vss    vss n w=12u  l=2.3636u ad=36p      pd=18u      as=89.4667p ps=32.2667u
m20 w3     i0     w12    vss n w=12u  l=2.3636u ad=100p     pd=37.3333u as=36p      ps=18u
m21 nq     w8     vss    vss n w=20u  l=2.3636u ad=118p     pd=36u      as=149.111p ps=53.7778u
m22 vss    w8     nq     vss n w=20u  l=2.3636u ad=149.111p pd=53.7778u as=118p     ps=36u
m23 w8     w3     vss    vss n w=10u  l=2.3636u ad=80p      pd=36u      as=74.5556p ps=26.8889u
C0  w10    w4     0.126f
C1  vss    w6     0.077f
C2  w3     vdd    0.280f
C3  vdd    i2     0.008f
C4  w6     i1     0.130f
C5  cmd0   w4     0.026f
C6  i0     cmd1   0.008f
C7  w10    w3     0.111f
C8  w3     cmd0   0.211f
C9  vss    w4     0.039f
C10 w10    i2     0.012f
C11 w2     vdd    0.304f
C12 w6     cmd1   0.045f
C13 i1     w4     0.159f
C14 cmd0   i2     0.013f
C15 vss    w3     0.337f
C16 w3     i1     0.114f
C17 w8     i0     0.029f
C18 vss    i2     0.008f
C19 w11    w10    0.012f
C20 w4     cmd1   0.391f
C21 i1     i2     0.057f
C22 nq     w8     0.075f
C23 w2     i1     0.022f
C24 vdd    cmd0   0.016f
C25 w8     w6     0.033f
C26 w3     cmd1   0.048f
C27 w11    vss    0.004f
C28 cmd1   i2     0.195f
C29 w5     w2     0.012f
C30 nq     i0     0.027f
C31 vdd    i1     0.017f
C32 i0     w6     0.288f
C33 w2     cmd1   0.106f
C34 w10    vss    0.293f
C35 w1     w2     0.019f
C36 w5     vdd    0.011f
C37 w3     w8     0.361f
C38 w10    i1     0.022f
C39 vss    cmd0   0.016f
C40 nq     w6     0.063f
C41 cmd0   i1     0.077f
C42 i0     w4     0.015f
C43 vdd    cmd1   0.107f
C44 w10    cmd1   0.005f
C45 w1     vdd    0.019f
C46 vss    i1     0.015f
C47 w3     i0     0.171f
C48 w6     w4     0.038f
C49 cmd0   cmd1   0.030f
C50 nq     w3     0.367f
C51 vss    cmd1   0.045f
C52 w8     vdd    0.081f
C53 w3     w6     0.359f
C54 i1     cmd1   0.140f
C55 w6     i2     0.022f
C56 vdd    i0     0.026f
C57 w8     cmd0   0.066f
C58 w3     w4     0.140f
C59 w12    vss    0.010f
C60 w9     w10    0.019f
C61 w4     i2     0.168f
C62 vss    w8     0.026f
C63 nq     vdd    0.142f
C64 i0     cmd0   0.328f
C65 w3     i2     0.014f
C66 w2     w4     0.068f
C67 vdd    w6     0.021f
C68 w9     vss    0.007f
C69 w10    w6     0.020f
C70 w3     w2     0.160f
C71 w7     vdd    0.011f
C72 vss    i0     0.022f
C73 nq     cmd0   0.003f
C74 i0     i1     0.029f
C75 vdd    w4     0.043f
C76 w2     i2     0.010f
C77 cmd0   w6     0.369f
C78 nq     vss    0.025f
C79 nq     vss    0.010f
C81 w3     vss    0.084f
C82 w8     vss    0.060f
C84 i0     vss    0.048f
C85 cmd0   vss    0.068f
C86 w6     vss    0.054f
C87 i1     vss    0.038f
C88 w4     vss    0.049f
C89 cmd1   vss    0.072f
C90 i2     vss    0.036f
.ends
