magic
tech scmos
timestamp 1180640047
<< checkpaint >>
rect -24 -26 94 126
<< ab >>
rect 0 0 70 100
<< pwell >>
rect -4 -6 74 49
<< nwell >>
rect -4 49 74 106
<< polysilicon >>
rect 15 76 17 81
rect 23 76 25 81
rect 35 76 37 81
rect 43 76 45 81
rect 57 74 59 79
rect 15 53 17 56
rect 8 52 17 53
rect 8 48 9 52
rect 13 50 17 52
rect 13 48 19 50
rect 8 47 19 48
rect 7 42 13 43
rect 7 38 8 42
rect 12 38 13 42
rect 7 37 13 38
rect 11 26 13 37
rect 17 37 19 47
rect 23 43 25 56
rect 35 53 37 56
rect 29 52 37 53
rect 29 48 30 52
rect 34 48 37 52
rect 29 47 37 48
rect 23 42 33 43
rect 23 41 28 42
rect 27 38 28 41
rect 32 38 33 42
rect 27 37 33 38
rect 17 34 21 37
rect 19 26 21 34
rect 31 26 33 37
rect 43 37 45 56
rect 57 53 59 56
rect 51 52 59 53
rect 51 48 52 52
rect 56 48 59 52
rect 51 47 59 48
rect 43 36 52 37
rect 43 33 47 36
rect 39 32 47 33
rect 51 32 52 36
rect 39 31 52 32
rect 39 26 41 31
rect 57 26 59 47
rect 11 12 13 17
rect 19 12 21 17
rect 31 12 33 17
rect 39 12 41 17
rect 57 12 59 17
<< ndiffusion >>
rect 3 17 11 26
rect 13 17 19 26
rect 21 22 31 26
rect 21 18 24 22
rect 28 18 31 22
rect 21 17 31 18
rect 33 17 39 26
rect 41 22 57 26
rect 41 18 48 22
rect 52 18 57 22
rect 41 17 57 18
rect 59 25 67 26
rect 59 21 62 25
rect 66 21 67 25
rect 59 20 67 21
rect 59 17 64 20
rect 3 11 9 17
rect 3 7 4 11
rect 8 7 9 11
rect 3 6 9 7
<< pdiffusion >>
rect 6 82 13 83
rect 6 78 8 82
rect 12 78 13 82
rect 47 82 55 83
rect 6 76 13 78
rect 47 78 48 82
rect 52 78 55 82
rect 47 76 55 78
rect 6 56 15 76
rect 17 56 23 76
rect 25 62 35 76
rect 25 58 28 62
rect 32 58 35 62
rect 25 56 35 58
rect 37 56 43 76
rect 45 74 55 76
rect 45 56 57 74
rect 59 70 64 74
rect 59 69 67 70
rect 59 65 62 69
rect 66 65 67 69
rect 59 61 67 65
rect 59 57 62 61
rect 66 57 67 61
rect 59 56 67 57
<< metal1 >>
rect -2 88 72 100
rect 8 82 12 88
rect 8 77 12 78
rect 48 82 52 88
rect 48 77 52 78
rect 7 68 53 72
rect 7 52 13 68
rect 7 48 9 52
rect 7 47 13 48
rect 18 53 22 63
rect 28 62 42 63
rect 32 58 42 62
rect 28 57 42 58
rect 18 52 34 53
rect 18 48 30 52
rect 18 47 34 48
rect 18 43 22 47
rect 7 42 22 43
rect 7 38 8 42
rect 12 38 22 42
rect 7 37 22 38
rect 27 42 33 43
rect 27 38 28 42
rect 32 38 33 42
rect 27 32 33 38
rect 7 28 33 32
rect 7 18 13 28
rect 38 22 42 57
rect 47 53 53 68
rect 62 69 66 70
rect 62 61 66 65
rect 47 52 57 53
rect 47 48 52 52
rect 56 48 57 52
rect 47 47 57 48
rect 62 36 66 57
rect 46 32 47 36
rect 51 32 66 36
rect 62 25 66 32
rect 23 18 24 22
rect 28 18 42 22
rect 23 17 42 18
rect 48 22 52 23
rect 62 20 66 21
rect 48 12 52 18
rect -2 11 72 12
rect -2 7 4 11
rect 8 7 72 11
rect -2 0 72 7
<< ntransistor >>
rect 11 17 13 26
rect 19 17 21 26
rect 31 17 33 26
rect 39 17 41 26
rect 57 17 59 26
<< ptransistor >>
rect 15 56 17 76
rect 23 56 25 76
rect 35 56 37 76
rect 43 56 45 76
rect 57 56 59 74
<< polycontact >>
rect 9 48 13 52
rect 8 38 12 42
rect 30 48 34 52
rect 28 38 32 42
rect 52 48 56 52
rect 47 32 51 36
<< ndcontact >>
rect 24 18 28 22
rect 48 18 52 22
rect 62 21 66 25
rect 4 7 8 11
<< pdcontact >>
rect 8 78 12 82
rect 48 78 52 82
rect 28 58 32 62
rect 62 65 66 69
rect 62 57 66 61
<< psubstratepcontact >>
rect 18 4 22 8
rect 28 4 32 8
<< nsubstratencontact >>
rect 8 92 12 96
rect 18 92 22 96
<< psubstratepdiff >>
rect 17 8 33 9
rect 17 4 18 8
rect 22 4 28 8
rect 32 4 33 8
rect 17 3 33 4
<< nsubstratendiff >>
rect 7 96 23 97
rect 7 92 8 96
rect 12 92 18 96
rect 22 92 23 96
rect 7 91 23 92
<< labels >>
rlabel polysilicon 47 34 47 34 6 sn
rlabel metal1 10 25 10 25 6 a0
rlabel metal1 10 25 10 25 6 a0
rlabel metal1 20 30 20 30 6 a0
rlabel metal1 20 30 20 30 6 a0
rlabel polycontact 10 40 10 40 6 a1
rlabel polycontact 10 40 10 40 6 a1
rlabel metal1 20 50 20 50 6 a1
rlabel metal1 20 50 20 50 6 a1
rlabel metal1 10 60 10 60 6 s
rlabel metal1 10 60 10 60 6 s
rlabel metal1 20 70 20 70 6 s
rlabel metal1 20 70 20 70 6 s
rlabel metal1 35 6 35 6 6 vss
rlabel metal1 35 6 35 6 6 vss
rlabel metal1 30 20 30 20 6 z
rlabel metal1 30 20 30 20 6 z
rlabel metal1 30 35 30 35 6 a0
rlabel metal1 30 35 30 35 6 a0
rlabel metal1 30 50 30 50 6 a1
rlabel metal1 30 50 30 50 6 a1
rlabel pdcontact 30 60 30 60 6 z
rlabel pdcontact 30 60 30 60 6 z
rlabel metal1 30 70 30 70 6 s
rlabel metal1 30 70 30 70 6 s
rlabel metal1 35 94 35 94 6 vdd
rlabel metal1 35 94 35 94 6 vdd
rlabel metal1 40 40 40 40 6 z
rlabel metal1 40 40 40 40 6 z
rlabel metal1 50 60 50 60 6 s
rlabel metal1 50 60 50 60 6 s
rlabel metal1 40 70 40 70 6 s
rlabel metal1 40 70 40 70 6 s
rlabel metal1 56 34 56 34 6 sn
rlabel metal1 64 45 64 45 6 sn
<< end >>
