.subckt oai22v0x05 a1 a2 b1 b2 vdd vss z
*   SPICE3 file   created from oai22v0x05.ext -      technology: scmos
m00 w1     b1     vdd    vdd p w=16u  l=2.3636u ad=48p      pd=22u      as=145.5p   ps=53u
m01 z      b2     w1     vdd p w=16u  l=2.3636u ad=64p      pd=24u      as=48p      ps=22u
m02 w2     a2     z      vdd p w=16u  l=2.3636u ad=48p      pd=22u      as=64p      ps=24u
m03 vdd    a1     w2     vdd p w=16u  l=2.3636u ad=145.5p   pd=53u      as=48p      ps=22u
m04 n3     b2     z      vss n w=7u   l=2.3636u ad=38.5p    pd=21.5u    as=45.5p    ps=23u
m05 vss    a2     n3     vss n w=7u   l=2.3636u ad=74.5p    pd=33u      as=38.5p    ps=21.5u
m06 z      b1     n3     vss n w=7u   l=2.3636u ad=45.5p    pd=23u      as=38.5p    ps=21.5u
m07 n3     a1     vss    vss n w=7u   l=2.3636u ad=38.5p    pd=21.5u    as=74.5p    ps=33u
C0  w2     vdd    0.003f
C1  a1     a2     0.110f
C2  w1     b2     0.005f
C3  z      b1     0.205f
C4  a1     b1     0.029f
C5  a2     b2     0.085f
C6  w1     vdd    0.003f
C7  n3     z      0.185f
C8  b2     b1     0.149f
C9  a2     vdd    0.019f
C10 vss    a2     0.047f
C11 n3     a1     0.021f
C12 b1     vdd    0.018f
C13 n3     b2     0.025f
C14 z      a1     0.048f
C15 vss    b1     0.020f
C16 n3     vdd    0.006f
C17 z      b2     0.090f
C18 vss    n3     0.305f
C19 z      vdd    0.212f
C20 a1     b2     0.059f
C21 vss    z      0.040f
C22 a2     b1     0.043f
C23 a1     vdd    0.067f
C24 vss    a1     0.014f
C25 b2     vdd    0.025f
C26 z      w1     0.012f
C27 n3     a2     0.133f
C28 vss    b2     0.013f
C29 w2     a1     0.023f
C30 z      a2     0.020f
C31 n3     b1     0.036f
C33 n3     vss    0.008f
C34 z      vss    0.019f
C35 a1     vss    0.028f
C36 a2     vss    0.026f
C37 b2     vss    0.024f
C38 b1     vss    0.027f
.ends
