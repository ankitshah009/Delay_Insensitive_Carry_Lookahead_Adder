magic
tech scmos
timestamp 1170759832
<< checkpaint >>
rect -22 -26 86 114
<< ab >>
rect 0 0 64 88
<< pwell >>
rect -4 -8 68 40
<< nwell >>
rect -4 40 68 96
<< polysilicon >>
rect 2 77 11 83
rect 9 74 11 77
rect 21 77 30 83
rect 34 77 43 83
rect 21 74 23 77
rect 41 74 43 77
rect 53 77 62 83
rect 53 74 55 77
rect 9 43 11 46
rect 21 43 23 46
rect 41 43 43 46
rect 53 43 55 46
rect 2 37 14 43
rect 18 37 30 43
rect 34 37 46 43
rect 50 37 62 43
rect 9 34 11 37
rect 21 34 23 37
rect 41 34 43 37
rect 53 34 55 37
rect 9 11 11 14
rect 2 5 11 11
rect 21 11 23 14
rect 41 11 43 14
rect 21 5 30 11
rect 34 5 43 11
rect 53 11 55 14
rect 53 5 62 11
<< ndiffusion >>
rect 2 14 9 34
rect 11 14 21 34
rect 23 14 30 34
rect 34 14 41 34
rect 43 14 53 34
rect 55 14 62 34
rect 13 2 19 14
rect 45 2 51 14
<< pdiffusion >>
rect 13 74 19 86
rect 45 74 51 86
rect 2 46 9 74
rect 11 46 21 74
rect 23 46 30 74
rect 34 46 41 74
rect 43 46 53 74
rect 55 46 62 74
<< metal1 >>
rect -2 86 2 90
rect 10 86 22 90
rect 30 86 34 90
rect 42 86 54 90
rect 62 86 66 90
rect 5 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 59 82
rect 13 6 14 10
rect 18 6 46 10
rect 50 6 51 10
rect -2 -2 2 2
rect 10 -2 22 2
rect 30 -2 34 2
rect 42 -2 54 2
rect 62 -2 66 2
<< metal2 >>
rect -2 86 6 90
rect 10 86 22 90
rect 26 86 38 90
rect 42 86 54 90
rect 58 86 66 90
rect -2 82 66 86
rect -2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 66 82
rect -2 76 66 78
rect -2 10 66 12
rect -2 6 14 10
rect 18 6 46 10
rect 50 6 66 10
rect -2 2 66 6
rect -2 -2 6 2
rect 10 -2 22 2
rect 26 -2 38 2
rect 42 -2 54 2
rect 58 -2 66 2
<< ntransistor >>
rect 9 14 11 34
rect 21 14 23 34
rect 41 14 43 34
rect 53 14 55 34
<< ptransistor >>
rect 9 46 11 74
rect 21 46 23 74
rect 41 46 43 74
rect 53 46 55 74
<< m2contact >>
rect 6 86 10 90
rect 22 86 26 90
rect 38 86 42 90
rect 54 86 58 90
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 14 6 18 10
rect 46 6 50 10
rect 6 -2 10 2
rect 22 -2 26 2
rect 38 -2 42 2
rect 54 -2 58 2
<< psubstratepcontact >>
rect 2 -2 6 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 58 -2 62 2
<< nsubstratencontact >>
rect 2 86 6 90
rect 26 86 30 90
rect 34 86 38 90
rect 58 86 62 90
<< psubstratepdiff >>
rect 0 2 7 3
rect 25 2 39 3
rect 57 2 64 3
rect 0 -2 2 2
rect 6 -2 7 2
rect 0 -3 7 -2
rect 25 -2 26 2
rect 30 -2 34 2
rect 38 -2 39 2
rect 25 -3 39 -2
rect 57 -2 58 2
rect 62 -2 64 2
rect 57 -3 64 -2
<< nsubstratendiff >>
rect 0 90 7 91
rect 0 86 2 90
rect 6 86 7 90
rect 25 90 39 91
rect 25 86 26 90
rect 30 86 34 90
rect 38 86 39 90
rect 57 90 64 91
rect 57 86 58 90
rect 62 86 64 90
rect 0 85 7 86
rect 25 85 39 86
rect 57 85 64 86
<< labels >>
rlabel metal2 32 6 32 6 6 vss
rlabel metal2 32 82 32 82 6 vdd
<< end >>
