magic
tech scmos
timestamp 1179386826
<< checkpaint >>
rect -22 -25 102 105
<< ab >>
rect 0 0 80 80
<< pwell >>
rect -4 -7 84 36
<< nwell >>
rect -4 36 84 87
<< polysilicon >>
rect 9 70 11 74
rect 16 70 18 74
rect 26 70 28 74
rect 33 70 35 74
rect 43 70 45 74
rect 50 70 52 74
rect 60 70 62 74
rect 67 70 69 74
rect 9 34 11 43
rect 16 40 18 43
rect 26 40 28 43
rect 33 40 35 43
rect 43 40 45 43
rect 16 38 29 40
rect 33 38 45 40
rect 50 39 52 43
rect 60 39 62 43
rect 50 38 62 39
rect 67 38 69 43
rect 23 34 24 38
rect 28 34 29 38
rect 9 33 19 34
rect 9 32 14 33
rect 13 29 14 32
rect 18 29 19 33
rect 13 28 19 29
rect 23 33 29 34
rect 36 37 42 38
rect 36 33 37 37
rect 41 33 42 37
rect 50 34 51 38
rect 55 34 62 38
rect 13 25 15 28
rect 23 25 25 33
rect 36 32 42 33
rect 47 32 62 34
rect 66 37 72 38
rect 66 33 67 37
rect 71 33 72 37
rect 66 32 72 33
rect 37 29 39 32
rect 47 29 49 32
rect 59 29 61 32
rect 69 29 71 32
rect 13 6 15 10
rect 23 6 25 10
rect 37 6 39 10
rect 47 6 49 10
rect 59 6 61 10
rect 69 6 71 10
<< ndiffusion >>
rect 27 25 37 29
rect 4 15 13 25
rect 4 11 7 15
rect 11 11 13 15
rect 4 10 13 11
rect 15 22 23 25
rect 15 18 17 22
rect 21 18 23 22
rect 15 10 23 18
rect 25 15 37 25
rect 25 11 29 15
rect 33 11 37 15
rect 25 10 37 11
rect 39 22 47 29
rect 39 18 41 22
rect 45 18 47 22
rect 39 10 47 18
rect 49 15 59 29
rect 49 11 52 15
rect 56 11 59 15
rect 49 10 59 11
rect 61 22 69 29
rect 61 18 63 22
rect 67 18 69 22
rect 61 10 69 18
rect 71 22 78 29
rect 71 18 73 22
rect 77 18 78 22
rect 71 15 78 18
rect 71 11 73 15
rect 77 11 78 15
rect 71 10 78 11
<< pdiffusion >>
rect 2 69 9 70
rect 2 65 3 69
rect 7 65 9 69
rect 2 62 9 65
rect 2 58 3 62
rect 7 58 9 62
rect 2 43 9 58
rect 11 43 16 70
rect 18 56 26 70
rect 18 52 20 56
rect 24 52 26 56
rect 18 48 26 52
rect 18 44 20 48
rect 24 44 26 48
rect 18 43 26 44
rect 28 43 33 70
rect 35 69 43 70
rect 35 65 37 69
rect 41 65 43 69
rect 35 62 43 65
rect 35 58 37 62
rect 41 58 43 62
rect 35 43 43 58
rect 45 43 50 70
rect 52 56 60 70
rect 52 52 54 56
rect 58 52 60 56
rect 52 48 60 52
rect 52 44 54 48
rect 58 44 60 48
rect 52 43 60 44
rect 62 43 67 70
rect 69 69 77 70
rect 69 65 71 69
rect 75 65 77 69
rect 69 62 77 65
rect 69 58 71 62
rect 75 58 77 62
rect 69 43 77 58
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect -2 69 82 78
rect -2 68 3 69
rect 2 65 3 68
rect 7 68 37 69
rect 7 65 8 68
rect 2 62 8 65
rect 2 58 3 62
rect 7 58 8 62
rect 36 65 37 68
rect 41 68 71 69
rect 41 65 42 68
rect 36 62 42 65
rect 36 58 37 62
rect 41 58 42 62
rect 70 65 71 68
rect 75 68 82 69
rect 75 65 76 68
rect 70 62 76 65
rect 70 58 71 62
rect 75 58 76 62
rect 18 56 24 57
rect 18 52 20 56
rect 54 56 58 57
rect 24 52 54 54
rect 58 52 63 54
rect 18 50 63 52
rect 18 48 24 50
rect 18 47 20 48
rect 2 44 20 47
rect 54 48 58 50
rect 2 42 24 44
rect 29 42 49 46
rect 54 43 58 44
rect 2 22 6 42
rect 29 38 33 42
rect 45 38 49 42
rect 23 34 24 38
rect 28 34 33 38
rect 37 37 41 38
rect 14 33 18 34
rect 45 34 51 38
rect 55 34 56 38
rect 65 37 71 38
rect 37 30 41 33
rect 65 33 67 37
rect 65 30 71 33
rect 18 29 71 30
rect 14 26 71 29
rect 2 18 17 22
rect 21 18 41 22
rect 45 18 63 22
rect 67 18 68 22
rect 72 18 73 22
rect 77 18 78 22
rect 72 15 78 18
rect 6 12 7 15
rect -2 11 7 12
rect 11 12 12 15
rect 28 12 29 15
rect 11 11 29 12
rect 33 12 34 15
rect 51 12 52 15
rect 33 11 52 12
rect 56 12 57 15
rect 72 12 73 15
rect 56 11 73 12
rect 77 12 78 15
rect 77 11 82 12
rect -2 2 82 11
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
<< ntransistor >>
rect 13 10 15 25
rect 23 10 25 25
rect 37 10 39 29
rect 47 10 49 29
rect 59 10 61 29
rect 69 10 71 29
<< ptransistor >>
rect 9 43 11 70
rect 16 43 18 70
rect 26 43 28 70
rect 33 43 35 70
rect 43 43 45 70
rect 50 43 52 70
rect 60 43 62 70
rect 67 43 69 70
<< polycontact >>
rect 24 34 28 38
rect 14 29 18 33
rect 37 33 41 37
rect 51 34 55 38
rect 67 33 71 37
<< ndcontact >>
rect 7 11 11 15
rect 17 18 21 22
rect 29 11 33 15
rect 41 18 45 22
rect 52 11 56 15
rect 63 18 67 22
rect 73 18 77 22
rect 73 11 77 15
<< pdcontact >>
rect 3 65 7 69
rect 3 58 7 62
rect 20 52 24 56
rect 20 44 24 48
rect 37 65 41 69
rect 37 58 41 62
rect 54 52 58 56
rect 54 44 58 48
rect 71 65 75 69
rect 71 58 75 62
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
<< psubstratepdiff >>
rect 0 2 80 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 80 2
rect 0 -3 80 -2
<< nsubstratendiff >>
rect 0 82 80 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 80 82
rect 0 77 80 78
<< labels >>
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 20 12 20 6 z
rlabel ndcontact 20 20 20 20 6 z
rlabel metal1 20 28 20 28 6 a
rlabel metal1 28 20 28 20 6 z
rlabel metal1 28 28 28 28 6 a
rlabel metal1 12 44 12 44 6 z
rlabel metal1 28 36 28 36 6 b
rlabel metal1 28 52 28 52 6 z
rlabel metal1 20 48 20 48 6 z
rlabel metal1 40 6 40 6 6 vss
rlabel metal1 36 20 36 20 6 z
rlabel metal1 36 28 36 28 6 a
rlabel ndcontact 44 20 44 20 6 z
rlabel metal1 44 28 44 28 6 a
rlabel metal1 36 44 36 44 6 b
rlabel metal1 44 44 44 44 6 b
rlabel metal1 36 52 36 52 6 z
rlabel metal1 44 52 44 52 6 z
rlabel metal1 40 74 40 74 6 vdd
rlabel metal1 52 20 52 20 6 z
rlabel metal1 52 28 52 28 6 a
rlabel metal1 60 20 60 20 6 z
rlabel metal1 60 28 60 28 6 a
rlabel polycontact 52 36 52 36 6 b
rlabel metal1 60 52 60 52 6 z
rlabel metal1 52 52 52 52 6 z
rlabel metal1 68 32 68 32 6 a
<< end >>
