magic
tech scmos
timestamp 1185094817
<< checkpaint >>
rect -22 -22 32 122
<< ab >>
rect 0 0 10 100
<< pwell >>
rect -4 -4 14 48
<< nwell >>
rect -4 48 14 104
<< metal1 >>
rect -2 88 12 100
rect -2 0 12 12
<< labels >>
rlabel metal1 5 6 5 6 6 vss
rlabel metal1 5 94 5 94 6 vdd
<< end >>
