magic
tech scmos
timestamp 1180639968
<< checkpaint >>
rect -24 -26 94 126
<< ab >>
rect 0 0 70 100
<< pwell >>
rect -4 -6 74 49
<< nwell >>
rect -4 49 74 106
<< polysilicon >>
rect 33 89 35 94
rect 45 89 47 94
rect 11 83 13 88
rect 57 89 59 94
rect 11 52 13 63
rect 33 52 35 63
rect 45 52 47 63
rect 57 52 59 63
rect 11 51 22 52
rect 11 50 17 51
rect 15 47 17 50
rect 21 47 22 51
rect 15 46 22 47
rect 33 51 41 52
rect 33 47 36 51
rect 40 47 41 51
rect 33 46 41 47
rect 45 51 53 52
rect 45 47 48 51
rect 52 47 53 51
rect 45 46 53 47
rect 57 51 63 52
rect 57 47 58 51
rect 62 47 63 51
rect 57 46 63 47
rect 15 37 17 46
rect 33 37 35 46
rect 45 37 47 46
rect 57 42 59 46
rect 53 40 59 42
rect 53 37 55 40
rect 15 22 17 27
rect 33 25 35 30
rect 45 20 47 25
rect 53 20 55 25
<< ndiffusion >>
rect 7 36 15 37
rect 7 32 8 36
rect 12 32 15 36
rect 7 31 15 32
rect 10 27 15 31
rect 17 32 33 37
rect 17 28 20 32
rect 24 30 33 32
rect 35 36 45 37
rect 35 32 38 36
rect 42 32 45 36
rect 35 30 45 32
rect 24 28 31 30
rect 17 27 31 28
rect 40 25 45 30
rect 47 25 53 37
rect 55 32 64 37
rect 55 28 58 32
rect 62 28 64 32
rect 55 25 64 28
<< pdiffusion >>
rect 49 92 55 93
rect 49 89 50 92
rect 6 73 11 83
rect 3 72 11 73
rect 3 68 4 72
rect 8 68 11 72
rect 3 67 11 68
rect 6 63 11 67
rect 13 82 21 83
rect 13 78 16 82
rect 20 78 21 82
rect 13 75 21 78
rect 13 63 19 75
rect 28 69 33 89
rect 25 68 33 69
rect 25 64 26 68
rect 30 64 33 68
rect 25 63 33 64
rect 35 82 45 89
rect 35 78 38 82
rect 42 78 45 82
rect 35 63 45 78
rect 47 88 50 89
rect 54 89 55 92
rect 54 88 57 89
rect 47 63 57 88
rect 59 83 64 89
rect 59 82 67 83
rect 59 78 62 82
rect 66 78 67 82
rect 59 77 67 78
rect 59 63 64 77
<< metal1 >>
rect -2 92 72 100
rect -2 88 50 92
rect 54 88 72 92
rect 16 82 20 88
rect 37 78 38 82
rect 42 78 62 82
rect 66 78 67 82
rect 16 77 20 78
rect 4 72 22 73
rect 8 68 22 72
rect 4 67 22 68
rect 26 68 30 69
rect 8 36 12 67
rect 26 51 30 64
rect 38 68 53 73
rect 38 52 42 68
rect 58 63 62 73
rect 16 47 17 51
rect 21 47 30 51
rect 26 42 30 47
rect 36 51 42 52
rect 40 47 42 51
rect 36 46 42 47
rect 48 57 62 63
rect 48 51 52 57
rect 48 46 52 47
rect 57 51 63 52
rect 57 47 58 51
rect 62 47 63 51
rect 57 42 63 47
rect 26 38 42 42
rect 38 36 42 38
rect 8 27 12 32
rect 20 32 24 33
rect 38 31 42 32
rect 47 38 63 42
rect 20 12 24 28
rect 47 18 53 38
rect 58 32 62 33
rect 58 12 62 28
rect -2 0 72 12
<< ntransistor >>
rect 15 27 17 37
rect 33 30 35 37
rect 45 25 47 37
rect 53 25 55 37
<< ptransistor >>
rect 11 63 13 83
rect 33 63 35 89
rect 45 63 47 89
rect 57 63 59 89
<< polycontact >>
rect 17 47 21 51
rect 36 47 40 51
rect 48 47 52 51
rect 58 47 62 51
<< ndcontact >>
rect 8 32 12 36
rect 20 28 24 32
rect 38 32 42 36
rect 58 28 62 32
<< pdcontact >>
rect 4 68 8 72
rect 16 78 20 82
rect 26 64 30 68
rect 38 78 42 82
rect 50 88 54 92
rect 62 78 66 82
<< psubstratepcontact >>
rect 8 4 12 8
rect 18 4 22 8
<< nsubstratencontact >>
rect 8 92 12 96
<< psubstratepdiff >>
rect 7 8 23 9
rect 7 4 8 8
rect 12 4 18 8
rect 22 4 23 8
rect 7 3 23 4
<< nsubstratendiff >>
rect 7 96 13 97
rect 7 92 8 96
rect 12 92 13 96
rect 7 91 13 92
<< labels >>
rlabel polycontact 18 49 18 49 6 zn
rlabel metal1 10 50 10 50 6 z
rlabel metal1 10 50 10 50 6 z
rlabel metal1 28 53 28 53 6 zn
rlabel metal1 23 49 23 49 6 zn
rlabel metal1 20 70 20 70 6 z
rlabel metal1 20 70 20 70 6 z
rlabel metal1 35 6 35 6 6 vss
rlabel metal1 35 6 35 6 6 vss
rlabel metal1 40 36 40 36 6 zn
rlabel metal1 50 30 50 30 6 a1
rlabel metal1 50 30 50 30 6 a1
rlabel metal1 50 70 50 70 6 b
rlabel metal1 50 55 50 55 6 a2
rlabel metal1 40 60 40 60 6 b
rlabel metal1 50 70 50 70 6 b
rlabel metal1 40 60 40 60 6 b
rlabel metal1 50 55 50 55 6 a2
rlabel metal1 35 94 35 94 6 vdd
rlabel metal1 35 94 35 94 6 vdd
rlabel metal1 60 45 60 45 6 a1
rlabel metal1 60 45 60 45 6 a1
rlabel metal1 60 65 60 65 6 a2
rlabel metal1 60 65 60 65 6 a2
rlabel metal1 52 80 52 80 6 n2
<< end >>
