magic
tech scmos
timestamp 1179385035
<< checkpaint >>
rect -22 -25 62 105
<< ab >>
rect 0 0 40 80
<< pwell >>
rect -4 -7 44 36
<< nwell >>
rect -4 36 44 87
<< polysilicon >>
rect 9 70 11 74
rect 20 58 22 63
rect 30 58 32 63
rect 9 39 11 42
rect 20 39 22 50
rect 30 47 32 50
rect 29 46 35 47
rect 29 42 30 46
rect 34 42 35 46
rect 29 41 35 42
rect 9 38 15 39
rect 9 34 10 38
rect 14 34 15 38
rect 9 33 15 34
rect 19 38 25 39
rect 19 34 20 38
rect 24 34 25 38
rect 19 33 25 34
rect 9 30 11 33
rect 22 25 24 33
rect 29 25 31 41
rect 9 11 11 16
rect 22 13 24 18
rect 29 13 31 18
<< ndiffusion >>
rect 2 29 9 30
rect 2 25 3 29
rect 7 25 9 29
rect 2 21 9 25
rect 2 17 3 21
rect 7 17 9 21
rect 2 16 9 17
rect 11 25 19 30
rect 11 18 22 25
rect 24 18 29 25
rect 31 23 38 25
rect 31 19 33 23
rect 37 19 38 23
rect 31 18 38 19
rect 11 16 19 18
rect 13 12 19 16
rect 13 8 14 12
rect 18 8 19 12
rect 13 7 19 8
<< pdiffusion >>
rect 32 70 38 71
rect 4 55 9 70
rect 2 54 9 55
rect 2 50 3 54
rect 7 50 9 54
rect 2 47 9 50
rect 2 43 3 47
rect 7 43 9 47
rect 2 42 9 43
rect 11 69 18 70
rect 11 65 13 69
rect 17 65 18 69
rect 32 66 33 70
rect 37 66 38 70
rect 32 65 38 66
rect 11 62 18 65
rect 11 58 13 62
rect 17 58 18 62
rect 34 58 38 65
rect 11 50 20 58
rect 22 55 30 58
rect 22 51 24 55
rect 28 51 30 55
rect 22 50 30 51
rect 32 50 38 58
rect 11 42 18 50
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect -2 70 42 78
rect -2 69 33 70
rect -2 68 13 69
rect 12 65 13 68
rect 17 68 33 69
rect 17 65 18 68
rect 32 66 33 68
rect 37 68 42 70
rect 37 66 38 68
rect 12 62 18 65
rect 12 58 13 62
rect 17 58 18 62
rect 2 54 7 55
rect 2 50 3 54
rect 2 47 7 50
rect 2 43 3 47
rect 2 42 7 43
rect 10 51 24 55
rect 28 51 29 55
rect 2 30 6 42
rect 10 38 14 51
rect 25 42 30 46
rect 34 42 38 55
rect 17 34 20 38
rect 24 34 31 38
rect 10 30 14 34
rect 2 29 7 30
rect 2 25 3 29
rect 10 26 22 30
rect 25 26 31 34
rect 2 23 7 25
rect 18 23 22 26
rect 2 21 14 23
rect 2 17 3 21
rect 7 17 14 21
rect 18 19 33 23
rect 37 19 38 23
rect -2 8 14 12
rect 18 8 42 12
rect -2 2 42 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
<< ntransistor >>
rect 9 16 11 30
rect 22 18 24 25
rect 29 18 31 25
<< ptransistor >>
rect 9 42 11 70
rect 20 50 22 58
rect 30 50 32 58
<< polycontact >>
rect 30 42 34 46
rect 10 34 14 38
rect 20 34 24 38
<< ndcontact >>
rect 3 25 7 29
rect 3 17 7 21
rect 33 19 37 23
rect 14 8 18 12
<< pdcontact >>
rect 3 50 7 54
rect 3 43 7 47
rect 13 65 17 69
rect 33 66 37 70
rect 13 58 17 62
rect 24 51 28 55
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
<< psubstratepdiff >>
rect 0 2 40 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 40 2
rect 0 -3 40 -2
<< nsubstratendiff >>
rect 0 82 40 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 40 82
rect 0 77 40 78
<< labels >>
rlabel polycontact 12 36 12 36 6 zn
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 20 12 20 6 z
rlabel metal1 12 40 12 40 6 zn
rlabel metal1 20 6 20 6 6 vss
rlabel metal1 20 36 20 36 6 a
rlabel metal1 28 32 28 32 6 a
rlabel metal1 28 44 28 44 6 b
rlabel metal1 19 53 19 53 6 zn
rlabel metal1 20 74 20 74 6 vdd
rlabel metal1 28 21 28 21 6 zn
rlabel metal1 36 52 36 52 6 b
<< end >>
