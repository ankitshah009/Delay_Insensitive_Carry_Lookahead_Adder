magic
tech scmos
timestamp 1185038932
<< checkpaint >>
rect -22 -24 82 124
<< ab >>
rect 0 0 60 100
<< pwell >>
rect -2 -4 62 49
<< nwell >>
rect -2 49 62 104
<< polysilicon >>
rect 47 95 49 98
rect 11 85 13 88
rect 23 85 25 88
rect 35 85 37 88
rect 11 43 13 65
rect 23 63 25 65
rect 17 62 25 63
rect 17 58 18 62
rect 22 61 25 62
rect 22 58 23 61
rect 17 57 23 58
rect 35 53 37 65
rect 35 52 43 53
rect 35 51 38 52
rect 37 48 38 51
rect 42 48 43 52
rect 37 47 43 48
rect 27 46 33 47
rect 7 42 13 43
rect 7 38 8 42
rect 12 38 13 42
rect 7 37 13 38
rect 11 25 13 37
rect 17 42 23 43
rect 17 38 18 42
rect 22 38 23 42
rect 27 42 28 46
rect 32 43 33 46
rect 47 43 49 55
rect 32 42 49 43
rect 27 41 49 42
rect 17 37 23 38
rect 17 35 25 37
rect 23 25 25 35
rect 37 32 43 33
rect 37 29 38 32
rect 35 28 38 29
rect 42 28 43 32
rect 35 27 43 28
rect 35 25 37 27
rect 47 25 49 41
rect 11 12 13 15
rect 23 12 25 15
rect 35 12 37 15
rect 47 2 49 5
<< ndiffusion >>
rect 15 32 21 33
rect 15 28 16 32
rect 20 28 21 32
rect 15 25 21 28
rect 3 22 11 25
rect 3 18 4 22
rect 8 18 11 22
rect 3 15 11 18
rect 13 15 23 25
rect 25 22 35 25
rect 25 18 28 22
rect 32 18 35 22
rect 25 15 35 18
rect 37 15 47 25
rect 39 12 47 15
rect 39 8 40 12
rect 44 8 47 12
rect 39 5 47 8
rect 49 22 57 25
rect 49 18 52 22
rect 56 18 57 22
rect 49 5 57 18
<< pdiffusion >>
rect 3 92 9 93
rect 3 88 4 92
rect 8 88 9 92
rect 39 92 47 95
rect 39 88 40 92
rect 44 88 47 92
rect 3 85 9 88
rect 39 85 47 88
rect 3 65 11 85
rect 13 65 23 85
rect 25 82 35 85
rect 25 78 28 82
rect 32 78 35 82
rect 25 72 35 78
rect 25 68 28 72
rect 32 68 35 72
rect 25 65 35 68
rect 37 65 47 85
rect 39 55 47 65
rect 49 82 57 95
rect 49 78 52 82
rect 56 78 57 82
rect 49 72 57 78
rect 49 68 52 72
rect 56 68 57 72
rect 49 62 57 68
rect 49 58 52 62
rect 56 58 57 62
rect 49 55 57 58
<< metal1 >>
rect -2 96 62 101
rect -2 92 16 96
rect 20 92 28 96
rect 32 92 62 96
rect -2 88 4 92
rect 8 88 40 92
rect 44 88 62 92
rect -2 87 62 88
rect 27 82 33 83
rect 47 82 57 83
rect 7 42 13 82
rect 7 38 8 42
rect 12 38 13 42
rect 7 37 13 38
rect 17 62 23 82
rect 27 78 28 82
rect 32 78 33 82
rect 27 77 33 78
rect 28 73 32 77
rect 27 72 33 73
rect 27 68 28 72
rect 32 68 33 72
rect 27 67 33 68
rect 17 58 18 62
rect 22 58 23 62
rect 17 42 23 58
rect 28 47 32 67
rect 37 52 43 82
rect 37 48 38 52
rect 42 48 43 52
rect 17 38 18 42
rect 22 38 23 42
rect 27 46 33 47
rect 27 42 28 46
rect 32 42 33 46
rect 27 41 33 42
rect 17 37 23 38
rect 15 32 21 33
rect 28 32 32 41
rect 15 28 16 32
rect 20 28 32 32
rect 37 32 43 48
rect 37 28 38 32
rect 42 28 43 32
rect 15 27 21 28
rect 3 22 9 23
rect 27 22 33 23
rect 3 18 4 22
rect 8 18 28 22
rect 32 18 33 22
rect 37 18 43 28
rect 47 78 52 82
rect 56 78 57 82
rect 47 77 57 78
rect 47 73 53 77
rect 47 72 57 73
rect 47 68 52 72
rect 56 68 57 72
rect 47 67 57 68
rect 47 63 53 67
rect 47 62 57 63
rect 47 58 52 62
rect 56 58 57 62
rect 47 57 57 58
rect 47 23 53 57
rect 47 22 57 23
rect 47 18 52 22
rect 56 18 57 22
rect 3 17 9 18
rect 27 17 33 18
rect 47 17 57 18
rect -2 12 62 13
rect -2 8 40 12
rect 44 8 62 12
rect -2 4 4 8
rect 8 4 16 8
rect 20 4 28 8
rect 32 4 62 8
rect -2 -1 62 4
<< ntransistor >>
rect 11 15 13 25
rect 23 15 25 25
rect 35 15 37 25
rect 47 5 49 25
<< ptransistor >>
rect 11 65 13 85
rect 23 65 25 85
rect 35 65 37 85
rect 47 55 49 95
<< polycontact >>
rect 18 58 22 62
rect 38 48 42 52
rect 8 38 12 42
rect 18 38 22 42
rect 28 42 32 46
rect 38 28 42 32
<< ndcontact >>
rect 16 28 20 32
rect 4 18 8 22
rect 28 18 32 22
rect 40 8 44 12
rect 52 18 56 22
<< pdcontact >>
rect 4 88 8 92
rect 40 88 44 92
rect 28 78 32 82
rect 28 68 32 72
rect 52 78 56 82
rect 52 68 56 72
rect 52 58 56 62
<< psubstratepcontact >>
rect 4 4 8 8
rect 16 4 20 8
rect 28 4 32 8
<< nsubstratencontact >>
rect 16 92 20 96
rect 28 92 32 96
<< psubstratepdiff >>
rect 3 8 33 9
rect 3 4 4 8
rect 8 4 16 8
rect 20 4 28 8
rect 32 4 33 8
rect 3 3 33 4
<< nsubstratendiff >>
rect 15 96 33 97
rect 15 92 16 96
rect 20 92 28 96
rect 32 92 33 96
rect 15 91 33 92
<< labels >>
rlabel metal1 10 60 10 60 6 i0
rlabel metal1 10 60 10 60 6 i0
rlabel polycontact 20 60 20 60 6 i1
rlabel polycontact 20 60 20 60 6 i1
rlabel psubstratepcontact 30 6 30 6 6 vss
rlabel psubstratepcontact 30 6 30 6 6 vss
rlabel polycontact 40 50 40 50 6 i2
rlabel polycontact 40 50 40 50 6 i2
rlabel nsubstratencontact 30 94 30 94 6 vdd
rlabel nsubstratencontact 30 94 30 94 6 vdd
rlabel metal1 50 50 50 50 6 q
rlabel metal1 50 50 50 50 6 q
<< end >>
