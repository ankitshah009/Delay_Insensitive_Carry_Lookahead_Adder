.subckt xaon22_x05 a1 a2 b1 b2 vdd vss z
*   SPICE3 file   created from xaon22_x05.ext -      technology: scmos
m00 vdd    a1     an     vdd p w=20u  l=2.3636u ad=178.5p   pd=39.5u    as=114p     ps=38.6667u
m01 an     a2     vdd    vdd p w=20u  l=2.3636u ad=114p     pd=38.6667u as=178.5p   ps=39.5u
m02 z      bn     an     vdd p w=20u  l=2.3636u ad=100p     pd=30u      as=114p     ps=38.6667u
m03 bn     an     z      vdd p w=20u  l=2.3636u ad=140.667p pd=41.3333u as=100p     ps=30u
m04 vdd    b1     bn     vdd p w=20u  l=2.3636u ad=178.5p   pd=39.5u    as=140.667p ps=41.3333u
m05 bn     b2     vdd    vdd p w=20u  l=2.3636u ad=140.667p pd=41.3333u as=178.5p   ps=39.5u
m06 w1     a1     vss    vss n w=16u  l=2.3636u ad=48p      pd=22u      as=144.39p  ps=43.7073u
m07 an     a2     w1     vss n w=16u  l=2.3636u ad=80p      pd=26u      as=48p      ps=22u
m08 w2     b2     an     vss n w=16u  l=2.3636u ad=48p      pd=22u      as=80p      ps=26u
m09 z      b1     w2     vss n w=16u  l=2.3636u ad=80p      pd=33.28u   as=48p      ps=22u
m10 w3     bn     z      vss n w=9u   l=2.3636u ad=27p      pd=15u      as=45p      ps=18.72u
m11 vss    an     w3     vss n w=9u   l=2.3636u ad=81.2195p pd=24.5854u as=27p      ps=15u
m12 w4     b1     vss    vss n w=16u  l=2.3636u ad=48p      pd=22u      as=144.39p  ps=43.7073u
m13 bn     b2     w4     vss n w=16u  l=2.3636u ad=98p      pd=48u      as=48p      ps=22u
C0  a1     vdd    0.007f
C1  vss    a2     0.007f
C2  b2     an     0.076f
C3  z      bn     0.067f
C4  b1     bn     0.279f
C5  b2     a2     0.025f
C6  z      a1     0.035f
C7  w2     z      0.005f
C8  b1     a1     0.006f
C9  an     a2     0.192f
C10 vss    z      0.040f
C11 w3     an     0.007f
C12 an     vdd    0.222f
C13 bn     a1     0.021f
C14 vss    b1     0.054f
C15 z      b2     0.015f
C16 a2     vdd    0.031f
C17 b2     b1     0.363f
C18 z      an     0.399f
C19 vss    bn     0.028f
C20 b2     bn     0.161f
C21 b1     an     0.092f
C22 z      a2     0.131f
C23 vss    a1     0.036f
C24 w4     b2     0.022f
C25 an     bn     0.478f
C26 b2     a1     0.009f
C27 z      vdd    0.015f
C28 b1     a2     0.019f
C29 an     a1     0.063f
C30 b1     vdd    0.050f
C31 bn     a2     0.069f
C32 w2     an     0.012f
C33 vss    b2     0.195f
C34 bn     vdd    0.221f
C35 a2     a1     0.148f
C36 z      b1     0.026f
C37 vss    an     0.303f
C39 z      vss    0.009f
C40 b2     vss    0.057f
C41 b1     vss    0.052f
C42 an     vss    0.039f
C43 bn     vss    0.053f
C44 a2     vss    0.038f
C45 a1     vss    0.033f
.ends
