magic
tech scmos
timestamp 1179385967
<< checkpaint >>
rect -22 -22 78 94
<< ab >>
rect 0 0 56 72
<< pwell >>
rect -4 -4 60 32
<< nwell >>
rect -4 32 60 76
<< polysilicon >>
rect 9 65 11 69
rect 19 65 21 69
rect 29 65 31 69
rect 39 57 41 61
rect 9 35 11 39
rect 19 35 21 39
rect 29 35 31 39
rect 39 35 41 39
rect 9 34 41 35
rect 9 33 28 34
rect 14 26 16 33
rect 24 30 28 33
rect 32 30 36 34
rect 40 30 41 34
rect 24 29 41 30
rect 24 26 26 29
rect 14 9 16 14
rect 24 9 26 14
<< ndiffusion >>
rect 6 19 14 26
rect 6 15 8 19
rect 12 15 14 19
rect 6 14 14 15
rect 16 25 24 26
rect 16 21 18 25
rect 22 21 24 25
rect 16 14 24 21
rect 26 19 34 26
rect 26 15 28 19
rect 32 15 34 19
rect 26 14 34 15
<< pdiffusion >>
rect 2 64 9 65
rect 2 60 3 64
rect 7 60 9 64
rect 2 57 9 60
rect 2 53 3 57
rect 7 53 9 57
rect 2 39 9 53
rect 11 51 19 65
rect 11 47 13 51
rect 17 47 19 51
rect 11 44 19 47
rect 11 40 13 44
rect 17 40 19 44
rect 11 39 19 40
rect 21 64 29 65
rect 21 60 23 64
rect 27 60 29 64
rect 21 57 29 60
rect 21 53 23 57
rect 27 53 29 57
rect 21 39 29 53
rect 31 57 36 65
rect 31 51 39 57
rect 31 47 33 51
rect 37 47 39 51
rect 31 44 39 47
rect 31 40 33 44
rect 37 40 39 44
rect 31 39 39 40
rect 41 56 48 57
rect 41 52 43 56
rect 47 52 48 56
rect 41 49 48 52
rect 41 45 43 49
rect 47 45 48 49
rect 41 39 48 45
<< metal1 >>
rect -2 68 58 72
rect -2 64 41 68
rect 45 64 48 68
rect 52 64 58 68
rect 3 57 7 60
rect 3 52 7 53
rect 23 57 27 60
rect 23 52 27 53
rect 42 56 48 64
rect 42 52 43 56
rect 47 52 48 56
rect 13 51 17 52
rect 13 44 17 47
rect 9 40 13 42
rect 33 51 39 52
rect 37 47 39 51
rect 33 44 39 47
rect 42 49 48 52
rect 42 45 43 49
rect 47 45 48 49
rect 17 40 33 42
rect 37 40 39 44
rect 9 38 39 40
rect 18 25 22 38
rect 27 30 28 34
rect 32 30 36 34
rect 40 30 47 34
rect 41 22 47 30
rect 18 20 22 21
rect 8 19 12 20
rect 8 8 12 15
rect 28 19 32 20
rect 28 8 32 15
rect -2 4 42 8
rect 46 4 58 8
rect -2 0 58 4
<< ntransistor >>
rect 14 14 16 26
rect 24 14 26 26
<< ptransistor >>
rect 9 39 11 65
rect 19 39 21 65
rect 29 39 31 65
rect 39 39 41 57
<< polycontact >>
rect 28 30 32 34
rect 36 30 40 34
<< ndcontact >>
rect 8 15 12 19
rect 18 21 22 25
rect 28 15 32 19
<< pdcontact >>
rect 3 60 7 64
rect 3 53 7 57
rect 13 47 17 51
rect 13 40 17 44
rect 23 60 27 64
rect 23 53 27 57
rect 33 47 37 51
rect 33 40 37 44
rect 43 52 47 56
rect 43 45 47 49
<< psubstratepcontact >>
rect 42 4 46 8
<< nsubstratencontact >>
rect 41 64 45 68
rect 48 64 52 68
<< psubstratepdiff >>
rect 41 8 47 24
rect 41 4 42 8
rect 46 4 47 8
rect 41 3 47 4
<< nsubstratendiff >>
rect 40 68 53 69
rect 40 64 41 68
rect 45 64 48 68
rect 52 64 53 68
rect 40 63 53 64
<< labels >>
rlabel metal1 20 32 20 32 6 z
rlabel metal1 12 40 12 40 6 z
rlabel metal1 28 4 28 4 6 vss
rlabel metal1 36 32 36 32 6 a
rlabel metal1 28 40 28 40 6 z
rlabel metal1 36 44 36 44 6 z
rlabel metal1 28 68 28 68 6 vdd
rlabel metal1 44 28 44 28 6 a
<< end >>
