magic
tech scmos
timestamp 1180600709
<< checkpaint >>
rect -22 -22 172 122
<< ab >>
rect 0 0 150 100
<< pwell >>
rect -4 -4 154 48
<< nwell >>
rect -4 48 154 104
<< polysilicon >>
rect 25 94 27 98
rect 37 94 39 98
rect 49 94 51 98
rect 57 94 59 98
rect 69 94 71 98
rect 81 94 83 98
rect 89 94 91 98
rect 113 94 115 98
rect 125 94 127 98
rect 13 70 15 74
rect 13 53 15 56
rect 5 52 15 53
rect 5 48 6 52
rect 10 48 15 52
rect 5 47 15 48
rect 13 37 15 47
rect 25 53 27 75
rect 37 73 39 76
rect 31 72 39 73
rect 31 68 32 72
rect 36 68 39 72
rect 31 67 39 68
rect 25 52 33 53
rect 25 48 28 52
rect 32 48 33 52
rect 25 47 33 48
rect 13 25 15 29
rect 25 23 27 47
rect 37 41 39 67
rect 49 63 51 75
rect 45 62 51 63
rect 45 58 46 62
rect 50 58 51 62
rect 45 57 51 58
rect 47 52 53 53
rect 47 48 48 52
rect 52 51 53 52
rect 57 51 59 75
rect 69 73 71 76
rect 81 73 83 76
rect 52 49 59 51
rect 52 48 53 49
rect 47 47 53 48
rect 37 39 51 41
rect 31 32 39 33
rect 31 28 32 32
rect 36 28 39 32
rect 31 27 39 28
rect 37 23 39 27
rect 49 23 51 39
rect 57 23 59 49
rect 67 71 71 73
rect 77 71 83 73
rect 67 33 69 71
rect 77 53 79 71
rect 89 63 91 76
rect 101 69 103 73
rect 83 62 91 63
rect 83 58 84 62
rect 88 58 91 62
rect 83 57 91 58
rect 137 76 139 80
rect 73 52 79 53
rect 73 48 74 52
rect 78 51 79 52
rect 101 51 103 55
rect 78 49 103 51
rect 78 48 79 49
rect 73 47 79 48
rect 77 39 79 47
rect 63 32 69 33
rect 63 28 64 32
rect 68 28 69 32
rect 63 27 69 28
rect 73 37 79 39
rect 83 42 91 43
rect 83 38 84 42
rect 88 38 91 42
rect 83 37 91 38
rect 101 37 103 49
rect 113 43 115 55
rect 125 43 127 55
rect 137 53 139 56
rect 131 52 139 53
rect 131 48 132 52
rect 136 51 139 52
rect 136 48 137 51
rect 131 47 137 48
rect 141 44 147 45
rect 141 43 142 44
rect 113 41 142 43
rect 73 23 75 37
rect 79 32 85 33
rect 79 28 80 32
rect 84 28 85 32
rect 79 27 85 28
rect 69 21 75 23
rect 69 18 71 21
rect 81 19 83 27
rect 89 19 91 37
rect 101 25 103 29
rect 113 27 115 41
rect 125 27 127 41
rect 141 40 142 41
rect 146 40 147 44
rect 141 39 147 40
rect 131 34 137 35
rect 131 30 132 34
rect 136 31 137 34
rect 136 30 139 31
rect 131 29 139 30
rect 25 7 27 11
rect 37 7 39 11
rect 49 7 51 11
rect 57 7 59 11
rect 137 26 139 29
rect 137 12 139 16
rect 69 2 71 6
rect 81 3 83 7
rect 89 3 91 7
rect 113 3 115 7
rect 125 3 127 7
<< ndiffusion >>
rect 5 29 13 37
rect 15 34 23 37
rect 15 30 18 34
rect 22 30 23 34
rect 15 29 23 30
rect 5 22 11 29
rect 41 32 47 33
rect 41 28 42 32
rect 46 28 47 32
rect 41 23 47 28
rect 5 18 6 22
rect 10 18 11 22
rect 5 17 11 18
rect 17 22 25 23
rect 17 18 18 22
rect 22 18 25 22
rect 17 11 25 18
rect 27 11 37 23
rect 39 11 49 23
rect 51 11 57 23
rect 59 22 67 23
rect 59 18 62 22
rect 66 18 67 22
rect 93 36 101 37
rect 93 32 94 36
rect 98 32 101 36
rect 93 29 101 32
rect 103 29 111 37
rect 105 27 111 29
rect 117 32 123 33
rect 117 28 118 32
rect 122 28 123 32
rect 117 27 123 28
rect 93 22 99 23
rect 93 19 94 22
rect 76 18 81 19
rect 59 11 69 18
rect 61 6 69 11
rect 71 12 81 18
rect 71 8 74 12
rect 78 8 81 12
rect 71 7 81 8
rect 83 7 89 19
rect 91 18 94 19
rect 98 18 99 22
rect 91 7 99 18
rect 105 12 113 27
rect 105 8 106 12
rect 110 8 113 12
rect 105 7 113 8
rect 115 7 125 27
rect 127 26 132 27
rect 127 16 137 26
rect 139 24 147 26
rect 139 20 142 24
rect 146 20 147 24
rect 139 16 147 20
rect 127 12 135 16
rect 127 8 130 12
rect 134 8 135 12
rect 127 7 135 8
rect 71 6 78 7
<< pdiffusion >>
rect 105 94 111 95
rect 129 94 135 95
rect 5 82 11 83
rect 5 78 6 82
rect 10 78 11 82
rect 5 70 11 78
rect 17 82 25 94
rect 17 78 18 82
rect 22 78 25 82
rect 17 75 25 78
rect 27 76 37 94
rect 39 76 49 94
rect 27 75 32 76
rect 5 56 13 70
rect 15 62 23 70
rect 15 58 18 62
rect 22 58 23 62
rect 15 56 23 58
rect 41 75 49 76
rect 51 75 57 94
rect 59 82 69 94
rect 59 78 62 82
rect 66 78 69 82
rect 59 76 69 78
rect 71 92 81 94
rect 71 88 74 92
rect 78 88 81 92
rect 71 76 81 88
rect 83 76 89 94
rect 91 82 99 94
rect 91 78 94 82
rect 98 78 99 82
rect 91 76 99 78
rect 105 90 106 94
rect 110 90 113 94
rect 59 75 64 76
rect 41 72 47 75
rect 41 68 42 72
rect 46 68 47 72
rect 41 67 47 68
rect 105 69 113 90
rect 93 62 101 69
rect 93 58 94 62
rect 98 58 101 62
rect 93 55 101 58
rect 103 55 113 69
rect 115 82 125 94
rect 115 78 118 82
rect 122 78 125 82
rect 115 72 125 78
rect 115 68 118 72
rect 122 68 125 72
rect 115 62 125 68
rect 115 58 118 62
rect 122 58 125 62
rect 115 55 125 58
rect 127 90 130 94
rect 134 90 135 94
rect 127 82 135 90
rect 127 78 130 82
rect 134 78 135 82
rect 127 76 135 78
rect 127 72 137 76
rect 127 68 130 72
rect 134 68 137 72
rect 127 62 137 68
rect 127 58 130 62
rect 134 58 137 62
rect 127 56 137 58
rect 139 72 147 76
rect 139 68 142 72
rect 146 68 147 72
rect 139 62 147 68
rect 139 58 142 62
rect 146 58 147 62
rect 139 56 147 58
rect 127 55 132 56
<< metal1 >>
rect -2 96 152 100
rect -2 94 142 96
rect -2 92 106 94
rect -2 88 74 92
rect 78 90 106 92
rect 110 90 130 94
rect 134 92 142 94
rect 146 92 152 96
rect 134 90 152 92
rect 78 88 152 90
rect 6 82 10 88
rect 94 82 98 83
rect 17 78 18 82
rect 22 78 62 82
rect 66 78 67 82
rect 6 77 10 78
rect 8 72 12 73
rect 94 72 98 78
rect 118 82 122 83
rect 118 72 122 78
rect 8 68 32 72
rect 36 68 37 72
rect 41 68 42 72
rect 46 68 112 72
rect 8 52 12 68
rect 5 48 6 52
rect 10 48 12 52
rect 8 27 12 48
rect 18 62 22 63
rect 22 58 46 62
rect 50 58 51 62
rect 18 34 22 58
rect 28 52 32 53
rect 39 48 48 52
rect 52 48 53 52
rect 28 41 32 48
rect 58 42 62 68
rect 52 38 62 42
rect 68 52 72 63
rect 84 62 88 63
rect 77 58 84 62
rect 93 58 94 62
rect 84 52 88 58
rect 68 48 74 52
rect 78 48 79 52
rect 84 48 93 52
rect 52 32 56 38
rect 68 37 72 48
rect 84 42 88 48
rect 77 38 84 42
rect 84 37 88 38
rect 98 37 102 62
rect 94 36 102 37
rect 98 33 102 36
rect 22 30 32 32
rect 18 28 32 30
rect 36 28 37 32
rect 41 28 42 32
rect 46 28 56 32
rect 63 28 64 32
rect 68 28 80 32
rect 84 28 98 32
rect 6 22 10 23
rect 108 22 112 68
rect 118 62 122 68
rect 118 32 122 58
rect 130 82 134 88
rect 130 72 134 78
rect 130 62 134 68
rect 130 57 134 58
rect 142 72 146 73
rect 142 62 146 68
rect 118 27 122 28
rect 132 52 136 53
rect 132 34 136 48
rect 132 22 136 30
rect 17 18 18 22
rect 22 18 62 22
rect 66 18 67 22
rect 93 18 94 22
rect 98 18 136 22
rect 142 44 146 58
rect 142 24 146 40
rect 142 19 146 20
rect 6 12 10 18
rect -2 8 74 12
rect 78 8 106 12
rect 110 8 130 12
rect 134 8 152 12
rect -2 0 152 8
<< ntransistor >>
rect 13 29 15 37
rect 25 11 27 23
rect 37 11 39 23
rect 49 11 51 23
rect 57 11 59 23
rect 101 29 103 37
rect 69 6 71 18
rect 81 7 83 19
rect 89 7 91 19
rect 113 7 115 27
rect 125 7 127 27
rect 137 16 139 26
<< ptransistor >>
rect 25 75 27 94
rect 37 76 39 94
rect 13 56 15 70
rect 49 75 51 94
rect 57 75 59 94
rect 69 76 71 94
rect 81 76 83 94
rect 89 76 91 94
rect 101 55 103 69
rect 113 55 115 94
rect 125 55 127 94
rect 137 56 139 76
<< polycontact >>
rect 6 48 10 52
rect 32 68 36 72
rect 28 48 32 52
rect 46 58 50 62
rect 48 48 52 52
rect 32 28 36 32
rect 84 58 88 62
rect 74 48 78 52
rect 64 28 68 32
rect 84 38 88 42
rect 132 48 136 52
rect 80 28 84 32
rect 142 40 146 44
rect 132 30 136 34
<< ndcontact >>
rect 18 30 22 34
rect 42 28 46 32
rect 6 18 10 22
rect 18 18 22 22
rect 62 18 66 22
rect 94 32 98 36
rect 118 28 122 32
rect 74 8 78 12
rect 94 18 98 22
rect 106 8 110 12
rect 142 20 146 24
rect 130 8 134 12
<< pdcontact >>
rect 6 78 10 82
rect 18 78 22 82
rect 18 58 22 62
rect 62 78 66 82
rect 74 88 78 92
rect 94 78 98 82
rect 106 90 110 94
rect 42 68 46 72
rect 94 58 98 62
rect 118 78 122 82
rect 118 68 122 72
rect 118 58 122 62
rect 130 90 134 94
rect 130 78 134 82
rect 130 68 134 72
rect 130 58 134 62
rect 142 68 146 72
rect 142 58 146 62
<< nsubstratencontact >>
rect 142 92 146 96
<< nsubstratendiff >>
rect 141 96 147 97
rect 141 92 142 96
rect 146 92 147 96
rect 141 86 147 92
<< labels >>
rlabel metal1 10 50 10 50 6 cmd1
rlabel metal1 20 70 20 70 6 cmd1
rlabel polycontact 30 50 30 50 6 i2
rlabel polycontact 50 50 50 50 6 i1
rlabel metal1 30 70 30 70 6 cmd1
rlabel metal1 75 6 75 6 6 vss
rlabel metal1 80 40 80 40 6 i0
rlabel metal1 70 50 70 50 6 cmd0
rlabel metal1 80 60 80 60 6 i0
rlabel metal1 75 94 75 94 6 vdd
rlabel metal1 90 50 90 50 6 i0
rlabel metal1 120 55 120 55 6 nq
<< end >>
