magic
tech scmos
timestamp 1179387446
<< checkpaint >>
rect -22 -25 166 105
<< ab >>
rect 0 0 144 80
<< pwell >>
rect -4 -7 148 36
<< nwell >>
rect -4 36 148 87
<< polysilicon >>
rect 18 69 20 74
rect 28 69 30 74
rect 38 72 50 74
rect 38 69 40 72
rect 48 69 50 72
rect 69 70 71 74
rect 79 70 81 74
rect 91 70 93 74
rect 101 70 103 74
rect 118 70 120 74
rect 128 70 130 74
rect 2 40 8 41
rect 2 36 3 40
rect 7 37 8 40
rect 18 39 20 42
rect 28 39 30 42
rect 38 39 40 42
rect 16 38 31 39
rect 16 37 26 38
rect 7 36 11 37
rect 2 35 11 36
rect 9 30 11 35
rect 16 30 18 37
rect 25 34 26 37
rect 30 34 31 38
rect 25 33 31 34
rect 35 38 41 39
rect 48 38 50 42
rect 69 39 71 42
rect 79 39 81 42
rect 91 39 93 42
rect 101 39 103 42
rect 69 38 87 39
rect 35 34 36 38
rect 40 34 41 38
rect 69 37 82 38
rect 35 33 41 34
rect 28 30 30 33
rect 35 30 37 33
rect 45 30 47 34
rect 55 30 57 35
rect 81 34 82 37
rect 86 34 87 38
rect 81 33 87 34
rect 91 38 104 39
rect 91 34 98 38
rect 102 34 104 38
rect 91 33 104 34
rect 108 38 114 39
rect 108 34 109 38
rect 113 34 114 38
rect 118 38 120 42
rect 128 39 130 42
rect 128 38 135 39
rect 118 35 121 38
rect 108 33 114 34
rect 85 30 87 33
rect 92 30 94 33
rect 102 30 104 33
rect 109 30 111 33
rect 119 30 121 35
rect 128 34 130 38
rect 134 34 135 38
rect 128 33 135 34
rect 129 30 131 33
rect 9 18 11 23
rect 16 18 18 23
rect 85 12 87 16
rect 92 12 94 16
rect 102 12 104 16
rect 109 12 111 16
rect 28 6 30 11
rect 35 6 37 11
rect 45 8 47 11
rect 55 8 57 11
rect 119 8 121 16
rect 129 8 131 16
rect 45 6 131 8
<< ndiffusion >>
rect 2 29 9 30
rect 2 25 3 29
rect 7 25 9 29
rect 2 23 9 25
rect 11 23 16 30
rect 18 23 28 30
rect 20 14 28 23
rect 20 10 21 14
rect 25 11 28 14
rect 30 11 35 30
rect 37 22 45 30
rect 37 18 39 22
rect 43 18 45 22
rect 37 11 45 18
rect 47 29 55 30
rect 47 25 49 29
rect 53 25 55 29
rect 47 11 55 25
rect 57 23 62 30
rect 57 22 64 23
rect 57 18 59 22
rect 63 18 64 22
rect 57 17 64 18
rect 78 21 85 30
rect 78 17 79 21
rect 83 17 85 21
rect 57 11 62 17
rect 78 16 85 17
rect 87 16 92 30
rect 94 21 102 30
rect 94 17 96 21
rect 100 17 102 21
rect 94 16 102 17
rect 104 16 109 30
rect 111 21 119 30
rect 111 17 113 21
rect 117 17 119 21
rect 111 16 119 17
rect 121 28 129 30
rect 121 24 123 28
rect 127 24 129 28
rect 121 21 129 24
rect 121 17 123 21
rect 127 17 129 21
rect 121 16 129 17
rect 131 28 138 30
rect 131 24 133 28
rect 137 24 138 28
rect 131 21 138 24
rect 131 17 133 21
rect 137 17 138 21
rect 131 16 138 17
rect 25 10 26 11
rect 20 9 26 10
<< pdiffusion >>
rect 62 69 69 70
rect 13 55 18 69
rect 11 54 18 55
rect 11 50 12 54
rect 16 50 18 54
rect 11 47 18 50
rect 11 43 12 47
rect 16 43 18 47
rect 11 42 18 43
rect 20 62 28 69
rect 20 58 22 62
rect 26 58 28 62
rect 20 42 28 58
rect 30 54 38 69
rect 30 50 32 54
rect 36 50 38 54
rect 30 42 38 50
rect 40 47 48 69
rect 40 43 42 47
rect 46 43 48 47
rect 40 42 48 43
rect 50 55 55 69
rect 62 65 63 69
rect 67 65 69 69
rect 50 54 57 55
rect 50 50 52 54
rect 56 50 57 54
rect 50 47 57 50
rect 50 43 52 47
rect 56 43 57 47
rect 50 42 57 43
rect 62 42 69 65
rect 71 54 79 70
rect 71 50 73 54
rect 77 50 79 54
rect 71 47 79 50
rect 71 43 73 47
rect 77 43 79 47
rect 71 42 79 43
rect 81 69 91 70
rect 81 65 84 69
rect 88 65 91 69
rect 81 42 91 65
rect 93 54 101 70
rect 93 50 95 54
rect 99 50 101 54
rect 93 42 101 50
rect 103 69 118 70
rect 103 65 105 69
rect 109 65 112 69
rect 116 65 118 69
rect 103 62 118 65
rect 103 58 112 62
rect 116 58 118 62
rect 103 42 118 58
rect 120 47 128 70
rect 120 43 122 47
rect 126 43 128 47
rect 120 42 128 43
rect 130 69 138 70
rect 130 65 133 69
rect 137 65 138 69
rect 130 42 138 65
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect 118 78 122 82
rect 126 78 130 82
rect 134 78 138 82
rect 142 78 146 82
rect -2 69 146 78
rect -2 68 63 69
rect 62 65 63 68
rect 67 68 84 69
rect 67 65 68 68
rect 83 65 84 68
rect 88 68 105 69
rect 88 65 89 68
rect 103 65 105 68
rect 109 65 112 69
rect 116 68 133 69
rect 116 65 117 68
rect 132 65 133 68
rect 137 68 146 69
rect 137 65 138 68
rect 111 62 117 65
rect 3 58 22 62
rect 26 58 107 62
rect 111 58 112 62
rect 116 58 117 62
rect 121 58 134 62
rect 3 40 7 58
rect 3 35 7 36
rect 10 50 12 54
rect 16 50 32 54
rect 36 50 52 54
rect 56 50 57 54
rect 10 47 16 50
rect 52 47 57 50
rect 10 43 12 47
rect 10 42 16 43
rect 26 43 42 47
rect 46 43 47 47
rect 56 43 57 47
rect 10 31 14 42
rect 2 29 14 31
rect 2 25 3 29
rect 7 25 14 29
rect 26 38 30 43
rect 52 42 57 43
rect 60 38 64 58
rect 103 54 107 58
rect 35 34 36 38
rect 40 34 64 38
rect 72 50 73 54
rect 77 50 95 54
rect 99 50 100 54
rect 103 50 126 54
rect 72 47 77 50
rect 72 43 73 47
rect 122 47 126 50
rect 26 29 30 34
rect 72 29 77 43
rect 81 42 119 46
rect 81 38 87 42
rect 108 38 114 42
rect 81 34 82 38
rect 86 34 87 38
rect 97 34 98 38
rect 102 34 103 38
rect 108 34 109 38
rect 113 34 114 38
rect 97 30 103 34
rect 26 25 49 29
rect 53 25 92 29
rect 97 26 111 30
rect 122 29 126 43
rect 130 38 134 58
rect 130 33 134 34
rect 122 28 127 29
rect 10 22 14 25
rect 10 18 39 22
rect 43 18 59 22
rect 63 18 64 22
rect 88 21 92 25
rect 122 24 123 28
rect 113 21 117 22
rect 78 17 79 21
rect 83 17 84 21
rect 88 17 96 21
rect 100 17 101 21
rect 20 12 21 14
rect -2 10 21 12
rect 25 12 26 14
rect 69 12 73 16
rect 78 12 84 17
rect 113 12 117 17
rect 122 21 127 24
rect 122 17 123 21
rect 122 16 127 17
rect 133 28 137 29
rect 133 21 137 24
rect 133 12 137 17
rect 25 10 146 12
rect -2 2 146 10
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 122 2
rect 126 -2 130 2
rect 134 -2 138 2
rect 142 -2 146 2
<< ntransistor >>
rect 9 23 11 30
rect 16 23 18 30
rect 28 11 30 30
rect 35 11 37 30
rect 45 11 47 30
rect 55 11 57 30
rect 85 16 87 30
rect 92 16 94 30
rect 102 16 104 30
rect 109 16 111 30
rect 119 16 121 30
rect 129 16 131 30
<< ptransistor >>
rect 18 42 20 69
rect 28 42 30 69
rect 38 42 40 69
rect 48 42 50 69
rect 69 42 71 70
rect 79 42 81 70
rect 91 42 93 70
rect 101 42 103 70
rect 118 42 120 70
rect 128 42 130 70
<< polycontact >>
rect 3 36 7 40
rect 26 34 30 38
rect 36 34 40 38
rect 82 34 86 38
rect 98 34 102 38
rect 109 34 113 38
rect 130 34 134 38
<< ndcontact >>
rect 3 25 7 29
rect 21 10 25 14
rect 39 18 43 22
rect 49 25 53 29
rect 59 18 63 22
rect 79 17 83 21
rect 96 17 100 21
rect 113 17 117 21
rect 123 24 127 28
rect 123 17 127 21
rect 133 24 137 28
rect 133 17 137 21
<< pdcontact >>
rect 12 50 16 54
rect 12 43 16 47
rect 22 58 26 62
rect 32 50 36 54
rect 42 43 46 47
rect 63 65 67 69
rect 52 50 56 54
rect 52 43 56 47
rect 73 50 77 54
rect 73 43 77 47
rect 84 65 88 69
rect 95 50 99 54
rect 105 65 109 69
rect 112 65 116 69
rect 112 58 116 62
rect 122 43 126 47
rect 133 65 137 69
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
rect 90 -2 94 2
rect 98 -2 102 2
rect 106 -2 110 2
rect 114 -2 118 2
rect 122 -2 126 2
rect 130 -2 134 2
rect 138 -2 142 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
rect 90 78 94 82
rect 98 78 102 82
rect 106 78 110 82
rect 114 78 118 82
rect 122 78 126 82
rect 130 78 134 82
rect 138 78 142 82
<< psubstratepdiff >>
rect 0 2 144 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 122 2
rect 126 -2 130 2
rect 134 -2 138 2
rect 142 -2 144 2
rect 0 -3 144 -2
<< nsubstratendiff >>
rect 0 82 144 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect 118 78 122 82
rect 126 78 130 82
rect 134 78 138 82
rect 142 78 144 82
rect 0 77 144 78
<< labels >>
rlabel polycontact 5 38 5 38 6 bn
rlabel polysilicon 29 40 29 40 6 an
rlabel ptransistor 39 53 39 53 6 bn
rlabel metal1 20 20 20 20 6 z
rlabel ndcontact 4 28 4 28 6 z
rlabel metal1 12 36 12 36 6 z
rlabel metal1 20 52 20 52 6 z
rlabel metal1 5 48 5 48 6 bn
rlabel metal1 28 20 28 20 6 z
rlabel metal1 36 20 36 20 6 z
rlabel metal1 44 20 44 20 6 z
rlabel metal1 52 20 52 20 6 z
rlabel polycontact 28 36 28 36 6 an
rlabel metal1 36 45 36 45 6 an
rlabel metal1 36 52 36 52 6 z
rlabel metal1 44 52 44 52 6 z
rlabel metal1 52 52 52 52 6 z
rlabel metal1 28 52 28 52 6 z
rlabel metal1 72 6 72 6 6 vss
rlabel ndcontact 60 20 60 20 6 z
rlabel metal1 49 36 49 36 6 bn
rlabel metal1 84 40 84 40 6 a2
rlabel metal1 74 39 74 39 6 an
rlabel metal1 72 74 72 74 6 vdd
rlabel metal1 94 19 94 19 6 an
rlabel metal1 59 27 59 27 6 an
rlabel metal1 108 28 108 28 6 a1
rlabel metal1 100 32 100 32 6 a1
rlabel metal1 100 44 100 44 6 a2
rlabel metal1 108 44 108 44 6 a2
rlabel metal1 92 44 92 44 6 a2
rlabel metal1 86 52 86 52 6 an
rlabel metal1 55 60 55 60 6 bn
rlabel metal1 116 44 116 44 6 a2
rlabel metal1 132 44 132 44 6 b
rlabel metal1 124 35 124 35 6 bn
rlabel metal1 124 60 124 60 6 b
<< end >>
