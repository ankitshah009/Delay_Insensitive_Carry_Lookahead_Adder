magic
tech scmos
timestamp 1179385766
<< checkpaint >>
rect -22 -22 86 94
<< ab >>
rect 0 0 64 72
<< pwell >>
rect -4 -4 68 32
<< nwell >>
rect -4 32 68 76
<< polysilicon >>
rect 9 51 11 61
rect 19 60 21 70
rect 39 60 41 70
rect 49 60 51 65
rect 19 59 28 60
rect 19 55 23 59
rect 27 55 28 59
rect 19 54 28 55
rect 19 51 21 54
rect 39 40 41 54
rect 49 50 51 54
rect 45 49 51 50
rect 45 45 46 49
rect 50 45 51 49
rect 45 44 51 45
rect 9 34 11 39
rect 19 34 21 39
rect 9 33 15 34
rect 9 29 10 33
rect 14 29 15 33
rect 9 28 15 29
rect 19 33 35 34
rect 19 29 30 33
rect 34 29 35 33
rect 19 28 35 29
rect 39 33 45 40
rect 39 29 40 33
rect 44 29 45 33
rect 9 24 11 28
rect 19 24 21 28
rect 39 27 45 29
rect 39 24 41 27
rect 49 24 51 44
rect 9 2 11 18
rect 19 2 21 18
rect 39 2 41 18
rect 49 13 51 18
<< ndiffusion >>
rect 2 23 9 24
rect 2 19 3 23
rect 7 19 9 23
rect 2 18 9 19
rect 11 23 19 24
rect 11 19 13 23
rect 17 19 19 23
rect 11 18 19 19
rect 21 23 28 24
rect 21 19 23 23
rect 27 19 28 23
rect 21 18 28 19
rect 32 23 39 24
rect 32 19 33 23
rect 37 19 39 23
rect 32 18 39 19
rect 41 23 49 24
rect 41 19 43 23
rect 47 19 49 23
rect 41 18 49 19
rect 51 23 58 24
rect 51 19 53 23
rect 57 19 58 23
rect 51 18 58 19
<< pdiffusion >>
rect 32 59 39 60
rect 32 55 33 59
rect 37 55 39 59
rect 32 54 39 55
rect 41 59 49 60
rect 41 55 43 59
rect 47 55 49 59
rect 41 54 49 55
rect 51 59 58 60
rect 51 55 53 59
rect 57 55 58 59
rect 51 54 58 55
rect 2 50 9 51
rect 2 46 3 50
rect 7 46 9 50
rect 2 39 9 46
rect 11 50 19 51
rect 11 46 13 50
rect 17 46 19 50
rect 11 39 19 46
rect 21 50 28 51
rect 21 46 23 50
rect 27 46 28 50
rect 21 39 28 46
<< metal1 >>
rect -2 68 66 72
rect -2 64 4 68
rect 8 64 12 68
rect 16 64 66 68
rect 2 50 8 59
rect 2 46 3 50
rect 7 46 8 50
rect 12 50 18 64
rect 42 59 48 64
rect 22 55 23 59
rect 27 55 33 59
rect 37 55 38 59
rect 42 55 43 59
rect 47 55 48 59
rect 42 54 48 55
rect 52 59 58 60
rect 52 55 53 59
rect 57 55 58 59
rect 52 54 58 55
rect 12 46 13 50
rect 17 46 18 50
rect 22 50 28 51
rect 22 46 23 50
rect 27 46 28 50
rect 2 42 8 46
rect 2 38 18 42
rect 22 38 28 46
rect 33 49 50 50
rect 33 45 46 49
rect 33 44 50 45
rect 2 24 6 38
rect 22 34 26 38
rect 32 34 36 40
rect 41 38 47 44
rect 54 34 58 54
rect 10 33 26 34
rect 14 29 26 33
rect 10 28 26 29
rect 30 33 36 34
rect 34 29 36 33
rect 30 28 36 29
rect 40 33 58 34
rect 44 29 58 33
rect 40 28 58 29
rect 22 24 26 28
rect 32 24 36 28
rect 2 23 8 24
rect 2 19 3 23
rect 7 19 8 23
rect 2 13 8 19
rect 12 23 18 24
rect 12 19 13 23
rect 17 19 18 23
rect 12 8 18 19
rect 22 23 28 24
rect 22 19 23 23
rect 27 19 28 23
rect 22 13 28 19
rect 32 23 38 24
rect 32 19 33 23
rect 37 19 38 23
rect 32 13 38 19
rect 42 23 48 24
rect 42 19 43 23
rect 47 19 48 23
rect 42 8 48 19
rect 52 23 58 28
rect 52 19 53 23
rect 57 19 58 23
rect 52 13 58 19
rect -2 4 24 8
rect 28 4 32 8
rect 36 4 66 8
rect -2 0 66 4
<< ntransistor >>
rect 9 18 11 24
rect 19 18 21 24
rect 39 18 41 24
rect 49 18 51 24
<< ptransistor >>
rect 39 54 41 60
rect 49 54 51 60
rect 9 39 11 51
rect 19 39 21 51
<< polycontact >>
rect 23 55 27 59
rect 46 45 50 49
rect 10 29 14 33
rect 30 29 34 33
rect 40 29 44 33
<< ndcontact >>
rect 3 19 7 23
rect 13 19 17 23
rect 23 19 27 23
rect 33 19 37 23
rect 43 19 47 23
rect 53 19 57 23
<< pdcontact >>
rect 33 55 37 59
rect 43 55 47 59
rect 53 55 57 59
rect 3 46 7 50
rect 13 46 17 50
rect 23 46 27 50
<< psubstratepcontact >>
rect 24 4 28 8
rect 32 4 36 8
<< nsubstratencontact >>
rect 4 64 8 68
rect 12 64 16 68
<< psubstratepdiff >>
rect 23 8 37 9
rect 23 4 24 8
rect 28 4 32 8
rect 36 4 37 8
rect 23 3 37 4
<< nsubstratendiff >>
rect 3 68 17 69
rect 3 64 4 68
rect 8 64 12 68
rect 16 64 17 68
rect 3 63 17 64
<< labels >>
rlabel polycontact 12 31 12 31 6 n3
rlabel polysilicon 27 31 27 31 6 n2
rlabel polysilicon 23 57 23 57 6 n2
rlabel polysilicon 42 33 42 33 6 n1
rlabel metal1 12 40 12 40 6 z
rlabel metal1 4 36 4 36 6 z
rlabel metal1 18 31 18 31 6 n3
rlabel metal1 25 44 25 44 6 n3
rlabel metal1 32 4 32 4 6 vss
rlabel metal1 36 48 36 48 6 a
rlabel metal1 44 44 44 44 6 a
rlabel metal1 30 57 30 57 6 n2
rlabel metal1 32 68 32 68 6 vdd
rlabel metal1 49 31 49 31 6 n1
<< end >>
