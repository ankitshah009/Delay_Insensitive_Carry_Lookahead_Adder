.subckt bf1v0x6 a vdd vss z
*   SPICE3 file   created from bf1v0x6.ext -      technology: scmos
m00 vdd    an     z      vdd p w=27u  l=2.3636u ad=124.615p pd=43.8462u as=125.667p ps=46u
m01 z      an     vdd    vdd p w=27u  l=2.3636u ad=125.667p pd=46u      as=124.615p ps=43.8462u
m02 vdd    an     z      vdd p w=27u  l=2.3636u ad=124.615p pd=43.8462u as=125.667p ps=46u
m03 an     a      vdd    vdd p w=18u  l=2.3636u ad=72p      pd=26u      as=83.0769p ps=29.2308u
m04 vdd    a      an     vdd p w=18u  l=2.3636u ad=83.0769p pd=29.2308u as=72p      ps=26u
m05 z      an     vss    vss n w=20u  l=2.3636u ad=80p      pd=28u      as=128.136p ps=40u
m06 vss    an     z      vss n w=20u  l=2.3636u ad=128.136p pd=40u      as=80p      ps=28u
m07 an     a      vss    vss n w=19u  l=2.3636u ad=121p     pd=52u      as=121.729p ps=38u
C0  vss    z      0.166f
C1  a      an     0.217f
C2  vss    vdd    0.010f
C3  z      vdd    0.109f
C4  vss    a      0.028f
C5  vss    an     0.128f
C6  a      z      0.013f
C7  z      an     0.137f
C8  a      vdd    0.020f
C9  an     vdd    0.121f
C11 a      vss    0.034f
C12 z      vss    0.006f
C13 an     vss    0.046f
.ends
