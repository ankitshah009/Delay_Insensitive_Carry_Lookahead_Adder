magic
tech scmos
timestamp 1179385884
<< checkpaint >>
rect -22 -22 54 94
<< ab >>
rect 0 0 32 72
<< pwell >>
rect -4 -4 36 32
<< nwell >>
rect -4 32 36 76
<< polysilicon >>
rect 9 66 11 70
rect 19 66 21 70
rect 9 35 11 38
rect 19 35 21 38
rect 9 34 21 35
rect 9 30 16 34
rect 20 30 21 34
rect 9 29 21 30
rect 9 26 11 29
rect 19 26 21 29
rect 9 2 11 7
rect 19 2 21 7
<< ndiffusion >>
rect 2 19 9 26
rect 2 15 3 19
rect 7 15 9 19
rect 2 12 9 15
rect 2 8 3 12
rect 7 8 9 12
rect 2 7 9 8
rect 11 25 19 26
rect 11 21 13 25
rect 17 21 19 25
rect 11 18 19 21
rect 11 14 13 18
rect 17 14 19 18
rect 11 7 19 14
rect 21 19 29 26
rect 21 15 23 19
rect 27 15 29 19
rect 21 12 29 15
rect 21 8 23 12
rect 27 8 29 12
rect 21 7 29 8
<< pdiffusion >>
rect 2 65 9 66
rect 2 61 3 65
rect 7 61 9 65
rect 2 58 9 61
rect 2 54 3 58
rect 7 54 9 58
rect 2 38 9 54
rect 11 58 19 66
rect 11 54 13 58
rect 17 54 19 58
rect 11 51 19 54
rect 11 47 13 51
rect 17 47 19 51
rect 11 38 19 47
rect 21 65 29 66
rect 21 61 23 65
rect 27 61 29 65
rect 21 58 29 61
rect 21 54 23 58
rect 27 54 29 58
rect 21 38 29 54
<< metal1 >>
rect -2 65 34 72
rect -2 64 3 65
rect 2 61 3 64
rect 7 64 23 65
rect 7 61 8 64
rect 2 58 8 61
rect 22 61 23 64
rect 27 64 34 65
rect 27 61 28 64
rect 2 54 3 58
rect 7 54 8 58
rect 13 58 17 59
rect 22 58 28 61
rect 22 54 23 58
rect 27 54 28 58
rect 13 51 17 54
rect 2 47 13 50
rect 2 46 17 47
rect 2 26 6 46
rect 26 34 30 43
rect 15 30 16 34
rect 20 30 30 34
rect 2 25 23 26
rect 2 22 13 25
rect 17 22 23 25
rect 2 15 3 19
rect 7 15 8 19
rect 2 12 8 15
rect 13 18 17 21
rect 13 13 17 14
rect 22 15 23 19
rect 27 15 28 19
rect 2 8 3 12
rect 7 8 8 12
rect 22 12 28 15
rect 22 8 23 12
rect 27 8 28 12
rect -2 0 34 8
<< ntransistor >>
rect 9 7 11 26
rect 19 7 21 26
<< ptransistor >>
rect 9 38 11 66
rect 19 38 21 66
<< polycontact >>
rect 16 30 20 34
<< ndcontact >>
rect 3 15 7 19
rect 3 8 7 12
rect 13 21 17 25
rect 13 14 17 18
rect 23 15 27 19
rect 23 8 27 12
<< pdcontact >>
rect 3 61 7 65
rect 3 54 7 58
rect 13 54 17 58
rect 13 47 17 51
rect 23 61 27 65
rect 23 54 27 58
<< labels >>
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 24 12 24 6 z
rlabel metal1 12 48 12 48 6 z
rlabel metal1 16 4 16 4 6 vss
rlabel metal1 20 32 20 32 6 a
rlabel metal1 20 24 20 24 6 z
rlabel metal1 16 68 16 68 6 vdd
rlabel metal1 28 40 28 40 6 a
<< end >>
