magic
tech scmos
timestamp 1185038947
<< checkpaint >>
rect -22 -24 72 124
<< ab >>
rect 0 0 50 100
<< pwell >>
rect -2 -4 52 49
<< nwell >>
rect -2 49 52 104
<< polysilicon >>
rect 23 95 25 98
rect 35 95 37 98
rect 11 75 13 78
rect 11 53 13 55
rect 11 52 19 53
rect 11 48 14 52
rect 18 48 19 52
rect 11 47 19 48
rect 23 43 25 55
rect 35 43 37 55
rect 3 42 37 43
rect 3 38 4 42
rect 8 38 37 42
rect 3 37 37 38
rect 11 32 19 33
rect 11 28 14 32
rect 18 28 19 32
rect 11 27 19 28
rect 11 25 13 27
rect 23 25 25 37
rect 35 25 37 37
rect 11 12 13 15
rect 23 2 25 5
rect 35 2 37 5
<< ndiffusion >>
rect 3 22 11 25
rect 3 18 4 22
rect 8 18 11 22
rect 3 15 11 18
rect 13 15 23 25
rect 15 12 23 15
rect 15 8 16 12
rect 20 8 23 12
rect 15 5 23 8
rect 25 22 35 25
rect 25 18 28 22
rect 32 18 35 22
rect 25 5 35 18
rect 37 22 45 25
rect 37 18 40 22
rect 44 18 45 22
rect 37 12 45 18
rect 37 8 40 12
rect 44 8 45 12
rect 37 5 45 8
<< pdiffusion >>
rect 15 92 23 95
rect 15 88 16 92
rect 20 88 23 92
rect 15 75 23 88
rect 3 72 11 75
rect 3 68 4 72
rect 8 68 11 72
rect 3 62 11 68
rect 3 58 4 62
rect 8 58 11 62
rect 3 55 11 58
rect 13 55 23 75
rect 25 82 35 95
rect 25 78 28 82
rect 32 78 35 82
rect 25 72 35 78
rect 25 68 28 72
rect 32 68 35 72
rect 25 62 35 68
rect 25 58 28 62
rect 32 58 35 62
rect 25 55 35 58
rect 37 92 45 95
rect 37 88 40 92
rect 44 88 45 92
rect 37 82 45 88
rect 37 78 40 82
rect 44 78 45 82
rect 37 72 45 78
rect 37 68 40 72
rect 44 68 45 72
rect 37 62 45 68
rect 37 58 40 62
rect 44 58 45 62
rect 37 55 45 58
<< metal1 >>
rect -2 96 52 101
rect -2 92 4 96
rect 8 92 52 96
rect -2 88 16 92
rect 20 88 40 92
rect 44 88 52 92
rect -2 87 52 88
rect 3 86 9 87
rect 3 82 4 86
rect 8 82 9 86
rect 27 82 33 83
rect 3 81 9 82
rect 3 72 9 73
rect 3 68 4 72
rect 8 68 9 72
rect 3 67 9 68
rect 4 63 8 67
rect 3 62 9 63
rect 3 58 4 62
rect 8 58 9 62
rect 3 57 9 58
rect 4 43 8 57
rect 17 53 23 82
rect 13 52 23 53
rect 13 48 14 52
rect 18 48 23 52
rect 13 47 23 48
rect 3 42 9 43
rect 3 38 4 42
rect 8 38 9 42
rect 3 37 9 38
rect 4 23 8 37
rect 17 33 23 47
rect 13 32 23 33
rect 13 28 14 32
rect 18 28 23 32
rect 13 27 23 28
rect 3 22 9 23
rect 3 18 4 22
rect 8 18 9 22
rect 17 18 23 27
rect 27 78 28 82
rect 32 78 33 82
rect 27 72 33 78
rect 27 68 28 72
rect 32 68 33 72
rect 27 62 33 68
rect 27 58 28 62
rect 32 58 33 62
rect 27 22 33 58
rect 39 82 45 87
rect 39 78 40 82
rect 44 78 45 82
rect 39 72 45 78
rect 39 68 40 72
rect 44 68 45 72
rect 39 62 45 68
rect 39 58 40 62
rect 44 58 45 62
rect 39 57 45 58
rect 27 18 28 22
rect 32 18 33 22
rect 3 17 9 18
rect 27 17 33 18
rect 39 22 45 23
rect 39 18 40 22
rect 44 18 45 22
rect 39 13 45 18
rect -2 12 52 13
rect -2 8 16 12
rect 20 8 40 12
rect 44 8 52 12
rect -2 -1 52 8
<< ntransistor >>
rect 11 15 13 25
rect 23 5 25 25
rect 35 5 37 25
<< ptransistor >>
rect 11 55 13 75
rect 23 55 25 95
rect 35 55 37 95
<< polycontact >>
rect 14 48 18 52
rect 4 38 8 42
rect 14 28 18 32
<< ndcontact >>
rect 4 18 8 22
rect 16 8 20 12
rect 28 18 32 22
rect 40 18 44 22
rect 40 8 44 12
<< pdcontact >>
rect 16 88 20 92
rect 4 68 8 72
rect 4 58 8 62
rect 28 78 32 82
rect 28 68 32 72
rect 28 58 32 62
rect 40 88 44 92
rect 40 78 44 82
rect 40 68 44 72
rect 40 58 44 62
<< nsubstratencontact >>
rect 4 92 8 96
rect 4 82 8 86
<< nsubstratendiff >>
rect 3 96 9 97
rect 3 92 4 96
rect 8 92 9 96
rect 3 86 9 92
rect 3 82 4 86
rect 8 82 9 86
rect 3 81 9 82
<< labels >>
rlabel metal1 20 50 20 50 6 i
rlabel metal1 20 50 20 50 6 i
rlabel metal1 25 6 25 6 6 vss
rlabel metal1 25 6 25 6 6 vss
rlabel metal1 30 50 30 50 6 q
rlabel metal1 30 50 30 50 6 q
rlabel metal1 25 94 25 94 6 vdd
rlabel metal1 25 94 25 94 6 vdd
<< end >>
