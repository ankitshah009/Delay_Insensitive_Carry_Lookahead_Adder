.subckt nd3v0x2 a b c vdd vss z
*   SPICE3 file   created from nd3v0x2.ext -      technology: scmos
m00 z      b      vdd    vdd p w=14u  l=2.3636u ad=65.3333p pd=20u      as=116.667p ps=33.3333u
m01 vdd    b      z      vdd p w=14u  l=2.3636u ad=116.667p pd=33.3333u as=65.3333p ps=20u
m02 z      c      vdd    vdd p w=28u  l=2.3636u ad=130.667p pd=40u      as=233.333p ps=66.6667u
m03 vdd    a      z      vdd p w=28u  l=2.3636u ad=233.333p pd=66.6667u as=130.667p ps=40u
m04 w1     a      vss    vss n w=14u  l=2.3636u ad=35p      pd=19u      as=126p     ps=46u
m05 w2     b      w1     vss n w=14u  l=2.3636u ad=35p      pd=19u      as=35p      ps=19u
m06 z      c      w2     vss n w=14u  l=2.3636u ad=56p      pd=22u      as=35p      ps=19u
m07 w3     c      z      vss n w=14u  l=2.3636u ad=35p      pd=19u      as=56p      ps=22u
m08 w4     b      w3     vss n w=14u  l=2.3636u ad=35p      pd=19u      as=35p      ps=19u
m09 vss    a      w4     vss n w=14u  l=2.3636u ad=126p     pd=46u      as=35p      ps=19u
C0  w4     a      0.007f
C1  w2     z      0.010f
C2  vss    z      0.240f
C3  w2     a      0.008f
C4  z      vdd    0.385f
C5  vss    a      0.106f
C6  z      c      0.102f
C7  vss    b      0.028f
C8  vdd    a      0.046f
C9  vdd    b      0.043f
C10 a      c      0.191f
C11 c      b      0.136f
C12 w3     a      0.007f
C13 w1     z      0.015f
C14 vss    vdd    0.005f
C15 vss    c      0.022f
C16 z      a      0.296f
C17 z      b      0.142f
C18 vdd    c      0.021f
C19 a      b      0.206f
C21 z      vss    0.013f
C23 a      vss    0.033f
C24 c      vss    0.022f
C25 b      vss    0.047f
.ends
