magic
tech scmos
timestamp 1179386978
<< checkpaint >>
rect -22 -25 94 105
<< ab >>
rect 0 0 72 80
<< pwell >>
rect -4 -7 76 36
<< nwell >>
rect -4 36 76 87
<< polysilicon >>
rect 9 64 11 69
rect 21 60 23 65
rect 9 37 11 52
rect 44 58 46 63
rect 54 58 56 63
rect 61 58 63 63
rect 21 47 23 50
rect 15 46 23 47
rect 44 46 46 50
rect 15 42 16 46
rect 20 44 23 46
rect 40 44 46 46
rect 20 42 21 44
rect 15 41 21 42
rect 9 36 15 37
rect 9 32 10 36
rect 14 32 15 36
rect 9 31 15 32
rect 9 28 11 31
rect 19 29 21 41
rect 40 39 42 44
rect 54 39 56 42
rect 25 38 42 39
rect 25 34 26 38
rect 30 37 42 38
rect 30 34 31 37
rect 25 33 31 34
rect 40 30 42 37
rect 49 38 56 39
rect 49 34 50 38
rect 54 34 56 38
rect 49 33 56 34
rect 61 39 63 42
rect 61 38 67 39
rect 61 34 62 38
rect 66 34 67 38
rect 61 33 67 34
rect 50 30 52 33
rect 19 26 22 29
rect 20 23 22 26
rect 61 23 63 33
rect 9 17 11 22
rect 40 18 42 23
rect 50 18 52 23
rect 20 12 22 17
rect 61 11 63 16
<< ndiffusion >>
rect 33 29 40 30
rect 2 27 9 28
rect 2 23 3 27
rect 7 23 9 27
rect 2 22 9 23
rect 11 23 17 28
rect 33 25 34 29
rect 38 25 40 29
rect 33 23 40 25
rect 42 29 50 30
rect 42 25 44 29
rect 48 25 50 29
rect 42 23 50 25
rect 52 23 59 30
rect 11 22 20 23
rect 13 18 14 22
rect 18 18 20 22
rect 13 17 20 18
rect 22 22 29 23
rect 22 18 24 22
rect 28 18 29 22
rect 54 21 61 23
rect 22 17 29 18
rect 54 17 55 21
rect 59 17 61 21
rect 54 16 61 17
rect 63 22 70 23
rect 63 18 65 22
rect 69 18 70 22
rect 63 16 70 18
<< pdiffusion >>
rect 13 72 19 73
rect 13 68 14 72
rect 18 68 19 72
rect 13 64 19 68
rect 35 72 42 73
rect 35 68 37 72
rect 41 68 42 72
rect 2 63 9 64
rect 2 59 3 63
rect 7 59 9 63
rect 2 58 9 59
rect 4 52 9 58
rect 11 60 19 64
rect 11 52 21 60
rect 13 50 21 52
rect 23 56 28 60
rect 35 58 42 68
rect 23 55 31 56
rect 23 51 26 55
rect 30 51 31 55
rect 23 50 31 51
rect 35 50 44 58
rect 46 55 54 58
rect 46 51 48 55
rect 52 51 54 55
rect 46 50 54 51
rect 49 42 54 50
rect 56 42 61 58
rect 63 57 70 58
rect 63 53 65 57
rect 69 53 70 57
rect 63 42 70 53
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect -2 72 74 78
rect -2 68 14 72
rect 18 68 37 72
rect 41 68 74 72
rect 2 59 3 63
rect 7 59 62 63
rect 2 28 6 59
rect 26 55 30 56
rect 10 46 14 55
rect 10 42 16 46
rect 20 42 23 46
rect 26 38 30 51
rect 10 36 23 38
rect 14 34 23 36
rect 2 27 7 28
rect 2 23 3 27
rect 10 25 14 32
rect 26 30 30 34
rect 24 26 30 30
rect 34 51 48 55
rect 52 51 54 55
rect 34 49 54 51
rect 34 29 38 49
rect 58 46 62 59
rect 65 57 69 68
rect 65 52 69 53
rect 50 42 62 46
rect 50 38 54 42
rect 66 39 70 47
rect 50 33 54 34
rect 58 38 70 39
rect 58 34 62 38
rect 66 34 70 38
rect 58 33 70 34
rect 2 22 7 23
rect 24 22 28 26
rect 13 18 14 22
rect 18 18 19 22
rect 13 12 19 18
rect 24 17 28 18
rect 43 25 44 29
rect 48 25 69 29
rect 34 17 38 25
rect 65 22 69 25
rect 54 17 55 21
rect 59 17 60 21
rect 65 17 69 18
rect 54 12 60 17
rect -2 2 74 12
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
<< ntransistor >>
rect 9 22 11 28
rect 40 23 42 30
rect 50 23 52 30
rect 20 17 22 23
rect 61 16 63 23
<< ptransistor >>
rect 9 52 11 64
rect 21 50 23 60
rect 44 50 46 58
rect 54 42 56 58
rect 61 42 63 58
<< polycontact >>
rect 16 42 20 46
rect 10 32 14 36
rect 26 34 30 38
rect 50 34 54 38
rect 62 34 66 38
<< ndcontact >>
rect 3 23 7 27
rect 34 25 38 29
rect 44 25 48 29
rect 14 18 18 22
rect 24 18 28 22
rect 55 17 59 21
rect 65 18 69 22
<< pdcontact >>
rect 14 68 18 72
rect 37 68 41 72
rect 3 59 7 63
rect 26 51 30 55
rect 48 51 52 55
rect 65 53 69 57
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
<< psubstratepdiff >>
rect 0 2 72 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 72 2
rect 0 -3 72 -2
<< nsubstratendiff >>
rect 0 82 72 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 72 82
rect 0 77 72 78
<< labels >>
rlabel polycontact 28 36 28 36 6 bn
rlabel polycontact 52 36 52 36 6 a2n
rlabel metal1 4 42 4 42 6 a2n
rlabel metal1 12 28 12 28 6 a2
rlabel metal1 20 44 20 44 6 b
rlabel metal1 20 36 20 36 6 a2
rlabel metal1 12 52 12 52 6 b
rlabel metal1 36 6 36 6 6 vss
rlabel metal1 26 23 26 23 6 bn
rlabel metal1 36 36 36 36 6 z
rlabel metal1 28 41 28 41 6 bn
rlabel metal1 36 74 36 74 6 vdd
rlabel metal1 52 39 52 39 6 a2n
rlabel metal1 52 52 52 52 6 z
rlabel metal1 44 52 44 52 6 z
rlabel metal1 56 27 56 27 6 n1
rlabel metal1 67 23 67 23 6 n1
rlabel metal1 60 36 60 36 6 a1
rlabel metal1 68 40 68 40 6 a1
rlabel metal1 32 61 32 61 6 a2n
<< end >>
