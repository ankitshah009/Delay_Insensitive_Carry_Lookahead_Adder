magic
tech scmos
timestamp 1179387801
<< checkpaint >>
rect -22 -22 142 94
<< ab >>
rect 0 0 120 72
<< pwell >>
rect -4 -4 124 32
<< nwell >>
rect -4 32 124 76
<< polysilicon >>
rect 17 63 19 68
rect 29 63 31 68
rect 39 63 41 68
rect 49 63 51 68
rect 77 66 79 70
rect 2 50 8 51
rect 2 46 3 50
rect 7 46 8 50
rect 2 45 8 46
rect 6 41 8 45
rect 89 61 91 66
rect 99 61 101 66
rect 109 61 111 66
rect 77 47 79 50
rect 65 46 79 47
rect 17 41 19 44
rect 6 39 19 41
rect 9 21 11 39
rect 29 34 31 44
rect 39 35 41 44
rect 49 41 51 44
rect 65 42 66 46
rect 70 45 79 46
rect 70 42 71 45
rect 65 41 71 42
rect 45 40 51 41
rect 45 36 46 40
rect 50 36 51 40
rect 89 37 91 45
rect 45 35 51 36
rect 55 36 91 37
rect 99 36 101 45
rect 17 33 31 34
rect 17 29 18 33
rect 22 32 31 33
rect 35 34 41 35
rect 22 29 23 32
rect 35 30 36 34
rect 40 30 41 34
rect 35 29 41 30
rect 17 28 23 29
rect 20 21 22 28
rect 39 27 41 29
rect 30 21 32 25
rect 39 24 42 27
rect 40 21 42 24
rect 47 21 49 35
rect 55 32 56 36
rect 60 35 91 36
rect 95 35 101 36
rect 109 35 111 45
rect 60 32 61 35
rect 55 31 61 32
rect 65 30 71 31
rect 65 26 66 30
rect 70 26 71 30
rect 65 25 71 26
rect 69 22 71 25
rect 81 19 83 35
rect 95 31 96 35
rect 100 31 101 35
rect 95 30 101 31
rect 99 25 101 30
rect 105 34 111 35
rect 105 30 106 34
rect 110 30 111 34
rect 105 29 111 30
rect 91 19 93 24
rect 99 22 103 25
rect 101 19 103 22
rect 108 19 110 29
rect 9 4 11 12
rect 20 8 22 12
rect 30 4 32 12
rect 40 7 42 12
rect 47 7 49 12
rect 9 2 32 4
rect 69 4 71 15
rect 81 8 83 12
rect 91 4 93 12
rect 101 7 103 12
rect 108 7 110 12
rect 69 2 93 4
<< ndiffusion >>
rect 62 21 69 22
rect 2 20 9 21
rect 2 16 3 20
rect 7 16 9 20
rect 2 15 9 16
rect 4 12 9 15
rect 11 17 20 21
rect 11 13 14 17
rect 18 13 20 17
rect 11 12 20 13
rect 22 17 30 21
rect 22 13 24 17
rect 28 13 30 17
rect 22 12 30 13
rect 32 18 40 21
rect 32 14 34 18
rect 38 14 40 18
rect 32 12 40 14
rect 42 12 47 21
rect 49 12 57 21
rect 62 17 63 21
rect 67 17 69 21
rect 62 15 69 17
rect 71 19 79 22
rect 71 15 81 19
rect 51 11 57 12
rect 51 7 52 11
rect 56 7 57 11
rect 51 6 57 7
rect 73 13 81 15
rect 73 9 74 13
rect 78 12 81 13
rect 83 18 91 19
rect 83 14 85 18
rect 89 14 91 18
rect 83 12 91 14
rect 93 18 101 19
rect 93 14 95 18
rect 99 14 101 18
rect 93 12 101 14
rect 103 12 108 19
rect 110 12 118 19
rect 78 9 79 12
rect 73 8 79 9
rect 112 8 118 12
rect 112 4 113 8
rect 117 4 118 8
rect 112 3 118 4
<< pdiffusion >>
rect 21 68 27 69
rect 21 64 22 68
rect 26 64 27 68
rect 21 63 27 64
rect 81 68 87 69
rect 81 66 82 68
rect 12 50 17 63
rect 10 49 17 50
rect 10 45 11 49
rect 15 45 17 49
rect 10 44 17 45
rect 19 44 29 63
rect 31 49 39 63
rect 31 45 33 49
rect 37 45 39 49
rect 31 44 39 45
rect 41 50 49 63
rect 41 46 43 50
rect 47 46 49 50
rect 41 44 49 46
rect 51 59 56 63
rect 72 60 77 66
rect 70 59 77 60
rect 51 58 58 59
rect 51 54 53 58
rect 57 54 58 58
rect 70 55 71 59
rect 75 55 77 59
rect 70 54 77 55
rect 51 53 58 54
rect 51 44 56 53
rect 72 50 77 54
rect 79 64 82 66
rect 86 64 87 68
rect 79 61 87 64
rect 79 50 89 61
rect 81 45 89 50
rect 91 50 99 61
rect 91 46 93 50
rect 97 46 99 50
rect 91 45 99 46
rect 101 51 109 61
rect 101 47 103 51
rect 107 47 109 51
rect 101 45 109 47
rect 111 59 118 61
rect 111 55 113 59
rect 117 55 118 59
rect 111 54 118 55
rect 111 45 116 54
<< metal1 >>
rect -2 68 122 72
rect -2 64 22 68
rect 26 64 61 68
rect 65 64 82 68
rect 86 64 122 68
rect 2 54 15 59
rect 26 54 53 58
rect 57 54 58 58
rect 70 55 71 59
rect 75 55 113 59
rect 117 55 118 59
rect 2 50 7 54
rect 26 50 30 54
rect 2 46 3 50
rect 2 45 7 46
rect 11 49 30 50
rect 15 46 30 49
rect 11 39 15 45
rect 3 35 15 39
rect 3 20 7 35
rect 18 33 22 35
rect 26 34 30 46
rect 33 49 37 50
rect 42 46 43 50
rect 47 46 58 50
rect 33 42 37 45
rect 33 40 50 42
rect 33 38 46 40
rect 26 30 36 34
rect 40 30 41 34
rect 18 27 22 29
rect 10 21 22 27
rect 46 26 50 36
rect 26 22 50 26
rect 54 36 58 46
rect 66 46 70 51
rect 66 38 79 42
rect 54 32 56 36
rect 60 32 61 36
rect 26 17 30 22
rect 54 18 58 32
rect 66 30 70 38
rect 84 35 88 55
rect 93 50 97 51
rect 102 47 103 51
rect 107 47 118 51
rect 93 43 97 46
rect 93 39 110 43
rect 66 25 70 26
rect 76 31 96 35
rect 100 31 101 35
rect 106 34 110 39
rect 76 21 80 31
rect 106 27 110 30
rect 3 15 7 16
rect 13 13 14 17
rect 18 13 19 17
rect 23 13 24 17
rect 28 13 30 17
rect 33 14 34 18
rect 38 14 58 18
rect 62 17 63 21
rect 67 17 80 21
rect 85 23 110 27
rect 85 18 89 23
rect 114 18 118 47
rect 94 14 95 18
rect 99 14 118 18
rect 85 13 89 14
rect 13 8 19 13
rect 51 8 52 11
rect -2 7 52 8
rect 56 8 57 11
rect 73 9 74 13
rect 78 9 79 13
rect 73 8 79 9
rect 56 7 62 8
rect -2 4 62 7
rect 66 4 113 8
rect 117 4 122 8
rect -2 0 122 4
<< ntransistor >>
rect 9 12 11 21
rect 20 12 22 21
rect 30 12 32 21
rect 40 12 42 21
rect 47 12 49 21
rect 69 15 71 22
rect 81 12 83 19
rect 91 12 93 19
rect 101 12 103 19
rect 108 12 110 19
<< ptransistor >>
rect 17 44 19 63
rect 29 44 31 63
rect 39 44 41 63
rect 49 44 51 63
rect 77 50 79 66
rect 89 45 91 61
rect 99 45 101 61
rect 109 45 111 61
<< polycontact >>
rect 3 46 7 50
rect 66 42 70 46
rect 46 36 50 40
rect 18 29 22 33
rect 36 30 40 34
rect 56 32 60 36
rect 66 26 70 30
rect 96 31 100 35
rect 106 30 110 34
<< ndcontact >>
rect 3 16 7 20
rect 14 13 18 17
rect 24 13 28 17
rect 34 14 38 18
rect 63 17 67 21
rect 52 7 56 11
rect 74 9 78 13
rect 85 14 89 18
rect 95 14 99 18
rect 113 4 117 8
<< pdcontact >>
rect 22 64 26 68
rect 11 45 15 49
rect 33 45 37 49
rect 43 46 47 50
rect 53 54 57 58
rect 71 55 75 59
rect 82 64 86 68
rect 93 46 97 50
rect 103 47 107 51
rect 113 55 117 59
<< psubstratepcontact >>
rect 62 4 66 8
<< nsubstratencontact >>
rect 61 64 65 68
<< psubstratepdiff >>
rect 61 8 67 9
rect 61 4 62 8
rect 66 4 67 8
rect 61 3 67 4
<< nsubstratendiff >>
rect 60 68 66 69
rect 60 64 61 68
rect 65 64 66 68
rect 60 63 66 64
<< labels >>
rlabel polycontact 38 32 38 32 6 bn
rlabel polycontact 48 38 48 38 6 an
rlabel polycontact 58 34 58 34 6 iz
rlabel polysilicon 109 21 109 21 6 zn
rlabel polycontact 98 33 98 33 6 cn
rlabel metal1 12 24 12 24 6 a
rlabel metal1 5 27 5 27 6 bn
rlabel metal1 13 42 13 42 6 bn
rlabel metal1 4 52 4 52 6 b
rlabel metal1 12 56 12 56 6 b
rlabel ndcontact 26 15 26 15 6 an
rlabel metal1 33 32 33 32 6 bn
rlabel metal1 20 28 20 28 6 a
rlabel metal1 35 44 35 44 6 an
rlabel metal1 60 4 60 4 6 vss
rlabel metal1 45 16 45 16 6 iz
rlabel metal1 48 32 48 32 6 an
rlabel metal1 68 40 68 40 6 c
rlabel metal1 56 32 56 32 6 iz
rlabel metal1 50 48 50 48 6 iz
rlabel metal1 42 56 42 56 6 bn
rlabel metal1 60 68 60 68 6 vdd
rlabel metal1 87 20 87 20 6 zn
rlabel metal1 71 19 71 19 6 cn
rlabel metal1 76 40 76 40 6 c
rlabel metal1 108 16 108 16 6 z
rlabel metal1 100 16 100 16 6 z
rlabel metal1 88 33 88 33 6 cn
rlabel metal1 116 36 116 36 6 z
rlabel metal1 95 45 95 45 6 zn
rlabel polycontact 108 33 108 33 6 zn
rlabel metal1 94 57 94 57 6 cn
<< end >>
