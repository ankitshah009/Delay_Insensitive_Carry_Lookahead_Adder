magic
tech scmos
timestamp 1180640139
<< checkpaint >>
rect -24 -26 84 126
<< ab >>
rect 0 0 60 100
<< pwell >>
rect -4 -6 64 49
<< nwell >>
rect -4 49 64 106
<< polysilicon >>
rect 31 93 33 98
rect 39 93 41 98
rect 47 93 49 98
rect 15 76 17 81
rect 15 49 17 56
rect 31 49 33 56
rect 39 53 41 56
rect 15 48 23 49
rect 15 45 18 48
rect 11 44 18 45
rect 22 44 23 48
rect 11 43 23 44
rect 27 48 33 49
rect 27 44 28 48
rect 32 44 33 48
rect 27 43 33 44
rect 37 52 43 53
rect 37 48 38 52
rect 42 48 43 52
rect 37 47 43 48
rect 11 27 13 43
rect 27 29 29 43
rect 37 30 39 47
rect 23 27 29 29
rect 35 27 39 30
rect 47 33 49 56
rect 47 32 53 33
rect 47 28 48 32
rect 52 28 53 32
rect 47 27 53 28
rect 23 24 25 27
rect 35 24 37 27
rect 47 24 49 27
rect 11 12 13 17
rect 23 12 25 17
rect 35 12 37 17
rect 47 12 49 17
<< ndiffusion >>
rect 6 23 11 27
rect 3 22 11 23
rect 3 18 4 22
rect 8 18 11 22
rect 3 17 11 18
rect 13 24 21 27
rect 13 17 23 24
rect 25 23 35 24
rect 25 19 28 23
rect 32 19 35 23
rect 25 17 35 19
rect 37 17 47 24
rect 49 22 57 24
rect 49 18 52 22
rect 56 18 57 22
rect 49 17 57 18
rect 15 12 21 17
rect 39 12 45 17
rect 15 8 16 12
rect 20 8 21 12
rect 15 7 21 8
rect 39 8 40 12
rect 44 8 45 12
rect 39 7 45 8
<< pdiffusion >>
rect 19 92 31 93
rect 19 88 22 92
rect 26 88 31 92
rect 19 76 31 88
rect 10 70 15 76
rect 7 69 15 70
rect 7 65 8 69
rect 12 65 15 69
rect 7 61 15 65
rect 7 57 8 61
rect 12 57 15 61
rect 7 56 15 57
rect 17 56 31 76
rect 33 56 39 93
rect 41 56 47 93
rect 49 81 54 93
rect 49 80 57 81
rect 49 76 52 80
rect 56 76 57 80
rect 49 72 57 76
rect 49 68 52 72
rect 56 68 57 72
rect 49 67 57 68
rect 49 56 54 67
<< metal1 >>
rect -2 92 62 100
rect -2 88 22 92
rect 26 88 62 92
rect 18 80 56 82
rect 18 78 52 80
rect 8 69 12 73
rect 8 61 12 65
rect 8 22 12 57
rect 18 48 22 78
rect 27 68 42 73
rect 18 32 22 44
rect 28 48 32 63
rect 38 52 42 68
rect 52 72 56 76
rect 52 67 56 68
rect 38 47 42 48
rect 28 42 32 44
rect 28 37 43 42
rect 48 32 52 53
rect 18 28 32 32
rect 28 23 32 28
rect 37 28 48 32
rect 37 27 52 28
rect 3 18 4 22
rect 8 18 23 22
rect 32 19 52 22
rect 28 18 52 19
rect 56 18 57 22
rect -2 8 16 12
rect 20 8 40 12
rect 44 8 62 12
rect -2 0 62 8
<< ntransistor >>
rect 11 17 13 27
rect 23 17 25 24
rect 35 17 37 24
rect 47 17 49 24
<< ptransistor >>
rect 15 56 17 76
rect 31 56 33 93
rect 39 56 41 93
rect 47 56 49 93
<< polycontact >>
rect 18 44 22 48
rect 28 44 32 48
rect 38 48 42 52
rect 48 28 52 32
<< ndcontact >>
rect 4 18 8 22
rect 28 19 32 23
rect 52 18 56 22
rect 16 8 20 12
rect 40 8 44 12
<< pdcontact >>
rect 22 88 26 92
rect 8 65 12 69
rect 8 57 12 61
rect 52 76 56 80
rect 52 68 56 72
<< psubstratepcontact >>
rect 28 4 32 8
<< nsubstratencontact >>
rect 8 92 12 96
<< psubstratepdiff >>
rect 27 8 33 9
rect 27 4 28 8
rect 32 4 33 8
rect 27 3 33 4
<< nsubstratendiff >>
rect 7 96 13 97
rect 7 92 8 96
rect 12 92 13 96
rect 7 91 13 92
<< labels >>
rlabel polycontact 19 46 19 46 6 zn
rlabel metal1 10 45 10 45 6 z
rlabel metal1 10 45 10 45 6 z
rlabel metal1 20 20 20 20 6 z
rlabel metal1 20 20 20 20 6 z
rlabel metal1 20 55 20 55 6 zn
rlabel metal1 30 6 30 6 6 vss
rlabel metal1 30 6 30 6 6 vss
rlabel metal1 30 25 30 25 6 zn
rlabel metal1 40 40 40 40 6 a
rlabel metal1 40 30 40 30 6 c
rlabel metal1 40 40 40 40 6 a
rlabel metal1 40 30 40 30 6 c
rlabel metal1 30 50 30 50 6 a
rlabel metal1 30 50 30 50 6 a
rlabel metal1 30 70 30 70 6 b
rlabel metal1 30 70 30 70 6 b
rlabel metal1 40 60 40 60 6 b
rlabel metal1 40 60 40 60 6 b
rlabel metal1 30 94 30 94 6 vdd
rlabel metal1 30 94 30 94 6 vdd
rlabel metal1 42 20 42 20 6 zn
rlabel metal1 50 40 50 40 6 c
rlabel metal1 50 40 50 40 6 c
rlabel metal1 54 74 54 74 6 zn
<< end >>
