magic
tech scmos
timestamp 1179386749
<< checkpaint >>
rect -22 -22 86 94
<< ab >>
rect 0 0 64 72
<< pwell >>
rect -4 -4 68 32
<< nwell >>
rect -4 32 68 76
<< polysilicon >>
rect 9 66 11 70
rect 16 66 18 70
rect 26 66 28 70
rect 33 66 35 70
rect 43 66 45 70
rect 50 66 52 70
rect 9 29 11 38
rect 16 35 18 38
rect 26 35 28 38
rect 16 34 28 35
rect 16 33 23 34
rect 22 30 23 33
rect 27 30 28 34
rect 22 29 28 30
rect 33 35 35 38
rect 43 35 45 38
rect 50 35 52 38
rect 33 34 45 35
rect 33 30 34 34
rect 38 33 45 34
rect 49 34 55 35
rect 38 30 39 33
rect 33 29 39 30
rect 49 30 50 34
rect 54 30 55 34
rect 49 29 55 30
rect 9 28 15 29
rect 9 24 10 28
rect 14 24 15 28
rect 23 24 25 29
rect 35 24 37 29
rect 49 25 51 29
rect 9 23 15 24
rect 13 20 15 23
rect 45 23 51 25
rect 45 20 47 23
rect 35 8 37 13
rect 45 8 47 13
rect 13 2 15 7
rect 23 2 25 7
<< ndiffusion >>
rect 18 20 23 24
rect 4 8 13 20
rect 4 4 6 8
rect 10 7 13 8
rect 15 18 23 20
rect 15 14 17 18
rect 21 14 23 18
rect 15 7 23 14
rect 25 13 35 24
rect 37 20 42 24
rect 37 18 45 20
rect 37 14 39 18
rect 43 14 45 18
rect 37 13 45 14
rect 47 18 55 20
rect 47 14 49 18
rect 53 14 55 18
rect 47 13 55 14
rect 25 8 33 13
rect 25 7 28 8
rect 10 4 11 7
rect 4 3 11 4
rect 27 4 28 7
rect 32 4 33 8
rect 27 3 33 4
<< pdiffusion >>
rect 4 51 9 66
rect 2 50 9 51
rect 2 46 3 50
rect 7 46 9 50
rect 2 43 9 46
rect 2 39 3 43
rect 7 39 9 43
rect 2 38 9 39
rect 11 38 16 66
rect 18 65 26 66
rect 18 61 20 65
rect 24 61 26 65
rect 18 58 26 61
rect 18 54 20 58
rect 24 54 26 58
rect 18 38 26 54
rect 28 38 33 66
rect 35 58 43 66
rect 35 54 37 58
rect 41 54 43 58
rect 35 51 43 54
rect 35 47 37 51
rect 41 47 43 51
rect 35 38 43 47
rect 45 38 50 66
rect 52 65 60 66
rect 52 61 54 65
rect 58 61 60 65
rect 52 58 60 61
rect 52 54 54 58
rect 58 54 60 58
rect 52 38 60 54
<< metal1 >>
rect -2 65 66 72
rect -2 64 20 65
rect 19 61 20 64
rect 24 64 54 65
rect 24 61 25 64
rect 19 58 25 61
rect 53 61 54 64
rect 58 64 66 65
rect 58 61 59 64
rect 19 54 20 58
rect 24 54 25 58
rect 37 58 41 59
rect 53 58 59 61
rect 53 54 54 58
rect 58 54 59 58
rect 37 51 41 54
rect 2 46 3 50
rect 7 47 37 50
rect 7 46 41 47
rect 2 43 7 46
rect 2 39 3 43
rect 2 38 7 39
rect 22 38 55 42
rect 2 18 6 38
rect 22 34 28 38
rect 49 34 55 38
rect 22 30 23 34
rect 27 30 28 34
rect 33 30 34 34
rect 38 30 39 34
rect 49 30 50 34
rect 54 30 55 34
rect 10 28 14 29
rect 33 26 39 30
rect 14 24 39 26
rect 10 22 39 24
rect 49 18 53 19
rect 2 14 17 18
rect 21 14 39 18
rect 43 14 44 18
rect 49 8 53 14
rect -2 4 6 8
rect 10 4 28 8
rect 32 4 56 8
rect 60 4 66 8
rect -2 0 66 4
<< ntransistor >>
rect 13 7 15 20
rect 23 7 25 24
rect 35 13 37 24
rect 45 13 47 20
<< ptransistor >>
rect 9 38 11 66
rect 16 38 18 66
rect 26 38 28 66
rect 33 38 35 66
rect 43 38 45 66
rect 50 38 52 66
<< polycontact >>
rect 23 30 27 34
rect 34 30 38 34
rect 50 30 54 34
rect 10 24 14 28
<< ndcontact >>
rect 6 4 10 8
rect 17 14 21 18
rect 39 14 43 18
rect 49 14 53 18
rect 28 4 32 8
<< pdcontact >>
rect 3 46 7 50
rect 3 39 7 43
rect 20 61 24 65
rect 20 54 24 58
rect 37 54 41 58
rect 37 47 41 51
rect 54 61 58 65
rect 54 54 58 58
<< psubstratepcontact >>
rect 56 4 60 8
<< psubstratepdiff >>
rect 55 8 61 9
rect 55 4 56 8
rect 60 4 61 8
rect 55 3 61 4
<< labels >>
rlabel metal1 12 16 12 16 6 z
rlabel metal1 4 32 4 32 6 z
rlabel metal1 12 48 12 48 6 z
rlabel ndcontact 20 16 20 16 6 z
rlabel metal1 28 16 28 16 6 z
rlabel metal1 20 24 20 24 6 b
rlabel metal1 28 24 28 24 6 b
rlabel metal1 28 40 28 40 6 a
rlabel metal1 20 48 20 48 6 z
rlabel metal1 28 48 28 48 6 z
rlabel metal1 32 4 32 4 6 vss
rlabel metal1 36 16 36 16 6 z
rlabel metal1 36 28 36 28 6 b
rlabel metal1 44 40 44 40 6 a
rlabel metal1 36 40 36 40 6 a
rlabel metal1 36 48 36 48 6 z
rlabel metal1 32 68 32 68 6 vdd
rlabel metal1 52 36 52 36 6 a
<< end >>
