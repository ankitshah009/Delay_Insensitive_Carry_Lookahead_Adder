magic
tech scmos
timestamp 1179385165
<< checkpaint >>
rect -22 -25 86 105
<< ab >>
rect 0 0 64 80
<< pwell >>
rect -4 -7 68 36
<< nwell >>
rect -4 36 68 87
<< polysilicon >>
rect 9 61 11 65
rect 20 64 22 69
rect 30 64 32 69
rect 42 64 44 69
rect 52 64 54 69
rect 9 39 11 43
rect 20 39 22 58
rect 30 47 32 58
rect 42 47 44 58
rect 29 46 35 47
rect 29 42 30 46
rect 34 42 35 46
rect 29 41 35 42
rect 42 46 48 47
rect 42 42 43 46
rect 47 42 48 46
rect 42 41 48 42
rect 9 38 15 39
rect 9 34 10 38
rect 14 34 15 38
rect 9 33 15 34
rect 19 38 25 39
rect 19 34 20 38
rect 24 34 25 38
rect 19 33 25 34
rect 9 25 11 33
rect 22 25 24 33
rect 29 25 31 41
rect 42 36 44 41
rect 36 34 44 36
rect 52 39 54 58
rect 52 38 58 39
rect 52 34 53 38
rect 57 34 58 38
rect 36 25 38 34
rect 52 33 58 34
rect 52 30 54 33
rect 43 28 54 30
rect 43 25 45 28
rect 9 11 11 16
rect 22 12 24 17
rect 29 12 31 17
rect 36 12 38 17
rect 43 12 45 17
<< ndiffusion >>
rect 4 22 9 25
rect 2 21 9 22
rect 2 17 3 21
rect 7 17 9 21
rect 2 16 9 17
rect 11 17 22 25
rect 24 17 29 25
rect 31 17 36 25
rect 38 17 43 25
rect 45 23 50 25
rect 45 22 52 23
rect 45 18 47 22
rect 51 18 52 22
rect 45 17 52 18
rect 11 16 20 17
rect 13 12 20 16
rect 13 8 14 12
rect 18 8 20 12
rect 13 7 20 8
<< pdiffusion >>
rect 34 72 40 73
rect 34 68 35 72
rect 39 68 40 72
rect 34 64 40 68
rect 13 63 20 64
rect 13 61 14 63
rect 4 56 9 61
rect 2 55 9 56
rect 2 51 3 55
rect 7 51 9 55
rect 2 48 9 51
rect 2 44 3 48
rect 7 44 9 48
rect 2 43 9 44
rect 11 59 14 61
rect 18 59 20 63
rect 11 58 20 59
rect 22 63 30 64
rect 22 59 24 63
rect 28 59 30 63
rect 22 58 30 59
rect 32 58 42 64
rect 44 63 52 64
rect 44 59 46 63
rect 50 59 52 63
rect 44 58 52 59
rect 54 63 61 64
rect 54 59 56 63
rect 60 59 61 63
rect 54 58 61 59
rect 11 43 18 58
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect -2 72 66 78
rect -2 68 35 72
rect 39 68 66 72
rect 14 63 18 68
rect 55 63 61 68
rect 2 55 7 63
rect 14 58 18 59
rect 23 59 24 63
rect 28 59 46 63
rect 50 59 51 63
rect 55 59 56 63
rect 60 59 61 63
rect 2 51 3 55
rect 23 54 27 59
rect 2 48 7 51
rect 2 44 3 48
rect 2 43 7 44
rect 11 50 27 54
rect 33 50 47 54
rect 2 22 6 43
rect 11 39 15 50
rect 33 46 37 50
rect 58 46 62 55
rect 25 42 30 46
rect 34 42 37 46
rect 41 42 43 46
rect 47 42 62 46
rect 10 38 15 39
rect 14 34 15 38
rect 19 34 20 38
rect 24 34 31 38
rect 41 34 53 38
rect 57 34 62 38
rect 10 33 15 34
rect 11 30 15 33
rect 27 30 31 34
rect 11 26 23 30
rect 27 26 47 30
rect 19 22 23 26
rect 2 21 15 22
rect 2 17 3 21
rect 7 17 15 21
rect 19 18 47 22
rect 51 18 52 22
rect 58 17 62 34
rect -2 8 14 12
rect 18 8 66 12
rect -2 2 66 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
<< ntransistor >>
rect 9 16 11 25
rect 22 17 24 25
rect 29 17 31 25
rect 36 17 38 25
rect 43 17 45 25
<< ptransistor >>
rect 9 43 11 61
rect 20 58 22 64
rect 30 58 32 64
rect 42 58 44 64
rect 52 58 54 64
<< polycontact >>
rect 30 42 34 46
rect 43 42 47 46
rect 10 34 14 38
rect 20 34 24 38
rect 53 34 57 38
<< ndcontact >>
rect 3 17 7 21
rect 47 18 51 22
rect 14 8 18 12
<< pdcontact >>
rect 35 68 39 72
rect 3 51 7 55
rect 3 44 7 48
rect 14 59 18 63
rect 24 59 28 63
rect 46 59 50 63
rect 56 59 60 63
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
<< psubstratepdiff >>
rect 0 2 64 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 64 2
rect 0 -3 64 -2
<< nsubstratendiff >>
rect 0 82 64 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 64 82
rect 0 77 64 78
<< labels >>
rlabel polycontact 12 36 12 36 6 zn
rlabel metal1 4 40 4 40 6 z
rlabel metal1 12 20 12 20 6 z
rlabel metal1 13 40 13 40 6 zn
rlabel metal1 32 6 32 6 6 vss
rlabel metal1 36 28 36 28 6 a
rlabel metal1 28 36 28 36 6 a
rlabel metal1 28 44 28 44 6 b
rlabel metal1 36 52 36 52 6 b
rlabel metal1 32 74 32 74 6 vdd
rlabel metal1 35 20 35 20 6 zn
rlabel metal1 44 28 44 28 6 a
rlabel metal1 44 36 44 36 6 d
rlabel polycontact 44 44 44 44 6 c
rlabel metal1 44 52 44 52 6 b
rlabel metal1 37 61 37 61 6 zn
rlabel metal1 60 24 60 24 6 d
rlabel metal1 52 36 52 36 6 d
rlabel metal1 52 44 52 44 6 c
rlabel metal1 60 52 60 52 6 c
<< end >>
