magic
tech scmos
timestamp 1179386652
<< checkpaint >>
rect -22 -22 102 94
<< ab >>
rect 0 0 80 72
<< pwell >>
rect -4 -4 84 32
<< nwell >>
rect -4 32 84 76
<< polysilicon >>
rect 9 65 11 70
rect 19 65 21 70
rect 32 65 34 70
rect 42 65 44 70
rect 64 50 70 51
rect 64 46 65 50
rect 69 46 70 50
rect 64 45 70 46
rect 54 42 60 43
rect 9 31 11 40
rect 19 37 21 40
rect 32 37 34 40
rect 19 36 25 37
rect 19 32 20 36
rect 24 32 25 36
rect 32 36 38 37
rect 32 33 33 36
rect 19 31 25 32
rect 29 32 33 33
rect 37 32 38 36
rect 29 31 38 32
rect 42 35 44 40
rect 54 38 55 42
rect 59 38 60 42
rect 54 37 60 38
rect 42 34 49 35
rect 9 30 15 31
rect 9 26 10 30
rect 14 27 15 30
rect 14 26 17 27
rect 9 25 17 26
rect 15 22 17 25
rect 22 22 24 31
rect 29 22 31 31
rect 42 30 44 34
rect 48 30 49 34
rect 42 29 49 30
rect 42 27 48 29
rect 54 28 56 37
rect 64 33 66 45
rect 36 25 48 27
rect 36 22 38 25
rect 46 22 48 25
rect 53 25 56 28
rect 60 31 66 33
rect 53 22 55 25
rect 60 22 62 31
rect 72 30 78 31
rect 72 27 73 30
rect 67 26 73 27
rect 77 26 78 30
rect 67 25 78 26
rect 67 22 69 25
rect 15 2 17 7
rect 22 2 24 7
rect 29 2 31 7
rect 36 2 38 7
rect 46 2 48 7
rect 53 2 55 7
rect 60 2 62 7
rect 67 2 69 7
<< ndiffusion >>
rect 6 8 15 22
rect 6 4 8 8
rect 12 7 15 8
rect 17 7 22 22
rect 24 7 29 22
rect 31 7 36 22
rect 38 18 46 22
rect 38 14 40 18
rect 44 14 46 18
rect 38 7 46 14
rect 48 7 53 22
rect 55 7 60 22
rect 62 7 67 22
rect 69 12 77 22
rect 69 8 71 12
rect 75 8 77 12
rect 69 7 77 8
rect 12 4 13 7
rect 6 3 13 4
<< pdiffusion >>
rect 24 65 30 67
rect 2 64 9 65
rect 2 60 3 64
rect 7 60 9 64
rect 2 57 9 60
rect 2 53 3 57
rect 7 53 9 57
rect 2 40 9 53
rect 11 58 19 65
rect 11 54 13 58
rect 17 54 19 58
rect 11 50 19 54
rect 11 46 13 50
rect 17 46 19 50
rect 11 40 19 46
rect 21 61 25 65
rect 29 61 32 65
rect 21 40 32 61
rect 34 58 42 65
rect 34 54 36 58
rect 40 54 42 58
rect 34 40 42 54
rect 44 64 52 65
rect 44 60 46 64
rect 50 60 52 64
rect 44 57 52 60
rect 44 53 46 57
rect 50 53 52 57
rect 44 40 52 53
<< metal1 >>
rect -2 68 82 72
rect -2 65 57 68
rect -2 64 25 65
rect 2 60 3 64
rect 7 60 8 64
rect 24 61 25 64
rect 29 64 57 65
rect 61 64 72 68
rect 76 64 82 68
rect 29 61 30 64
rect 2 57 8 60
rect 45 60 46 64
rect 50 60 51 64
rect 2 53 3 57
rect 7 53 8 57
rect 12 54 13 58
rect 17 54 36 58
rect 40 54 41 58
rect 45 57 51 60
rect 12 50 18 54
rect 45 53 46 57
rect 50 53 51 57
rect 58 50 62 59
rect 2 46 13 50
rect 17 46 18 50
rect 24 46 65 50
rect 69 46 71 50
rect 2 18 6 46
rect 24 42 28 46
rect 17 38 28 42
rect 33 38 55 42
rect 59 38 60 42
rect 64 38 71 42
rect 20 36 24 38
rect 20 31 24 32
rect 33 36 39 38
rect 37 32 39 36
rect 64 34 68 38
rect 10 30 14 31
rect 33 30 39 32
rect 43 30 44 34
rect 48 30 68 34
rect 72 30 78 31
rect 72 26 73 30
rect 77 26 78 30
rect 10 22 78 26
rect 58 21 78 22
rect 2 14 40 18
rect 44 14 47 18
rect 58 13 62 21
rect 71 12 75 13
rect -2 4 8 8
rect 12 4 82 8
rect -2 0 82 4
<< ntransistor >>
rect 15 7 17 22
rect 22 7 24 22
rect 29 7 31 22
rect 36 7 38 22
rect 46 7 48 22
rect 53 7 55 22
rect 60 7 62 22
rect 67 7 69 22
<< ptransistor >>
rect 9 40 11 65
rect 19 40 21 65
rect 32 40 34 65
rect 42 40 44 65
<< polycontact >>
rect 65 46 69 50
rect 20 32 24 36
rect 33 32 37 36
rect 55 38 59 42
rect 10 26 14 30
rect 44 30 48 34
rect 73 26 77 30
<< ndcontact >>
rect 8 4 12 8
rect 40 14 44 18
rect 71 8 75 12
<< pdcontact >>
rect 3 60 7 64
rect 3 53 7 57
rect 13 54 17 58
rect 13 46 17 50
rect 25 61 29 65
rect 36 54 40 58
rect 46 60 50 64
rect 46 53 50 57
<< nsubstratencontact >>
rect 57 64 61 68
rect 72 64 76 68
<< nsubstratendiff >>
rect 56 68 77 69
rect 56 64 57 68
rect 61 64 72 68
rect 76 64 77 68
rect 56 63 77 64
<< labels >>
rlabel metal1 4 32 4 32 6 z
rlabel metal1 20 16 20 16 6 z
rlabel metal1 28 16 28 16 6 z
rlabel metal1 12 16 12 16 6 z
rlabel metal1 20 24 20 24 6 a
rlabel metal1 28 24 28 24 6 a
rlabel metal1 20 40 20 40 6 b
rlabel metal1 12 48 12 48 6 z
rlabel metal1 28 48 28 48 6 b
rlabel metal1 20 56 20 56 6 z
rlabel metal1 28 56 28 56 6 z
rlabel metal1 40 4 40 4 6 vss
rlabel metal1 36 16 36 16 6 z
rlabel metal1 44 16 44 16 6 z
rlabel metal1 36 24 36 24 6 a
rlabel metal1 44 24 44 24 6 a
rlabel metal1 44 40 44 40 6 c
rlabel metal1 36 36 36 36 6 c
rlabel metal1 36 48 36 48 6 b
rlabel metal1 44 48 44 48 6 b
rlabel metal1 36 56 36 56 6 z
rlabel metal1 40 68 40 68 6 vdd
rlabel metal1 52 24 52 24 6 a
rlabel metal1 60 20 60 20 6 a
rlabel metal1 60 32 60 32 6 d
rlabel metal1 52 32 52 32 6 d
rlabel metal1 52 40 52 40 6 c
rlabel metal1 52 48 52 48 6 b
rlabel metal1 60 52 60 52 6 b
rlabel metal1 68 24 68 24 6 a
rlabel metal1 76 24 76 24 6 a
rlabel metal1 68 40 68 40 6 d
rlabel polycontact 68 48 68 48 6 b
<< end >>
