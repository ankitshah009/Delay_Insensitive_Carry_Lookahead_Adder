magic
tech scmos
timestamp 1179386761
<< checkpaint >>
rect -22 -25 102 105
<< ab >>
rect 0 0 80 80
<< pwell >>
rect -4 -7 84 36
<< nwell >>
rect -4 36 84 87
<< polysilicon >>
rect 9 70 11 74
rect 16 70 18 74
rect 26 70 28 74
rect 33 70 35 74
rect 43 70 45 74
rect 50 70 52 74
rect 60 70 62 74
rect 67 70 69 74
rect 9 33 11 42
rect 16 39 18 42
rect 26 39 28 42
rect 16 38 28 39
rect 16 37 23 38
rect 22 34 23 37
rect 27 34 28 38
rect 33 39 35 42
rect 43 39 45 42
rect 33 37 45 39
rect 50 39 52 42
rect 60 39 62 42
rect 50 38 62 39
rect 22 33 28 34
rect 35 36 41 37
rect 9 32 18 33
rect 9 31 13 32
rect 12 28 13 31
rect 17 28 18 32
rect 12 27 18 28
rect 13 24 15 27
rect 23 24 25 33
rect 35 32 36 36
rect 40 32 41 36
rect 50 34 51 38
rect 55 37 62 38
rect 55 34 56 37
rect 50 33 56 34
rect 35 31 41 32
rect 45 31 56 33
rect 67 31 69 42
rect 35 28 37 31
rect 45 28 47 31
rect 63 30 69 31
rect 13 6 15 11
rect 23 6 25 11
rect 63 26 64 30
rect 68 26 69 30
rect 63 25 69 26
rect 35 6 37 11
rect 45 6 47 11
<< ndiffusion >>
rect 27 24 35 28
rect 4 12 13 24
rect 4 8 6 12
rect 10 11 13 12
rect 15 22 23 24
rect 15 18 17 22
rect 21 18 23 22
rect 15 11 23 18
rect 25 12 35 24
rect 25 11 28 12
rect 10 8 11 11
rect 4 7 11 8
rect 27 8 28 11
rect 32 11 35 12
rect 37 22 45 28
rect 37 18 39 22
rect 43 18 45 22
rect 37 11 45 18
rect 47 23 55 28
rect 47 19 49 23
rect 53 19 55 23
rect 47 16 55 19
rect 47 12 49 16
rect 53 12 55 16
rect 47 11 55 12
rect 32 8 33 11
rect 27 7 33 8
<< pdiffusion >>
rect 2 69 9 70
rect 2 65 3 69
rect 7 65 9 69
rect 2 62 9 65
rect 2 58 3 62
rect 7 58 9 62
rect 2 42 9 58
rect 11 42 16 70
rect 18 54 26 70
rect 18 50 20 54
rect 24 50 26 54
rect 18 47 26 50
rect 18 43 20 47
rect 24 43 26 47
rect 18 42 26 43
rect 28 42 33 70
rect 35 69 43 70
rect 35 65 37 69
rect 41 65 43 69
rect 35 62 43 65
rect 35 58 37 62
rect 41 58 43 62
rect 35 42 43 58
rect 45 42 50 70
rect 52 54 60 70
rect 52 50 54 54
rect 58 50 60 54
rect 52 47 60 50
rect 52 43 54 47
rect 58 43 60 47
rect 52 42 60 43
rect 62 42 67 70
rect 69 69 77 70
rect 69 65 71 69
rect 75 65 77 69
rect 69 62 77 65
rect 69 58 71 62
rect 75 58 77 62
rect 69 42 77 58
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect -2 69 82 78
rect -2 68 3 69
rect 2 65 3 68
rect 7 68 37 69
rect 7 65 8 68
rect 2 62 8 65
rect 2 58 3 62
rect 7 58 8 62
rect 36 65 37 68
rect 41 68 71 69
rect 41 65 42 68
rect 36 62 42 65
rect 36 58 37 62
rect 41 58 42 62
rect 70 65 71 68
rect 75 68 82 69
rect 75 65 76 68
rect 70 62 76 65
rect 70 58 71 62
rect 75 58 76 62
rect 19 50 20 54
rect 24 50 54 54
rect 58 50 59 54
rect 19 47 24 50
rect 2 43 20 47
rect 54 47 59 50
rect 2 42 24 43
rect 28 42 50 46
rect 58 46 59 47
rect 58 43 63 46
rect 54 42 63 43
rect 2 22 6 42
rect 28 38 32 42
rect 22 34 23 38
rect 27 34 32 38
rect 46 38 50 42
rect 36 36 40 37
rect 13 32 17 33
rect 46 34 51 38
rect 55 34 63 38
rect 36 30 40 32
rect 17 28 64 30
rect 13 26 64 28
rect 68 26 70 30
rect 2 18 17 22
rect 21 18 39 22
rect 43 18 44 22
rect 48 19 49 23
rect 53 19 54 23
rect 48 16 54 19
rect 66 17 70 26
rect 48 12 49 16
rect 53 12 54 16
rect -2 8 6 12
rect 10 8 28 12
rect 32 8 82 12
rect -2 2 82 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
<< ntransistor >>
rect 13 11 15 24
rect 23 11 25 24
rect 35 11 37 28
rect 45 11 47 28
<< ptransistor >>
rect 9 42 11 70
rect 16 42 18 70
rect 26 42 28 70
rect 33 42 35 70
rect 43 42 45 70
rect 50 42 52 70
rect 60 42 62 70
rect 67 42 69 70
<< polycontact >>
rect 23 34 27 38
rect 13 28 17 32
rect 36 32 40 36
rect 51 34 55 38
rect 64 26 68 30
<< ndcontact >>
rect 6 8 10 12
rect 17 18 21 22
rect 28 8 32 12
rect 39 18 43 22
rect 49 19 53 23
rect 49 12 53 16
<< pdcontact >>
rect 3 65 7 69
rect 3 58 7 62
rect 20 50 24 54
rect 20 43 24 47
rect 37 65 41 69
rect 37 58 41 62
rect 54 50 58 54
rect 54 43 58 47
rect 71 65 75 69
rect 71 58 75 62
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
<< psubstratepdiff >>
rect 0 2 80 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 80 2
rect 0 -3 80 -2
<< nsubstratendiff >>
rect 0 82 80 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 80 82
rect 0 77 80 78
<< labels >>
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 20 12 20 6 z
rlabel ndcontact 20 20 20 20 6 z
rlabel metal1 20 28 20 28 6 a
rlabel metal1 28 20 28 20 6 z
rlabel metal1 28 28 28 28 6 a
rlabel metal1 12 44 12 44 6 z
rlabel metal1 20 44 20 44 6 z
rlabel metal1 28 36 28 36 6 b
rlabel metal1 28 52 28 52 6 z
rlabel metal1 40 6 40 6 6 vss
rlabel metal1 36 20 36 20 6 z
rlabel metal1 36 28 36 28 6 a
rlabel metal1 44 28 44 28 6 a
rlabel metal1 36 44 36 44 6 b
rlabel metal1 44 44 44 44 6 b
rlabel metal1 36 52 36 52 6 z
rlabel metal1 44 52 44 52 6 z
rlabel metal1 40 74 40 74 6 vdd
rlabel metal1 52 28 52 28 6 a
rlabel metal1 60 28 60 28 6 a
rlabel polycontact 52 36 52 36 6 b
rlabel metal1 60 36 60 36 6 b
rlabel metal1 60 44 60 44 6 z
rlabel metal1 52 52 52 52 6 z
rlabel metal1 68 20 68 20 6 a
<< end >>
