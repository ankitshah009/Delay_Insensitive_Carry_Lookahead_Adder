magic
tech scmos
timestamp 1179386258
<< checkpaint >>
rect -22 -22 86 94
<< ab >>
rect 0 0 64 72
<< pwell >>
rect -4 -4 68 32
<< nwell >>
rect -4 32 68 76
<< polysilicon >>
rect 9 66 11 70
rect 19 66 21 70
rect 29 66 31 70
rect 39 66 41 70
rect 49 66 51 70
rect 9 35 11 42
rect 19 35 21 42
rect 29 35 31 42
rect 39 35 41 42
rect 49 36 51 39
rect 9 34 15 35
rect 9 30 10 34
rect 14 30 15 34
rect 9 29 15 30
rect 19 34 31 35
rect 19 30 26 34
rect 30 30 31 34
rect 19 29 31 30
rect 35 34 41 35
rect 35 30 36 34
rect 40 30 41 34
rect 45 35 51 36
rect 45 31 46 35
rect 50 31 51 35
rect 45 30 51 31
rect 35 29 41 30
rect 12 26 14 29
rect 19 26 21 29
rect 29 26 31 29
rect 36 26 38 29
rect 47 26 49 30
rect 47 7 49 12
rect 12 2 14 6
rect 19 2 21 6
rect 29 2 31 6
rect 36 2 38 6
<< ndiffusion >>
rect 4 11 12 26
rect 4 7 6 11
rect 10 7 12 11
rect 4 6 12 7
rect 14 6 19 26
rect 21 18 29 26
rect 21 14 23 18
rect 27 14 29 18
rect 21 6 29 14
rect 31 6 36 26
rect 38 18 47 26
rect 38 14 40 18
rect 44 14 47 18
rect 38 12 47 14
rect 49 25 56 26
rect 49 21 51 25
rect 55 21 56 25
rect 49 18 56 21
rect 49 14 51 18
rect 55 14 56 18
rect 49 12 56 14
rect 38 11 45 12
rect 38 7 40 11
rect 44 7 45 11
rect 38 6 45 7
<< pdiffusion >>
rect 2 65 9 66
rect 2 61 3 65
rect 7 61 9 65
rect 2 58 9 61
rect 2 54 3 58
rect 7 54 9 58
rect 2 42 9 54
rect 11 57 19 66
rect 11 53 13 57
rect 17 53 19 57
rect 11 50 19 53
rect 11 46 13 50
rect 17 46 19 50
rect 11 42 19 46
rect 21 65 29 66
rect 21 61 23 65
rect 27 61 29 65
rect 21 58 29 61
rect 21 54 23 58
rect 27 54 29 58
rect 21 42 29 54
rect 31 57 39 66
rect 31 53 33 57
rect 37 53 39 57
rect 31 50 39 53
rect 31 46 33 50
rect 37 46 39 50
rect 31 42 39 46
rect 41 65 49 66
rect 41 61 43 65
rect 47 61 49 65
rect 41 58 49 61
rect 41 54 43 58
rect 47 54 49 58
rect 41 42 49 54
rect 43 39 49 42
rect 51 52 56 66
rect 51 51 58 52
rect 51 47 53 51
rect 57 47 58 51
rect 51 44 58 47
rect 51 40 53 44
rect 57 40 58 44
rect 51 39 58 40
<< metal1 >>
rect -2 65 66 72
rect -2 64 3 65
rect 2 61 3 64
rect 7 64 23 65
rect 7 61 8 64
rect 2 58 8 61
rect 22 61 23 64
rect 27 64 43 65
rect 27 61 28 64
rect 22 58 28 61
rect 42 61 43 64
rect 47 64 66 65
rect 47 61 48 64
rect 2 54 3 58
rect 7 54 8 58
rect 13 57 17 58
rect 22 54 23 58
rect 27 54 28 58
rect 33 57 38 59
rect 13 50 17 53
rect 37 53 38 57
rect 42 58 48 61
rect 42 54 43 58
rect 47 54 48 58
rect 33 50 38 53
rect 53 51 57 52
rect 2 46 13 50
rect 17 46 33 50
rect 37 46 38 50
rect 2 18 6 46
rect 42 42 46 51
rect 53 44 57 47
rect 10 34 14 35
rect 17 34 23 42
rect 33 38 50 42
rect 46 35 50 38
rect 17 30 26 34
rect 30 30 31 34
rect 35 30 36 34
rect 40 30 41 34
rect 46 30 50 31
rect 10 26 14 30
rect 35 26 41 30
rect 53 26 57 40
rect 10 25 57 26
rect 10 22 51 25
rect 55 22 57 25
rect 51 18 55 21
rect 2 14 23 18
rect 27 14 31 18
rect 39 14 40 18
rect 44 14 45 18
rect 39 11 45 14
rect 51 13 55 14
rect 5 8 6 11
rect -2 7 6 8
rect 10 8 11 11
rect 39 8 40 11
rect 10 7 40 8
rect 44 8 45 11
rect 44 7 66 8
rect -2 0 66 7
<< ntransistor >>
rect 12 6 14 26
rect 19 6 21 26
rect 29 6 31 26
rect 36 6 38 26
rect 47 12 49 26
<< ptransistor >>
rect 9 42 11 66
rect 19 42 21 66
rect 29 42 31 66
rect 39 42 41 66
rect 49 39 51 66
<< polycontact >>
rect 10 30 14 34
rect 26 30 30 34
rect 36 30 40 34
rect 46 31 50 35
<< ndcontact >>
rect 6 7 10 11
rect 23 14 27 18
rect 40 14 44 18
rect 51 21 55 25
rect 51 14 55 18
rect 40 7 44 11
<< pdcontact >>
rect 3 61 7 65
rect 3 54 7 58
rect 13 53 17 57
rect 13 46 17 50
rect 23 61 27 65
rect 23 54 27 58
rect 33 53 37 57
rect 33 46 37 50
rect 43 61 47 65
rect 43 54 47 58
rect 53 47 57 51
rect 53 40 57 44
<< labels >>
rlabel polycontact 12 32 12 32 6 an
rlabel polycontact 38 32 38 32 6 an
rlabel metal1 12 16 12 16 6 z
rlabel metal1 12 28 12 28 6 an
rlabel metal1 4 32 4 32 6 z
rlabel metal1 12 48 12 48 6 z
rlabel metal1 20 16 20 16 6 z
rlabel metal1 28 16 28 16 6 z
rlabel polycontact 28 32 28 32 6 b
rlabel metal1 20 36 20 36 6 b
rlabel metal1 20 48 20 48 6 z
rlabel metal1 28 48 28 48 6 z
rlabel metal1 32 4 32 4 6 vss
rlabel metal1 38 28 38 28 6 an
rlabel metal1 36 40 36 40 6 a
rlabel metal1 44 44 44 44 6 a
rlabel pdcontact 36 56 36 56 6 z
rlabel metal1 32 68 32 68 6 vdd
rlabel metal1 53 19 53 19 6 an
rlabel metal1 55 37 55 37 6 an
<< end >>
