magic
tech scmos
timestamp 1185094761
<< checkpaint >>
rect -22 -22 72 122
<< ab >>
rect 0 0 50 100
<< pwell >>
rect -4 -4 54 48
<< nwell >>
rect -4 48 54 104
<< polysilicon >>
rect 15 78 17 82
rect 23 78 25 82
rect 37 73 39 78
rect 15 43 17 56
rect 23 52 25 56
rect 37 52 39 56
rect 23 49 27 52
rect 13 42 21 43
rect 13 38 16 42
rect 20 38 21 42
rect 13 37 21 38
rect 25 42 27 49
rect 32 51 39 52
rect 32 47 33 51
rect 37 47 39 51
rect 32 46 39 47
rect 25 41 32 42
rect 25 37 27 41
rect 31 37 32 41
rect 13 23 15 37
rect 25 36 32 37
rect 25 23 27 36
rect 37 26 39 46
rect 13 12 15 17
rect 25 12 27 17
rect 37 12 39 17
<< ndiffusion >>
rect 30 23 37 26
rect 4 17 13 23
rect 15 22 25 23
rect 15 18 18 22
rect 22 18 25 22
rect 15 17 25 18
rect 27 22 37 23
rect 27 18 30 22
rect 34 18 37 22
rect 27 17 37 18
rect 39 25 47 26
rect 39 21 42 25
rect 46 21 47 25
rect 39 20 47 21
rect 39 17 44 20
rect 4 12 11 17
rect 4 8 6 12
rect 10 8 11 12
rect 4 7 11 8
<< pdiffusion >>
rect 10 70 15 78
rect 7 69 15 70
rect 7 65 8 69
rect 12 65 15 69
rect 7 61 15 65
rect 7 57 8 61
rect 12 57 15 61
rect 7 56 15 57
rect 17 56 23 78
rect 25 73 35 78
rect 25 72 37 73
rect 25 68 28 72
rect 32 68 37 72
rect 25 56 37 68
rect 39 70 44 73
rect 39 69 47 70
rect 39 65 42 69
rect 46 65 47 69
rect 39 61 47 65
rect 39 57 42 61
rect 46 57 47 61
rect 39 56 47 57
<< metal1 >>
rect -2 96 52 100
rect -2 92 8 96
rect 12 92 18 96
rect 22 92 52 96
rect -2 88 52 92
rect 8 69 12 73
rect 8 61 12 65
rect 18 63 22 73
rect 28 72 32 88
rect 28 67 32 68
rect 42 69 46 70
rect 18 57 32 63
rect 8 23 12 57
rect 18 44 22 53
rect 28 51 32 57
rect 42 61 46 65
rect 28 47 33 51
rect 37 47 38 51
rect 16 42 22 44
rect 20 38 22 42
rect 42 41 46 57
rect 18 32 22 38
rect 26 37 27 41
rect 31 37 46 41
rect 18 27 33 32
rect 42 25 46 37
rect 8 22 22 23
rect 8 18 18 22
rect 8 17 22 18
rect 30 22 34 23
rect 42 20 46 21
rect 30 12 34 18
rect -2 8 6 12
rect 10 8 52 12
rect -2 4 18 8
rect 22 4 28 8
rect 32 4 52 8
rect -2 0 52 4
<< ntransistor >>
rect 13 17 15 23
rect 25 17 27 23
rect 37 17 39 26
<< ptransistor >>
rect 15 56 17 78
rect 23 56 25 78
rect 37 56 39 73
<< polycontact >>
rect 16 38 20 42
rect 33 47 37 51
rect 27 37 31 41
<< ndcontact >>
rect 18 18 22 22
rect 30 18 34 22
rect 42 21 46 25
rect 6 8 10 12
<< pdcontact >>
rect 8 65 12 69
rect 8 57 12 61
rect 28 68 32 72
rect 42 65 46 69
rect 42 57 46 61
<< psubstratepcontact >>
rect 18 4 22 8
rect 28 4 32 8
<< nsubstratencontact >>
rect 8 92 12 96
rect 18 92 22 96
<< psubstratepdiff >>
rect 17 8 33 9
rect 17 4 18 8
rect 22 4 28 8
rect 32 4 33 8
rect 17 3 33 4
<< nsubstratendiff >>
rect 7 96 23 97
rect 7 92 8 96
rect 12 92 18 96
rect 22 92 23 96
rect 7 91 23 92
<< labels >>
rlabel polycontact 28 39 28 39 6 an
rlabel ndcontact 20 20 20 20 6 z
rlabel metal1 10 45 10 45 6 z
rlabel metal1 20 40 20 40 6 b
rlabel metal1 20 65 20 65 6 a
rlabel metal1 25 6 25 6 6 vss
rlabel metal1 30 30 30 30 6 b
rlabel metal1 30 55 30 55 6 a
rlabel metal1 25 94 25 94 6 vdd
rlabel metal1 36 39 36 39 6 an
rlabel metal1 44 45 44 45 6 an
<< end >>
