.subckt cgi2v0x1 a b c vdd vss z
*   SPICE3 file   created from cgi2v0x1.ext -      technology: scmos
m00 vdd    a      n1     vdd p w=27u  l=2.3636u ad=135p     pd=46u      as=125.667p ps=46u
m01 w1     a      vdd    vdd p w=27u  l=2.3636u ad=67.5p    pd=32u      as=135p     ps=46u
m02 z      b      w1     vdd p w=27u  l=2.3636u ad=108p     pd=35u      as=67.5p    ps=32u
m03 n1     c      z      vdd p w=27u  l=2.3636u ad=125.667p pd=46u      as=108p     ps=35u
m04 vdd    b      n1     vdd p w=27u  l=2.3636u ad=135p     pd=46u      as=125.667p ps=46u
m05 vss    a      n3     vss n w=12u  l=2.3636u ad=94p      pd=35.3333u as=56p      ps=26u
m06 w2     a      vss    vss n w=12u  l=2.3636u ad=30p      pd=17u      as=94p      ps=35.3333u
m07 z      b      w2     vss n w=12u  l=2.3636u ad=48p      pd=20u      as=30p      ps=17u
m08 n3     c      z      vss n w=12u  l=2.3636u ad=56p      pd=26u      as=48p      ps=20u
m09 vss    b      n3     vss n w=12u  l=2.3636u ad=94p      pd=35.3333u as=56p      ps=26u
C0  a      vdd    0.022f
C1  vss    c      0.082f
C2  n3     b      0.013f
C3  z      n1     0.191f
C4  n3     vdd    0.005f
C5  z      b      0.119f
C6  vss    a      0.020f
C7  w2     n3     0.006f
C8  z      vdd    0.062f
C9  n1     b      0.082f
C10 n3     vss    0.337f
C11 w2     z      0.008f
C12 c      a      0.043f
C13 n1     vdd    0.405f
C14 vss    z      0.068f
C15 b      vdd    0.044f
C16 z      w1     0.007f
C17 n3     c      0.097f
C18 vss    n1     0.018f
C19 z      c      0.116f
C20 vss    b      0.033f
C21 w1     n1     0.023f
C22 n3     a      0.041f
C23 vss    vdd    0.004f
C24 n1     c      0.026f
C25 z      a      0.098f
C26 n1     a      0.042f
C27 c      b      0.232f
C28 w1     vdd    0.004f
C29 n3     z      0.177f
C30 b      a      0.125f
C31 c      vdd    0.025f
C32 n3     n1     0.038f
C33 n3     vss    0.003f
C35 z      vss    0.003f
C36 c      vss    0.019f
C37 b      vss    0.040f
C38 a      vss    0.042f
.ends
