magic
tech scmos
timestamp 1179385909
<< checkpaint >>
rect -22 -25 46 105
<< ab >>
rect 0 0 24 80
<< pwell >>
rect -4 -7 28 36
<< nwell >>
rect -4 36 28 87
<< polysilicon >>
rect 9 61 11 65
rect 9 39 11 42
rect 9 38 15 39
rect 9 34 10 38
rect 14 34 15 38
rect 9 33 15 34
rect 9 30 11 33
rect 9 6 11 11
<< ndiffusion >>
rect 2 29 9 30
rect 2 25 3 29
rect 7 25 9 29
rect 2 22 9 25
rect 2 18 3 22
rect 7 18 9 22
rect 2 17 9 18
rect 4 11 9 17
rect 11 23 19 30
rect 11 19 13 23
rect 17 19 19 23
rect 11 16 19 19
rect 11 12 13 16
rect 17 12 19 16
rect 11 11 19 12
<< pdiffusion >>
rect 13 62 19 63
rect 13 61 14 62
rect 4 56 9 61
rect 2 55 9 56
rect 2 51 3 55
rect 7 51 9 55
rect 2 48 9 51
rect 2 44 3 48
rect 7 44 9 48
rect 2 42 9 44
rect 11 58 14 61
rect 18 58 19 62
rect 11 42 19 58
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect -2 68 26 78
rect 13 62 19 68
rect 13 58 14 62
rect 18 58 19 62
rect 2 51 3 55
rect 7 51 14 55
rect 2 49 14 51
rect 2 48 7 49
rect 2 44 3 48
rect 2 43 7 44
rect 2 30 6 43
rect 18 39 22 47
rect 10 38 22 39
rect 14 34 22 38
rect 10 33 22 34
rect 2 29 7 30
rect 2 25 3 29
rect 2 22 7 25
rect 2 18 3 22
rect 2 17 7 18
rect 12 19 13 23
rect 17 19 18 23
rect 12 16 18 19
rect 12 12 13 16
rect 17 12 18 16
rect -2 2 26 12
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
<< ntransistor >>
rect 9 11 11 30
<< ptransistor >>
rect 9 42 11 61
<< polycontact >>
rect 10 34 14 38
<< ndcontact >>
rect 3 25 7 29
rect 3 18 7 22
rect 13 19 17 23
rect 13 12 17 16
<< pdcontact >>
rect 3 51 7 55
rect 3 44 7 48
rect 14 58 18 62
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
<< psubstratepdiff >>
rect 0 2 24 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 24 2
rect 0 -3 24 -2
<< nsubstratendiff >>
rect 0 82 24 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 24 82
rect 0 77 24 78
<< labels >>
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 6 12 6 6 vss
rlabel polycontact 12 36 12 36 6 a
rlabel metal1 12 52 12 52 6 z
rlabel metal1 12 74 12 74 6 vdd
rlabel metal1 20 40 20 40 6 a
<< end >>
