magic
tech scmos
timestamp 1179386424
<< checkpaint >>
rect -22 -22 118 94
<< ab >>
rect 0 0 96 72
<< pwell >>
rect -4 -4 100 32
<< nwell >>
rect -4 32 100 76
<< polysilicon >>
rect 9 66 11 70
rect 19 66 21 70
rect 29 66 31 70
rect 39 66 41 70
rect 49 66 51 70
rect 59 66 61 70
rect 70 53 72 58
rect 80 53 82 58
rect 9 35 11 40
rect 19 35 21 40
rect 29 35 31 40
rect 39 35 41 40
rect 49 35 51 40
rect 9 34 15 35
rect 9 30 10 34
rect 14 30 15 34
rect 9 29 15 30
rect 19 34 31 35
rect 19 30 26 34
rect 30 30 31 34
rect 19 29 31 30
rect 35 34 51 35
rect 35 30 36 34
rect 40 33 51 34
rect 59 35 61 40
rect 70 35 72 40
rect 80 35 82 40
rect 59 34 72 35
rect 40 30 41 33
rect 35 29 41 30
rect 59 30 60 34
rect 64 33 72 34
rect 76 34 82 35
rect 64 30 65 33
rect 59 29 65 30
rect 76 30 77 34
rect 81 30 82 34
rect 76 29 82 30
rect 12 26 14 29
rect 19 26 21 29
rect 29 26 31 29
rect 36 26 38 29
rect 12 2 14 7
rect 19 2 21 7
rect 29 2 31 7
rect 36 2 38 7
<< ndiffusion >>
rect 3 8 12 26
rect 3 4 5 8
rect 9 7 12 8
rect 14 7 19 26
rect 21 18 29 26
rect 21 14 23 18
rect 27 14 29 18
rect 21 7 29 14
rect 31 7 36 26
rect 38 8 47 26
rect 38 7 41 8
rect 9 4 10 7
rect 3 3 10 4
rect 40 4 41 7
rect 45 4 47 8
rect 40 3 47 4
<< pdiffusion >>
rect 2 65 9 66
rect 2 61 3 65
rect 7 61 9 65
rect 2 58 9 61
rect 2 54 3 58
rect 7 54 9 58
rect 2 40 9 54
rect 11 57 19 66
rect 11 53 13 57
rect 17 53 19 57
rect 11 50 19 53
rect 11 46 13 50
rect 17 46 19 50
rect 11 40 19 46
rect 21 65 29 66
rect 21 61 23 65
rect 27 61 29 65
rect 21 58 29 61
rect 21 54 23 58
rect 27 54 29 58
rect 21 40 29 54
rect 31 58 39 66
rect 31 54 33 58
rect 37 54 39 58
rect 31 50 39 54
rect 31 46 33 50
rect 37 46 39 50
rect 31 40 39 46
rect 41 65 49 66
rect 41 61 43 65
rect 47 61 49 65
rect 41 58 49 61
rect 41 54 43 58
rect 47 54 49 58
rect 41 40 49 54
rect 51 58 59 66
rect 51 54 53 58
rect 57 54 59 58
rect 51 50 59 54
rect 51 46 53 50
rect 57 46 59 50
rect 51 40 59 46
rect 61 65 68 66
rect 61 61 63 65
rect 67 61 68 65
rect 61 58 68 61
rect 61 54 63 58
rect 67 54 68 58
rect 61 53 68 54
rect 61 40 70 53
rect 72 52 80 53
rect 72 48 74 52
rect 78 48 80 52
rect 72 45 80 48
rect 72 41 74 45
rect 78 41 80 45
rect 72 40 80 41
rect 82 52 90 53
rect 82 48 84 52
rect 88 48 90 52
rect 82 40 90 48
<< metal1 >>
rect -2 68 98 72
rect -2 65 76 68
rect -2 64 3 65
rect 2 61 3 64
rect 7 64 23 65
rect 7 61 8 64
rect 2 58 8 61
rect 22 61 23 64
rect 27 64 43 65
rect 27 61 28 64
rect 22 58 28 61
rect 42 61 43 64
rect 47 64 63 65
rect 47 61 48 64
rect 2 54 3 58
rect 7 54 8 58
rect 13 57 17 58
rect 22 54 23 58
rect 27 54 28 58
rect 33 58 38 59
rect 37 54 38 58
rect 42 58 48 61
rect 62 61 63 64
rect 67 64 76 65
rect 80 64 84 68
rect 88 64 98 68
rect 67 61 68 64
rect 42 54 43 58
rect 47 54 48 58
rect 53 58 57 59
rect 62 58 68 61
rect 62 54 63 58
rect 67 54 68 58
rect 13 50 17 53
rect 33 50 38 54
rect 53 50 57 54
rect 74 52 78 53
rect 2 46 13 50
rect 17 46 33 50
rect 37 46 53 50
rect 57 48 74 50
rect 57 46 78 48
rect 84 52 88 64
rect 84 47 88 48
rect 2 18 6 46
rect 74 45 78 46
rect 25 38 49 42
rect 74 40 78 41
rect 10 34 14 35
rect 25 34 31 38
rect 45 34 49 38
rect 25 30 26 34
rect 30 30 31 34
rect 35 30 36 34
rect 40 30 41 34
rect 45 30 60 34
rect 64 30 65 34
rect 73 30 77 34
rect 81 30 87 34
rect 10 26 14 30
rect 35 26 41 30
rect 73 26 79 30
rect 10 22 79 26
rect 2 14 23 18
rect 27 14 31 18
rect -2 4 5 8
rect 9 4 41 8
rect 45 4 76 8
rect 80 4 84 8
rect 88 4 98 8
rect -2 0 98 4
<< ntransistor >>
rect 12 7 14 26
rect 19 7 21 26
rect 29 7 31 26
rect 36 7 38 26
<< ptransistor >>
rect 9 40 11 66
rect 19 40 21 66
rect 29 40 31 66
rect 39 40 41 66
rect 49 40 51 66
rect 59 40 61 66
rect 70 40 72 53
rect 80 40 82 53
<< polycontact >>
rect 10 30 14 34
rect 26 30 30 34
rect 36 30 40 34
rect 60 30 64 34
rect 77 30 81 34
<< ndcontact >>
rect 5 4 9 8
rect 23 14 27 18
rect 41 4 45 8
<< pdcontact >>
rect 3 61 7 65
rect 3 54 7 58
rect 13 53 17 57
rect 13 46 17 50
rect 23 61 27 65
rect 23 54 27 58
rect 33 54 37 58
rect 33 46 37 50
rect 43 61 47 65
rect 43 54 47 58
rect 53 54 57 58
rect 53 46 57 50
rect 63 61 67 65
rect 63 54 67 58
rect 74 48 78 52
rect 74 41 78 45
rect 84 48 88 52
<< psubstratepcontact >>
rect 76 4 80 8
rect 84 4 88 8
<< nsubstratencontact >>
rect 76 64 80 68
rect 84 64 88 68
<< psubstratepdiff >>
rect 75 8 89 24
rect 75 4 76 8
rect 80 4 84 8
rect 88 4 89 8
rect 75 3 89 4
<< nsubstratendiff >>
rect 75 68 89 69
rect 75 64 76 68
rect 80 64 84 68
rect 88 64 89 68
rect 75 61 89 64
<< labels >>
rlabel metal1 12 16 12 16 6 z
rlabel polycontact 12 32 12 32 6 a
rlabel metal1 4 32 4 32 6 z
rlabel metal1 12 48 12 48 6 z
rlabel metal1 28 16 28 16 6 z
rlabel metal1 20 16 20 16 6 z
rlabel metal1 20 24 20 24 6 a
rlabel metal1 28 24 28 24 6 a
rlabel polycontact 28 32 28 32 6 b
rlabel metal1 28 36 28 36 6 b
rlabel metal1 20 48 20 48 6 z
rlabel metal1 28 48 28 48 6 z
rlabel metal1 48 4 48 4 6 vss
rlabel metal1 36 24 36 24 6 a
rlabel metal1 44 24 44 24 6 a
rlabel metal1 52 24 52 24 6 a
rlabel metal1 52 32 52 32 6 b
rlabel metal1 36 40 36 40 6 b
rlabel metal1 44 40 44 40 6 b
rlabel metal1 36 52 36 52 6 z
rlabel metal1 44 48 44 48 6 z
rlabel metal1 52 48 52 48 6 z
rlabel metal1 48 68 48 68 6 vdd
rlabel metal1 60 24 60 24 6 a
rlabel metal1 68 24 68 24 6 a
rlabel metal1 76 28 76 28 6 a
rlabel metal1 60 32 60 32 6 b
rlabel metal1 60 48 60 48 6 z
rlabel metal1 68 48 68 48 6 z
rlabel metal1 76 48 76 48 6 z
rlabel metal1 84 32 84 32 6 a
<< end >>
