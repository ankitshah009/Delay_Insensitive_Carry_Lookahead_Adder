magic
tech scmos
timestamp 1179385619
<< checkpaint >>
rect -22 -22 134 94
<< ab >>
rect 0 0 112 72
<< pwell >>
rect -4 -4 116 32
<< nwell >>
rect -4 32 116 76
<< polysilicon >>
rect 25 68 110 70
rect 15 59 17 64
rect 25 60 27 68
rect 56 65 58 68
rect 35 60 37 64
rect 77 60 79 64
rect 87 60 89 68
rect 97 60 99 64
rect 56 40 58 43
rect 56 38 61 40
rect 15 35 17 38
rect 2 34 17 35
rect 2 30 3 34
rect 7 30 17 34
rect 25 35 27 38
rect 25 33 30 35
rect 2 29 17 30
rect 12 22 14 29
rect 28 27 30 33
rect 35 34 37 38
rect 59 36 61 38
rect 59 35 65 36
rect 77 35 79 38
rect 35 33 55 34
rect 35 32 50 33
rect 43 29 50 32
rect 54 29 55 33
rect 43 28 55 29
rect 59 31 60 35
rect 64 31 65 35
rect 59 30 65 31
rect 73 34 79 35
rect 73 30 74 34
rect 78 30 79 34
rect 87 33 89 38
rect 97 35 99 38
rect 94 33 99 35
rect 22 22 24 27
rect 28 25 34 27
rect 32 22 34 25
rect 12 7 14 12
rect 22 4 24 12
rect 32 8 34 12
rect 43 4 45 28
rect 59 26 61 30
rect 73 29 79 30
rect 94 29 96 33
rect 108 29 110 68
rect 73 27 83 29
rect 81 24 83 27
rect 91 27 96 29
rect 101 27 110 29
rect 91 24 93 27
rect 101 24 103 27
rect 59 11 61 16
rect 81 9 83 14
rect 91 4 93 14
rect 101 9 103 14
rect 22 2 93 4
<< ndiffusion >>
rect 3 17 12 22
rect 3 13 5 17
rect 9 13 12 17
rect 3 12 12 13
rect 14 21 22 22
rect 14 17 16 21
rect 20 17 22 21
rect 14 12 22 17
rect 24 21 32 22
rect 24 17 26 21
rect 30 17 32 21
rect 24 12 32 17
rect 34 19 39 22
rect 34 18 41 19
rect 34 14 36 18
rect 40 14 41 18
rect 34 12 41 14
rect 52 25 59 26
rect 52 21 53 25
rect 57 21 59 25
rect 52 20 59 21
rect 54 16 59 20
rect 61 24 66 26
rect 61 19 81 24
rect 61 16 71 19
rect 63 15 71 16
rect 75 15 81 19
rect 63 14 81 15
rect 83 23 91 24
rect 83 19 85 23
rect 89 19 91 23
rect 83 14 91 19
rect 93 19 101 24
rect 93 15 95 19
rect 99 15 101 19
rect 93 14 101 15
rect 103 23 110 24
rect 103 19 105 23
rect 109 19 110 23
rect 103 18 110 19
rect 103 14 108 18
<< pdiffusion >>
rect 20 59 25 60
rect 7 58 15 59
rect 7 54 9 58
rect 13 54 15 58
rect 7 51 15 54
rect 7 47 9 51
rect 13 47 15 51
rect 7 38 15 47
rect 17 50 25 59
rect 17 46 19 50
rect 23 46 25 50
rect 17 43 25 46
rect 17 39 19 43
rect 23 39 25 43
rect 17 38 25 39
rect 27 50 35 60
rect 27 46 29 50
rect 33 46 35 50
rect 27 43 35 46
rect 27 39 29 43
rect 33 39 35 43
rect 27 38 35 39
rect 37 51 42 60
rect 37 50 44 51
rect 37 46 39 50
rect 43 46 44 50
rect 51 49 56 65
rect 37 43 44 46
rect 49 48 56 49
rect 49 44 50 48
rect 54 44 56 48
rect 49 43 56 44
rect 58 64 75 65
rect 58 60 63 64
rect 67 60 75 64
rect 58 43 77 60
rect 37 39 39 43
rect 43 39 44 43
rect 37 38 44 39
rect 67 38 77 43
rect 79 50 87 60
rect 79 46 81 50
rect 85 46 87 50
rect 79 43 87 46
rect 79 39 81 43
rect 85 39 87 43
rect 79 38 87 39
rect 89 50 97 60
rect 89 46 91 50
rect 95 46 97 50
rect 89 43 97 46
rect 89 39 91 43
rect 95 39 97 43
rect 89 38 97 39
rect 99 59 106 60
rect 99 55 101 59
rect 105 55 106 59
rect 99 52 106 55
rect 99 48 101 52
rect 105 48 106 52
rect 99 47 106 48
rect 99 38 104 47
<< metal1 >>
rect -2 68 114 72
rect -2 64 4 68
rect 8 64 114 68
rect 9 58 13 64
rect 62 60 63 64
rect 67 60 68 64
rect 9 51 13 54
rect 9 46 13 47
rect 19 57 52 59
rect 72 57 101 59
rect 19 55 101 57
rect 105 55 106 59
rect 19 50 23 55
rect 48 53 76 55
rect 100 52 106 55
rect 19 43 23 46
rect 2 37 14 43
rect 2 34 7 37
rect 19 34 23 39
rect 2 30 3 34
rect 2 21 7 30
rect 16 30 23 34
rect 26 50 33 51
rect 26 46 29 50
rect 26 43 33 46
rect 26 39 29 43
rect 26 38 33 39
rect 39 50 43 51
rect 81 50 85 51
rect 39 43 43 46
rect 16 21 20 30
rect 4 13 5 17
rect 9 13 10 17
rect 16 16 20 17
rect 26 27 30 38
rect 39 35 43 39
rect 50 48 54 49
rect 65 46 78 50
rect 39 31 46 35
rect 26 21 38 27
rect 42 18 46 31
rect 50 33 54 44
rect 57 35 63 42
rect 57 31 60 35
rect 64 31 70 35
rect 57 29 70 31
rect 74 34 78 46
rect 74 29 78 30
rect 81 43 85 46
rect 50 25 54 29
rect 81 26 85 39
rect 90 50 95 51
rect 90 46 91 50
rect 100 48 101 52
rect 90 43 95 46
rect 90 39 91 43
rect 90 35 95 39
rect 90 29 102 35
rect 50 21 53 25
rect 57 21 58 25
rect 62 23 89 26
rect 62 22 85 23
rect 62 18 66 22
rect 98 19 102 29
rect 26 13 30 17
rect 35 14 36 18
rect 40 14 66 18
rect 70 15 71 19
rect 75 15 76 19
rect 85 18 89 19
rect 4 8 10 13
rect 47 8 48 11
rect -2 7 48 8
rect 52 8 53 11
rect 70 8 76 15
rect 94 15 95 19
rect 99 15 102 19
rect 105 23 109 52
rect 105 18 109 19
rect 94 13 102 15
rect 52 7 114 8
rect -2 0 114 7
<< ntransistor >>
rect 12 12 14 22
rect 22 12 24 22
rect 32 12 34 22
rect 59 16 61 26
rect 81 14 83 24
rect 91 14 93 24
rect 101 14 103 24
<< ptransistor >>
rect 15 38 17 59
rect 25 38 27 60
rect 35 38 37 60
rect 56 43 58 65
rect 77 38 79 60
rect 87 38 89 60
rect 97 38 99 60
<< polycontact >>
rect 3 30 7 34
rect 50 29 54 33
rect 60 31 64 35
rect 74 30 78 34
<< ndcontact >>
rect 5 13 9 17
rect 16 17 20 21
rect 26 17 30 21
rect 36 14 40 18
rect 53 21 57 25
rect 71 15 75 19
rect 85 19 89 23
rect 95 15 99 19
rect 105 19 109 23
<< pdcontact >>
rect 9 54 13 58
rect 9 47 13 51
rect 19 46 23 50
rect 19 39 23 43
rect 29 46 33 50
rect 29 39 33 43
rect 39 46 43 50
rect 50 44 54 48
rect 63 60 67 64
rect 39 39 43 43
rect 81 46 85 50
rect 81 39 85 43
rect 91 46 95 50
rect 91 39 95 43
rect 101 55 105 59
rect 101 48 105 52
<< psubstratepcontact >>
rect 48 7 52 11
<< nsubstratencontact >>
rect 4 64 8 68
<< psubstratepdiff >>
rect 47 11 53 12
rect 47 7 48 11
rect 52 7 53 11
rect 47 6 53 7
<< nsubstratendiff >>
rect 3 68 9 69
rect 3 64 4 68
rect 8 64 9 68
rect 3 63 9 64
<< labels >>
rlabel polysilicon 49 31 49 31 6 sn
rlabel polycontact 4 32 4 32 6 a0
rlabel metal1 18 25 18 25 6 a0n
rlabel metal1 12 40 12 40 6 a0
rlabel metal1 36 24 36 24 6 z0
rlabel metal1 28 32 28 32 6 z0
rlabel pdcontact 41 41 41 41 6 a1n
rlabel metal1 21 44 21 44 6 a0n
rlabel metal1 56 4 56 4 6 vss
rlabel metal1 50 16 50 16 6 a1n
rlabel metal1 60 36 60 36 6 s
rlabel metal1 52 35 52 35 6 sn
rlabel metal1 56 68 56 68 6 vdd
rlabel metal1 75 24 75 24 6 a1n
rlabel metal1 68 32 68 32 6 s
rlabel metal1 76 36 76 36 6 a1
rlabel metal1 83 36 83 36 6 a1n
rlabel metal1 68 48 68 48 6 a1
rlabel metal1 100 24 100 24 6 z1
rlabel pdcontact 92 40 92 40 6 z1
rlabel metal1 107 35 107 35 6 a0n
rlabel metal1 89 57 89 57 6 a0n
<< end >>
