.subckt a2_x4 i0 i1 q vdd vss
*   SPICE3 file   created from a2_x4.ext -      technology: scmos
m00 w1     i0     vdd    vdd p w=20u  l=2.3636u ad=101.5p   pd=31u      as=146.78p  ps=44.4068u
m01 vdd    i1     w1     vdd p w=20u  l=2.3636u ad=146.78p  pd=44.4068u as=101.5p   ps=31u
m02 q      w1     vdd    vdd p w=39u  l=2.3636u ad=195p     pd=49u      as=286.22p  ps=86.5932u
m03 vdd    w1     q      vdd p w=39u  l=2.3636u ad=286.22p  pd=86.5932u as=195p     ps=49u
m04 w2     i0     w1     vss n w=18u  l=2.3636u ad=90p      pd=28u      as=144p     ps=52u
m05 vss    i1     w2     vss n w=18u  l=2.3636u ad=108.321p pd=36u      as=90p      ps=28u
m06 q      w1     vss    vss n w=19u  l=2.3636u ad=95p      pd=29u      as=114.339p ps=38u
m07 vss    w1     q      vss n w=19u  l=2.3636u ad=114.339p pd=38u      as=95p      ps=29u
C0  vdd    w1     0.085f
C1  vss    i1     0.063f
C2  w2     w1     0.019f
C3  q      i0     0.054f
C4  vss    vdd    0.004f
C5  i1     vdd    0.134f
C6  q      w1     0.121f
C7  i0     w1     0.323f
C8  w2     vss    0.019f
C9  vss    q      0.082f
C10 q      i1     0.334f
C11 vss    i0     0.013f
C12 q      vdd    0.168f
C13 i1     i0     0.130f
C14 vss    w1     0.123f
C15 i0     vdd    0.033f
C16 i1     w1     0.442f
C18 q      vss    0.014f
C19 i1     vss    0.039f
C20 i0     vss    0.034f
C22 w1     vss    0.066f
.ends
