magic
tech scmos
timestamp 1185094714
<< checkpaint >>
rect -22 -22 62 122
<< ab >>
rect 0 0 40 100
<< pwell >>
rect -4 -4 44 48
<< nwell >>
rect -4 48 44 104
<< polysilicon >>
rect 13 94 15 98
rect 25 94 27 98
rect 13 53 15 56
rect 25 53 27 56
rect 13 52 27 53
rect 13 48 20 52
rect 24 48 27 52
rect 13 47 27 48
rect 13 36 15 47
rect 25 36 27 47
rect 13 12 15 17
rect 25 12 27 17
<< ndiffusion >>
rect 4 32 13 36
rect 4 28 6 32
rect 10 28 13 32
rect 4 22 13 28
rect 4 18 6 22
rect 10 18 13 22
rect 4 17 13 18
rect 15 32 25 36
rect 15 28 18 32
rect 22 28 25 32
rect 15 22 25 28
rect 15 18 18 22
rect 22 18 25 22
rect 15 17 25 18
rect 27 32 36 36
rect 27 28 30 32
rect 34 28 36 32
rect 27 22 36 28
rect 27 18 30 22
rect 34 18 36 22
rect 27 17 36 18
<< pdiffusion >>
rect 4 92 13 94
rect 4 88 6 92
rect 10 88 13 92
rect 4 82 13 88
rect 4 78 6 82
rect 10 78 13 82
rect 4 72 13 78
rect 4 68 6 72
rect 10 68 13 72
rect 4 56 13 68
rect 15 72 25 94
rect 15 68 18 72
rect 22 68 25 72
rect 15 62 25 68
rect 15 58 18 62
rect 22 58 25 62
rect 15 56 25 58
rect 27 92 36 94
rect 27 88 30 92
rect 34 88 36 92
rect 27 82 36 88
rect 27 78 30 82
rect 34 78 36 82
rect 27 72 36 78
rect 27 68 30 72
rect 34 68 36 72
rect 27 56 36 68
<< metal1 >>
rect -2 92 42 100
rect -2 88 6 92
rect 10 88 30 92
rect 34 88 42 92
rect 6 82 10 88
rect 6 72 10 78
rect 30 82 34 88
rect 6 67 10 68
rect 18 72 22 73
rect 18 63 22 68
rect 30 72 34 78
rect 30 67 34 68
rect 8 62 22 63
rect 8 58 18 62
rect 8 57 22 58
rect 8 43 12 57
rect 28 52 32 63
rect 17 48 20 52
rect 24 48 32 52
rect 8 37 22 43
rect 28 37 32 48
rect 6 32 10 33
rect 6 22 10 28
rect 6 12 10 18
rect 18 32 22 37
rect 18 22 22 28
rect 18 17 22 18
rect 30 32 34 33
rect 30 22 34 28
rect 30 12 34 18
rect -2 8 42 12
rect -2 4 8 8
rect 12 4 18 8
rect 22 4 42 8
rect -2 0 42 4
<< ntransistor >>
rect 13 17 15 36
rect 25 17 27 36
<< ptransistor >>
rect 13 56 15 94
rect 25 56 27 94
<< polycontact >>
rect 20 48 24 52
<< ndcontact >>
rect 6 28 10 32
rect 6 18 10 22
rect 18 28 22 32
rect 18 18 22 22
rect 30 28 34 32
rect 30 18 34 22
<< pdcontact >>
rect 6 88 10 92
rect 6 78 10 82
rect 6 68 10 72
rect 18 68 22 72
rect 18 58 22 62
rect 30 88 34 92
rect 30 78 34 82
rect 30 68 34 72
<< psubstratepcontact >>
rect 8 4 12 8
rect 18 4 22 8
<< psubstratepdiff >>
rect 7 8 23 9
rect 7 4 8 8
rect 12 4 18 8
rect 22 4 23 8
rect 7 3 23 4
<< labels >>
rlabel metal1 10 50 10 50 6 z
rlabel psubstratepcontact 20 6 20 6 6 vss
rlabel ndcontact 20 30 20 30 6 z
rlabel metal1 20 50 20 50 6 a
rlabel metal1 20 65 20 65 6 z
rlabel metal1 20 94 20 94 6 vdd
rlabel metal1 30 50 30 50 6 a
<< end >>
