magic
tech scmos
timestamp 1185094678
<< checkpaint >>
rect -22 -22 102 122
<< ab >>
rect 0 0 80 100
<< pwell >>
rect -4 -4 84 48
<< nwell >>
rect -4 48 84 104
<< polysilicon >>
rect 11 83 13 88
rect 23 83 25 88
rect 31 83 33 88
rect 43 83 45 88
rect 55 83 57 88
rect 67 83 69 88
rect 11 53 13 63
rect 23 53 25 63
rect 11 52 27 53
rect 11 48 16 52
rect 20 48 27 52
rect 11 47 27 48
rect 13 26 15 47
rect 25 33 27 47
rect 31 42 33 63
rect 43 54 45 63
rect 43 53 49 54
rect 43 49 44 53
rect 48 49 49 53
rect 43 48 49 49
rect 31 41 41 42
rect 31 37 36 41
rect 40 37 41 41
rect 31 36 41 37
rect 33 33 35 36
rect 45 33 47 48
rect 55 42 57 63
rect 67 52 69 57
rect 63 51 69 52
rect 63 47 64 51
rect 68 47 69 51
rect 63 46 69 47
rect 53 41 59 42
rect 53 37 54 41
rect 58 37 59 41
rect 67 37 69 46
rect 53 36 59 37
rect 57 33 59 36
rect 25 19 27 24
rect 33 19 35 24
rect 45 19 47 24
rect 57 19 59 24
rect 13 12 15 17
rect 67 19 69 24
<< ndiffusion >>
rect 61 33 67 37
rect 17 26 25 33
rect 8 23 13 26
rect 5 22 13 23
rect 5 18 6 22
rect 10 18 13 22
rect 5 17 13 18
rect 15 24 25 26
rect 27 24 33 33
rect 35 32 45 33
rect 35 28 38 32
rect 42 28 45 32
rect 35 24 45 28
rect 47 29 57 33
rect 47 25 50 29
rect 54 25 57 29
rect 47 24 57 25
rect 59 24 67 33
rect 69 36 77 37
rect 69 32 72 36
rect 76 32 77 36
rect 69 31 77 32
rect 69 24 74 31
rect 15 17 23 24
rect 17 12 23 17
rect 17 8 18 12
rect 22 8 23 12
rect 61 17 65 24
rect 61 16 67 17
rect 61 12 62 16
rect 66 12 67 16
rect 61 11 67 12
rect 17 7 23 8
<< pdiffusion >>
rect 3 82 11 83
rect 3 78 4 82
rect 8 78 11 82
rect 3 74 11 78
rect 3 70 4 74
rect 8 70 11 74
rect 3 69 11 70
rect 6 63 11 69
rect 13 82 23 83
rect 13 78 16 82
rect 20 78 23 82
rect 13 63 23 78
rect 25 63 31 83
rect 33 72 43 83
rect 33 68 36 72
rect 40 68 43 72
rect 33 63 43 68
rect 45 82 55 83
rect 45 78 48 82
rect 52 78 55 82
rect 45 63 55 78
rect 57 82 67 83
rect 57 78 60 82
rect 64 78 67 82
rect 57 63 67 78
rect 59 57 67 63
rect 69 63 74 83
rect 69 62 77 63
rect 69 58 72 62
rect 76 58 77 62
rect 69 57 77 58
<< metal1 >>
rect -2 96 82 100
rect -2 92 8 96
rect 12 92 18 96
rect 22 92 82 96
rect -2 88 82 92
rect 4 82 8 83
rect 4 74 8 78
rect 16 82 20 88
rect 60 82 64 88
rect 16 77 20 78
rect 26 78 48 82
rect 52 78 53 82
rect 26 72 30 78
rect 60 77 64 78
rect 8 70 30 72
rect 4 68 30 70
rect 36 72 42 73
rect 40 68 42 72
rect 36 63 42 68
rect 8 53 12 63
rect 28 57 42 63
rect 8 52 22 53
rect 8 48 16 52
rect 20 48 22 52
rect 8 47 22 48
rect 8 37 12 47
rect 28 32 32 57
rect 38 49 44 53
rect 48 49 52 73
rect 38 47 52 49
rect 58 67 72 73
rect 58 52 62 67
rect 72 62 76 63
rect 58 51 68 52
rect 58 47 64 51
rect 58 46 68 47
rect 72 42 76 58
rect 36 41 76 42
rect 40 37 54 41
rect 58 37 76 41
rect 36 36 76 37
rect 28 28 38 32
rect 42 28 43 32
rect 72 31 76 32
rect 28 27 43 28
rect 49 25 50 29
rect 54 25 55 29
rect 49 22 55 25
rect 5 18 6 22
rect 10 18 55 22
rect 62 16 66 17
rect -2 8 18 12
rect 22 8 82 12
rect -2 4 38 8
rect 42 4 48 8
rect 52 4 82 8
rect -2 0 82 4
<< ntransistor >>
rect 13 17 15 26
rect 25 24 27 33
rect 33 24 35 33
rect 45 24 47 33
rect 57 24 59 33
rect 67 24 69 37
<< ptransistor >>
rect 11 63 13 83
rect 23 63 25 83
rect 31 63 33 83
rect 43 63 45 83
rect 55 63 57 83
rect 67 57 69 83
<< polycontact >>
rect 16 48 20 52
rect 44 49 48 53
rect 36 37 40 41
rect 64 47 68 51
rect 54 37 58 41
<< ndcontact >>
rect 6 18 10 22
rect 38 28 42 32
rect 50 25 54 29
rect 72 32 76 36
rect 18 8 22 12
rect 62 12 66 16
<< pdcontact >>
rect 4 78 8 82
rect 4 70 8 74
rect 16 78 20 82
rect 36 68 40 72
rect 48 78 52 82
rect 60 78 64 82
rect 72 58 76 62
<< psubstratepcontact >>
rect 38 4 42 8
rect 48 4 52 8
<< nsubstratencontact >>
rect 8 92 12 96
rect 18 92 22 96
<< psubstratepdiff >>
rect 37 8 53 9
rect 37 4 38 8
rect 42 4 48 8
rect 52 4 53 8
rect 37 3 53 4
<< nsubstratendiff >>
rect 7 96 23 97
rect 7 92 8 96
rect 12 92 18 96
rect 22 92 23 96
rect 7 91 23 92
<< labels >>
rlabel polysilicon 36 39 36 39 6 an
rlabel polycontact 56 39 56 39 6 an
rlabel metal1 10 50 10 50 6 b
rlabel metal1 6 75 6 75 6 n2
rlabel metal1 20 50 20 50 6 b
rlabel psubstratepcontact 40 6 40 6 6 vss
rlabel ndcontact 40 30 40 30 6 z
rlabel metal1 30 45 30 45 6 z
rlabel metal1 40 50 40 50 6 c
rlabel metal1 40 65 40 65 6 z
rlabel metal1 40 94 40 94 6 vdd
rlabel metal1 52 23 52 23 6 n4
rlabel metal1 30 20 30 20 6 n4
rlabel metal1 60 60 60 60 6 a
rlabel metal1 50 60 50 60 6 c
rlabel metal1 39 80 39 80 6 n2
rlabel polycontact 56 39 56 39 6 an
rlabel metal1 74 47 74 47 6 an
rlabel metal1 70 70 70 70 6 a
<< end >>
