magic
tech scmos
timestamp 1179387215
<< checkpaint >>
rect -22 -25 78 105
<< ab >>
rect 0 0 56 80
<< pwell >>
rect -4 -7 60 36
<< nwell >>
rect -4 36 60 87
<< polysilicon >>
rect 24 69 26 74
rect 31 69 33 74
rect 38 69 40 74
rect 13 61 15 67
rect 13 46 15 49
rect 9 45 15 46
rect 9 41 10 45
rect 14 41 15 45
rect 9 40 15 41
rect 9 22 11 40
rect 24 39 26 44
rect 19 38 26 39
rect 19 34 20 38
rect 24 36 26 38
rect 24 34 25 36
rect 19 33 25 34
rect 19 22 21 33
rect 31 31 33 44
rect 38 41 40 44
rect 38 40 47 41
rect 38 39 42 40
rect 41 36 42 39
rect 46 36 47 40
rect 41 35 47 36
rect 29 30 36 31
rect 29 26 31 30
rect 35 26 36 30
rect 29 25 36 26
rect 29 22 31 25
rect 41 22 43 35
rect 9 11 11 16
rect 19 11 21 16
rect 29 11 31 16
rect 41 11 43 16
<< ndiffusion >>
rect 2 21 9 22
rect 2 17 3 21
rect 7 17 9 21
rect 2 16 9 17
rect 11 21 19 22
rect 11 17 13 21
rect 17 17 19 21
rect 11 16 19 17
rect 21 21 29 22
rect 21 17 23 21
rect 27 17 29 21
rect 21 16 29 17
rect 31 16 41 22
rect 43 21 50 22
rect 43 17 45 21
rect 49 17 50 21
rect 43 16 50 17
rect 33 12 39 16
rect 33 8 34 12
rect 38 8 39 12
rect 33 7 39 8
<< pdiffusion >>
rect 17 68 24 69
rect 17 64 18 68
rect 22 64 24 68
rect 17 61 24 64
rect 6 60 13 61
rect 6 56 7 60
rect 11 56 13 60
rect 6 55 13 56
rect 8 49 13 55
rect 15 49 24 61
rect 17 44 24 49
rect 26 44 31 69
rect 33 44 38 69
rect 40 64 45 69
rect 40 63 47 64
rect 40 59 42 63
rect 46 59 47 63
rect 40 58 47 59
rect 40 44 45 58
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect -2 68 58 78
rect 18 63 22 64
rect 2 60 15 62
rect 2 56 7 60
rect 11 56 15 60
rect 26 59 42 63
rect 46 59 47 63
rect 2 21 6 56
rect 26 55 30 59
rect 18 51 30 55
rect 18 48 22 51
rect 34 49 46 55
rect 10 45 22 48
rect 14 44 22 45
rect 10 29 14 41
rect 26 39 30 47
rect 42 40 46 49
rect 17 38 30 39
rect 17 34 20 38
rect 24 34 30 38
rect 34 30 38 39
rect 42 35 46 36
rect 10 25 26 29
rect 30 26 31 30
rect 35 26 47 30
rect 22 21 26 25
rect 2 17 3 21
rect 7 17 8 21
rect 12 17 13 21
rect 17 17 18 21
rect 22 17 23 21
rect 27 17 45 21
rect 49 17 50 21
rect 12 12 18 17
rect -2 8 34 12
rect 38 8 58 12
rect -2 2 58 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
<< ntransistor >>
rect 9 16 11 22
rect 19 16 21 22
rect 29 16 31 22
rect 41 16 43 22
<< ptransistor >>
rect 13 49 15 61
rect 24 44 26 69
rect 31 44 33 69
rect 38 44 40 69
<< polycontact >>
rect 10 41 14 45
rect 20 34 24 38
rect 42 36 46 40
rect 31 26 35 30
<< ndcontact >>
rect 3 17 7 21
rect 13 17 17 21
rect 23 17 27 21
rect 45 17 49 21
rect 34 8 38 12
<< pdcontact >>
rect 18 64 22 68
rect 7 56 11 60
rect 42 59 46 63
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
<< psubstratepdiff >>
rect 0 2 56 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 56 2
rect 0 -3 56 -2
<< nsubstratendiff >>
rect 0 82 56 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 56 82
rect 0 77 56 78
<< labels >>
rlabel polycontact 12 43 12 43 6 zn
rlabel metal1 4 36 4 36 6 z
rlabel metal1 20 36 20 36 6 a
rlabel metal1 12 36 12 36 6 zn
rlabel metal1 12 60 12 60 6 z
rlabel metal1 28 6 28 6 6 vss
rlabel metal1 36 32 36 32 6 b
rlabel metal1 28 44 28 44 6 a
rlabel metal1 36 52 36 52 6 c
rlabel metal1 28 74 28 74 6 vdd
rlabel metal1 36 19 36 19 6 zn
rlabel metal1 44 28 44 28 6 b
rlabel metal1 44 48 44 48 6 c
rlabel metal1 36 61 36 61 6 zn
<< end >>
