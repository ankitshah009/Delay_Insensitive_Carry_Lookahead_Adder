.subckt bf1_x8 a vdd vss z
*   SPICE3 file   created from bf1_x8.ext -      technology: scmos
m00 z      an     vdd    vdd p w=39u  l=2.3636u ad=195p     pd=52.7172u as=243.703p ps=66.8038u
m01 vdd    an     z      vdd p w=39u  l=2.3636u ad=243.703p pd=66.8038u as=195p     ps=52.7172u
m02 z      an     vdd    vdd p w=39u  l=2.3636u ad=195p     pd=52.7172u as=243.703p ps=66.8038u
m03 vdd    an     z      vdd p w=28u  l=2.3636u ad=174.967p pd=47.9617u as=140p     ps=37.8483u
m04 an     a      vdd    vdd p w=28u  l=2.3636u ad=140p     pd=40.25u   as=174.967p ps=47.9617u
m05 vdd    a      an     vdd p w=36u  l=2.3636u ad=224.957p pd=61.6651u as=180p     ps=51.75u
m06 z      an     vss    vss n w=18u  l=2.3636u ad=90p      pd=28u      as=111.462p ps=37.0385u
m07 vss    an     z      vss n w=18u  l=2.3636u ad=111.462p pd=37.0385u as=90p      ps=28u
m08 z      an     vss    vss n w=18u  l=2.3636u ad=90p      pd=28u      as=111.462p ps=37.0385u
m09 vss    an     z      vss n w=18u  l=2.3636u ad=111.462p pd=37.0385u as=90p      ps=28u
m10 an     a      vss    vss n w=16u  l=2.3636u ad=80p      pd=26u      as=99.0769p ps=32.9231u
m11 vss    a      an     vss n w=16u  l=2.3636u ad=99.0769p pd=32.9231u as=80p      ps=26u
C0  vss    z      0.451f
C1  vss    an     0.236f
C2  a      vdd    0.040f
C3  z      an     0.327f
C4  vss    a      0.047f
C5  vss    vdd    0.014f
C6  a      z      0.011f
C7  a      an     0.239f
C8  z      vdd    0.239f
C9  vdd    an     0.121f
C11 a      vss    0.052f
C12 z      vss    0.024f
C14 an     vss    0.087f
.ends
