magic
tech scmos
timestamp 1179387200
<< checkpaint >>
rect -22 -25 62 105
<< ab >>
rect 0 0 40 80
<< pwell >>
rect -4 -7 44 36
<< nwell >>
rect -4 36 44 87
<< polysilicon >>
rect 9 63 11 68
rect 19 63 25 64
rect 19 59 20 63
rect 24 59 25 63
rect 19 58 25 59
rect 22 55 24 58
rect 29 55 31 60
rect 9 41 11 45
rect 9 40 15 41
rect 9 36 10 40
rect 14 36 15 40
rect 22 37 24 45
rect 9 35 15 36
rect 19 35 24 37
rect 29 39 31 45
rect 29 38 35 39
rect 9 30 11 35
rect 19 30 21 35
rect 29 34 30 38
rect 34 34 35 38
rect 29 33 35 34
rect 29 30 31 33
rect 9 16 11 21
rect 19 19 21 24
rect 29 19 31 24
<< ndiffusion >>
rect 2 29 9 30
rect 2 25 3 29
rect 7 25 9 29
rect 2 24 9 25
rect 4 21 9 24
rect 11 24 19 30
rect 21 29 29 30
rect 21 25 23 29
rect 27 25 29 29
rect 21 24 29 25
rect 31 29 38 30
rect 31 25 33 29
rect 37 25 38 29
rect 31 24 38 25
rect 11 21 17 24
rect 13 17 17 21
rect 13 16 19 17
rect 13 12 14 16
rect 18 12 19 16
rect 13 11 19 12
<< pdiffusion >>
rect 13 72 19 73
rect 13 68 14 72
rect 18 68 19 72
rect 13 66 19 68
rect 13 63 17 66
rect 4 58 9 63
rect 2 57 9 58
rect 2 53 3 57
rect 7 53 9 57
rect 2 50 9 53
rect 2 46 3 50
rect 7 46 9 50
rect 2 45 9 46
rect 11 55 17 63
rect 11 45 22 55
rect 24 45 29 55
rect 31 54 38 55
rect 31 50 33 54
rect 37 50 38 54
rect 31 49 38 50
rect 31 45 36 49
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect -2 72 42 78
rect -2 68 14 72
rect 18 68 42 72
rect 2 58 6 63
rect 10 59 20 63
rect 24 59 25 63
rect 2 57 7 58
rect 2 53 3 57
rect 2 50 7 53
rect 2 46 3 50
rect 10 57 25 59
rect 10 49 14 57
rect 18 50 33 54
rect 37 50 38 54
rect 2 45 7 46
rect 2 31 6 45
rect 18 41 22 50
rect 10 40 22 41
rect 14 36 22 40
rect 34 39 38 47
rect 10 35 22 36
rect 2 29 14 31
rect 2 25 3 29
rect 7 25 14 29
rect 18 29 22 35
rect 26 38 38 39
rect 26 34 30 38
rect 34 34 38 38
rect 26 33 38 34
rect 18 25 23 29
rect 27 25 28 29
rect 32 25 33 29
rect 37 25 38 29
rect 14 16 18 17
rect 32 12 38 25
rect -2 2 42 12
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
<< ntransistor >>
rect 9 21 11 30
rect 19 24 21 30
rect 29 24 31 30
<< ptransistor >>
rect 9 45 11 63
rect 22 45 24 55
rect 29 45 31 55
<< polycontact >>
rect 20 59 24 63
rect 10 36 14 40
rect 30 34 34 38
<< ndcontact >>
rect 3 25 7 29
rect 23 25 27 29
rect 33 25 37 29
rect 14 12 18 16
<< pdcontact >>
rect 14 68 18 72
rect 3 53 7 57
rect 3 46 7 50
rect 33 50 37 54
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
<< psubstratepdiff >>
rect 0 2 40 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 40 2
rect 0 -3 40 -2
<< nsubstratendiff >>
rect 0 82 40 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 40 82
rect 0 77 40 78
<< labels >>
rlabel polycontact 12 38 12 38 6 zn
rlabel metal1 4 44 4 44 6 z
rlabel metal1 12 28 12 28 6 z
rlabel metal1 12 56 12 56 6 a
rlabel metal1 20 6 20 6 6 vss
rlabel metal1 23 27 23 27 6 zn
rlabel metal1 28 36 28 36 6 b
rlabel metal1 16 38 16 38 6 zn
rlabel metal1 20 60 20 60 6 a
rlabel metal1 20 74 20 74 6 vdd
rlabel metal1 36 40 36 40 6 b
rlabel metal1 28 52 28 52 6 zn
<< end >>
