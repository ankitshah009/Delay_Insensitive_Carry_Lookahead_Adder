magic
tech scmos
timestamp 1179385205
<< checkpaint >>
rect -22 -25 190 105
<< ab >>
rect 0 0 168 80
<< pwell >>
rect -4 -7 172 36
<< nwell >>
rect -4 36 172 87
<< polysilicon >>
rect 9 70 11 74
rect 16 70 18 74
rect 26 70 28 74
rect 33 70 35 74
rect 43 70 45 74
rect 50 70 52 74
rect 60 70 62 74
rect 67 70 69 74
rect 77 70 79 74
rect 107 70 109 74
rect 117 70 119 74
rect 127 70 129 74
rect 137 70 139 74
rect 147 70 149 74
rect 157 70 159 74
rect 87 56 89 61
rect 97 56 99 61
rect 9 29 11 42
rect 16 39 18 42
rect 26 39 28 42
rect 16 38 28 39
rect 16 34 18 38
rect 22 37 28 38
rect 22 34 23 37
rect 33 35 35 42
rect 43 35 45 42
rect 50 39 52 42
rect 60 39 62 42
rect 50 38 62 39
rect 16 33 23 34
rect 32 33 46 35
rect 50 34 51 38
rect 55 37 62 38
rect 55 34 56 37
rect 50 33 56 34
rect 32 31 34 33
rect 28 30 34 31
rect 44 30 46 33
rect 54 30 56 33
rect 67 32 69 42
rect 77 39 79 42
rect 87 39 89 42
rect 97 39 99 42
rect 107 39 109 42
rect 117 39 119 42
rect 77 38 119 39
rect 77 37 82 38
rect 81 34 82 37
rect 86 37 114 38
rect 86 34 87 37
rect 81 33 87 34
rect 113 34 114 37
rect 118 34 119 38
rect 127 39 129 42
rect 137 39 139 42
rect 147 39 149 42
rect 157 39 159 42
rect 127 38 159 39
rect 127 37 131 38
rect 113 33 119 34
rect 130 34 131 37
rect 135 37 159 38
rect 135 34 136 37
rect 130 33 136 34
rect 66 31 72 32
rect 28 29 29 30
rect 9 27 29 29
rect 28 26 29 27
rect 33 26 34 30
rect 28 25 34 26
rect 66 27 67 31
rect 71 27 72 31
rect 66 26 72 27
rect 91 31 109 33
rect 113 31 126 33
rect 91 30 97 31
rect 91 26 92 30
rect 96 26 97 30
rect 107 28 109 31
rect 114 28 116 31
rect 124 28 126 31
rect 131 28 133 33
rect 91 25 97 26
rect 44 6 46 10
rect 54 6 56 10
rect 107 6 109 11
rect 114 6 116 11
rect 124 6 126 11
rect 131 6 133 11
<< ndiffusion >>
rect 36 12 44 30
rect 36 8 37 12
rect 41 10 44 12
rect 46 22 54 30
rect 46 18 48 22
rect 52 18 54 22
rect 46 10 54 18
rect 56 12 64 30
rect 56 10 59 12
rect 41 8 42 10
rect 36 7 42 8
rect 58 8 59 10
rect 63 8 64 12
rect 58 7 64 8
rect 99 12 107 28
rect 99 8 100 12
rect 104 11 107 12
rect 109 11 114 28
rect 116 22 124 28
rect 116 18 118 22
rect 122 18 124 22
rect 116 11 124 18
rect 126 11 131 28
rect 133 23 146 28
rect 133 19 140 23
rect 144 19 146 23
rect 133 16 146 19
rect 133 12 140 16
rect 144 12 146 16
rect 133 11 146 12
rect 104 8 105 11
rect 99 7 105 8
<< pdiffusion >>
rect 4 64 9 70
rect 2 63 9 64
rect 2 59 3 63
rect 7 59 9 63
rect 2 58 9 59
rect 4 42 9 58
rect 11 42 16 70
rect 18 54 26 70
rect 18 50 20 54
rect 24 50 26 54
rect 18 42 26 50
rect 28 42 33 70
rect 35 63 43 70
rect 35 59 37 63
rect 41 59 43 63
rect 35 42 43 59
rect 45 42 50 70
rect 52 54 60 70
rect 52 50 54 54
rect 58 50 60 54
rect 52 47 60 50
rect 52 43 54 47
rect 58 43 60 47
rect 52 42 60 43
rect 62 42 67 70
rect 69 62 77 70
rect 69 58 71 62
rect 75 58 77 62
rect 69 55 77 58
rect 69 51 71 55
rect 75 51 77 55
rect 69 48 77 51
rect 69 44 71 48
rect 75 44 77 48
rect 69 42 77 44
rect 79 69 86 70
rect 79 65 81 69
rect 85 65 86 69
rect 79 64 86 65
rect 100 69 107 70
rect 100 65 101 69
rect 105 65 107 69
rect 100 64 107 65
rect 79 56 85 64
rect 101 56 107 64
rect 79 55 87 56
rect 79 51 81 55
rect 85 51 87 55
rect 79 42 87 51
rect 89 54 97 56
rect 89 50 91 54
rect 95 50 97 54
rect 89 47 97 50
rect 89 43 91 47
rect 95 43 97 47
rect 89 42 97 43
rect 99 55 107 56
rect 99 51 101 55
rect 105 51 107 55
rect 99 42 107 51
rect 109 62 117 70
rect 109 58 111 62
rect 115 58 117 62
rect 109 55 117 58
rect 109 51 111 55
rect 115 51 117 55
rect 109 48 117 51
rect 109 44 111 48
rect 115 44 117 48
rect 109 42 117 44
rect 119 69 127 70
rect 119 65 121 69
rect 125 65 127 69
rect 119 62 127 65
rect 119 58 121 62
rect 125 58 127 62
rect 119 42 127 58
rect 129 61 137 70
rect 129 57 131 61
rect 135 57 137 61
rect 129 54 137 57
rect 129 50 131 54
rect 135 50 137 54
rect 129 42 137 50
rect 139 69 147 70
rect 139 65 141 69
rect 145 65 147 69
rect 139 62 147 65
rect 139 58 141 62
rect 145 58 147 62
rect 139 42 147 58
rect 149 62 157 70
rect 149 58 151 62
rect 155 58 157 62
rect 149 55 157 58
rect 149 51 151 55
rect 155 51 157 55
rect 149 48 157 51
rect 149 44 151 48
rect 155 44 157 48
rect 149 42 157 44
rect 159 69 166 70
rect 159 65 161 69
rect 165 65 166 69
rect 159 62 166 65
rect 159 58 161 62
rect 165 58 166 62
rect 159 42 166 58
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect 118 78 122 82
rect 126 78 130 82
rect 134 78 138 82
rect 142 78 146 82
rect 150 78 154 82
rect 158 78 162 82
rect 166 78 170 82
rect -2 69 170 78
rect -2 68 81 69
rect 80 65 81 68
rect 85 68 101 69
rect 85 65 86 68
rect 2 59 3 63
rect 7 59 37 63
rect 41 62 75 63
rect 41 59 71 62
rect 71 55 75 58
rect 2 50 20 54
rect 24 50 54 54
rect 58 50 59 54
rect 2 22 6 50
rect 53 47 59 50
rect 17 38 23 46
rect 53 43 54 47
rect 58 43 59 47
rect 80 55 86 65
rect 100 65 101 68
rect 105 68 121 69
rect 105 65 106 68
rect 100 55 106 65
rect 120 65 121 68
rect 125 68 141 69
rect 125 65 126 68
rect 80 51 81 55
rect 85 51 86 55
rect 91 54 95 55
rect 71 48 75 51
rect 100 51 101 55
rect 105 51 106 55
rect 111 62 115 63
rect 120 62 126 65
rect 140 65 141 68
rect 145 68 161 69
rect 145 65 146 68
rect 140 62 146 65
rect 165 68 170 69
rect 120 58 121 62
rect 125 58 126 62
rect 131 61 135 62
rect 111 55 115 58
rect 140 58 141 62
rect 145 58 146 62
rect 151 62 155 63
rect 131 54 135 57
rect 151 55 155 58
rect 161 62 165 65
rect 161 57 165 58
rect 115 51 131 54
rect 91 47 95 50
rect 111 50 131 51
rect 135 51 151 54
rect 135 50 155 51
rect 111 48 115 50
rect 75 44 91 47
rect 71 43 91 44
rect 95 44 111 47
rect 151 48 155 50
rect 95 43 115 44
rect 130 39 134 47
rect 151 43 155 44
rect 17 34 18 38
rect 22 34 51 38
rect 55 34 56 38
rect 17 26 23 34
rect 66 31 71 39
rect 130 38 135 39
rect 66 30 67 31
rect 28 26 29 30
rect 33 27 67 30
rect 33 26 71 27
rect 81 34 82 38
rect 86 34 114 38
rect 118 34 119 38
rect 130 34 131 38
rect 81 26 87 34
rect 130 33 135 34
rect 130 30 134 33
rect 91 26 92 30
rect 96 26 134 30
rect 2 18 48 22
rect 52 18 118 22
rect 122 18 123 22
rect 130 17 134 26
rect 139 19 140 23
rect 144 19 145 23
rect 139 16 145 19
rect 139 12 140 16
rect 144 12 145 16
rect -2 8 37 12
rect 41 8 59 12
rect 63 8 100 12
rect 104 8 170 12
rect -2 2 170 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 122 2
rect 126 -2 130 2
rect 134 -2 138 2
rect 142 -2 146 2
rect 150 -2 154 2
rect 158 -2 162 2
rect 166 -2 170 2
<< ntransistor >>
rect 44 10 46 30
rect 54 10 56 30
rect 107 11 109 28
rect 114 11 116 28
rect 124 11 126 28
rect 131 11 133 28
<< ptransistor >>
rect 9 42 11 70
rect 16 42 18 70
rect 26 42 28 70
rect 33 42 35 70
rect 43 42 45 70
rect 50 42 52 70
rect 60 42 62 70
rect 67 42 69 70
rect 77 42 79 70
rect 87 42 89 56
rect 97 42 99 56
rect 107 42 109 70
rect 117 42 119 70
rect 127 42 129 70
rect 137 42 139 70
rect 147 42 149 70
rect 157 42 159 70
<< polycontact >>
rect 18 34 22 38
rect 51 34 55 38
rect 82 34 86 38
rect 114 34 118 38
rect 131 34 135 38
rect 29 26 33 30
rect 67 27 71 31
rect 92 26 96 30
<< ndcontact >>
rect 37 8 41 12
rect 48 18 52 22
rect 59 8 63 12
rect 100 8 104 12
rect 118 18 122 22
rect 140 19 144 23
rect 140 12 144 16
<< pdcontact >>
rect 3 59 7 63
rect 20 50 24 54
rect 37 59 41 63
rect 54 50 58 54
rect 54 43 58 47
rect 71 58 75 62
rect 71 51 75 55
rect 71 44 75 48
rect 81 65 85 69
rect 101 65 105 69
rect 81 51 85 55
rect 91 50 95 54
rect 91 43 95 47
rect 101 51 105 55
rect 111 58 115 62
rect 111 51 115 55
rect 111 44 115 48
rect 121 65 125 69
rect 121 58 125 62
rect 131 57 135 61
rect 131 50 135 54
rect 141 65 145 69
rect 141 58 145 62
rect 151 58 155 62
rect 151 51 155 55
rect 151 44 155 48
rect 161 65 165 69
rect 161 58 165 62
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
rect 90 -2 94 2
rect 98 -2 102 2
rect 106 -2 110 2
rect 114 -2 118 2
rect 122 -2 126 2
rect 130 -2 134 2
rect 138 -2 142 2
rect 146 -2 150 2
rect 154 -2 158 2
rect 162 -2 166 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
rect 90 78 94 82
rect 98 78 102 82
rect 106 78 110 82
rect 114 78 118 82
rect 122 78 126 82
rect 130 78 134 82
rect 138 78 142 82
rect 146 78 150 82
rect 154 78 158 82
rect 162 78 166 82
<< psubstratepdiff >>
rect 0 2 168 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 122 2
rect 126 -2 130 2
rect 134 -2 138 2
rect 142 -2 146 2
rect 150 -2 154 2
rect 158 -2 162 2
rect 166 -2 168 2
rect 0 -3 168 -2
<< nsubstratendiff >>
rect 0 82 168 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect 118 78 122 82
rect 126 78 130 82
rect 134 78 138 82
rect 142 78 146 82
rect 150 78 154 82
rect 158 78 162 82
rect 166 78 168 82
rect 0 77 168 78
<< labels >>
rlabel metal1 20 20 20 20 6 z
rlabel metal1 12 20 12 20 6 z
rlabel polycontact 20 36 20 36 6 c
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 52 12 52 6 z
rlabel metal1 20 52 20 52 6 z
rlabel metal1 28 20 28 20 6 z
rlabel metal1 52 20 52 20 6 z
rlabel metal1 44 20 44 20 6 z
rlabel metal1 36 20 36 20 6 z
rlabel metal1 36 28 36 28 6 b
rlabel metal1 44 28 44 28 6 b
rlabel metal1 52 28 52 28 6 b
rlabel metal1 28 36 28 36 6 c
rlabel polycontact 52 36 52 36 6 c
rlabel metal1 44 36 44 36 6 c
rlabel metal1 36 36 36 36 6 c
rlabel metal1 28 52 28 52 6 z
rlabel metal1 36 52 36 52 6 z
rlabel metal1 44 52 44 52 6 z
rlabel metal1 52 52 52 52 6 z
rlabel metal1 76 20 76 20 6 z
rlabel metal1 68 20 68 20 6 z
rlabel metal1 60 20 60 20 6 z
rlabel metal1 60 28 60 28 6 b
rlabel metal1 68 32 68 32 6 b
rlabel pdcontact 73 53 73 53 6 n1
rlabel pdcontact 38 61 38 61 6 n1
rlabel metal1 84 6 84 6 6 vss
rlabel metal1 84 20 84 20 6 z
rlabel metal1 108 20 108 20 6 z
rlabel metal1 100 20 100 20 6 z
rlabel metal1 92 20 92 20 6 z
rlabel metal1 100 28 100 28 6 a1
rlabel metal1 108 28 108 28 6 a1
rlabel metal1 84 32 84 32 6 a2
rlabel metal1 108 36 108 36 6 a2
rlabel metal1 100 36 100 36 6 a2
rlabel metal1 92 36 92 36 6 a2
rlabel metal1 93 49 93 49 6 n1
rlabel metal1 84 74 84 74 6 vdd
rlabel metal1 116 20 116 20 6 z
rlabel metal1 124 28 124 28 6 a1
rlabel metal1 116 28 116 28 6 a1
rlabel polycontact 116 36 116 36 6 a2
rlabel metal1 132 32 132 32 6 a1
rlabel metal1 133 56 133 56 6 n1
rlabel pdcontact 133 52 133 52 6 n1
<< end >>
