magic
tech scmos
timestamp 1179386987
<< checkpaint >>
rect -22 -25 86 105
<< ab >>
rect 0 0 64 80
<< pwell >>
rect -4 -7 68 36
<< nwell >>
rect -4 36 68 87
<< polysilicon >>
rect 19 66 21 71
rect 26 66 28 71
rect 9 58 11 63
rect 40 62 42 67
rect 9 38 11 50
rect 9 37 15 38
rect 9 33 10 37
rect 14 33 15 37
rect 9 32 15 33
rect 19 32 21 50
rect 26 47 28 50
rect 40 47 42 50
rect 26 46 33 47
rect 26 42 27 46
rect 31 42 33 46
rect 40 46 55 47
rect 40 45 50 46
rect 26 41 33 42
rect 49 42 50 45
rect 54 42 55 46
rect 49 41 55 42
rect 9 23 11 32
rect 19 31 25 32
rect 19 27 20 31
rect 24 27 25 31
rect 19 26 25 27
rect 19 23 21 26
rect 31 23 33 41
rect 51 30 53 41
rect 51 19 53 24
rect 9 11 11 16
rect 19 11 21 16
rect 31 11 33 16
<< ndiffusion >>
rect 44 29 51 30
rect 44 25 45 29
rect 49 25 51 29
rect 44 24 51 25
rect 53 29 60 30
rect 53 25 55 29
rect 59 25 60 29
rect 53 24 60 25
rect 2 22 9 23
rect 2 18 3 22
rect 7 18 9 22
rect 2 16 9 18
rect 11 21 19 23
rect 11 17 13 21
rect 17 17 19 21
rect 11 16 19 17
rect 21 16 31 23
rect 33 21 40 23
rect 33 17 35 21
rect 39 17 40 21
rect 33 16 40 17
rect 23 12 29 16
rect 23 8 24 12
rect 28 8 29 12
rect 23 7 29 8
<< pdiffusion >>
rect 14 58 19 66
rect 2 57 9 58
rect 2 53 3 57
rect 7 53 9 57
rect 2 50 9 53
rect 11 55 19 58
rect 11 51 13 55
rect 17 51 19 55
rect 11 50 19 51
rect 21 50 26 66
rect 28 62 37 66
rect 28 61 40 62
rect 28 57 34 61
rect 38 57 40 61
rect 28 50 40 57
rect 42 56 47 62
rect 42 55 49 56
rect 42 51 44 55
rect 48 51 49 55
rect 42 50 49 51
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect -2 68 66 78
rect 3 57 7 68
rect 34 61 38 68
rect 34 56 38 57
rect 3 52 7 53
rect 10 51 13 55
rect 17 51 22 55
rect 10 49 22 51
rect 10 47 14 49
rect 2 43 14 47
rect 26 46 30 55
rect 42 51 44 55
rect 48 51 49 55
rect 2 23 6 43
rect 26 42 27 46
rect 31 42 39 46
rect 10 37 23 38
rect 14 34 23 37
rect 10 25 14 33
rect 42 31 46 51
rect 50 46 62 47
rect 54 42 62 46
rect 50 41 62 42
rect 58 33 62 41
rect 19 27 20 31
rect 24 29 46 31
rect 24 27 45 29
rect 42 25 45 27
rect 49 25 50 29
rect 54 25 55 29
rect 59 25 60 29
rect 2 22 7 23
rect 2 18 3 22
rect 2 17 7 18
rect 12 17 13 21
rect 17 17 35 21
rect 39 17 40 21
rect 54 12 60 25
rect -2 8 24 12
rect 28 8 66 12
rect -2 2 66 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
<< ntransistor >>
rect 51 24 53 30
rect 9 16 11 23
rect 19 16 21 23
rect 31 16 33 23
<< ptransistor >>
rect 9 50 11 58
rect 19 50 21 66
rect 26 50 28 66
rect 40 50 42 62
<< polycontact >>
rect 10 33 14 37
rect 27 42 31 46
rect 50 42 54 46
rect 20 27 24 31
<< ndcontact >>
rect 45 25 49 29
rect 55 25 59 29
rect 3 18 7 22
rect 13 17 17 21
rect 35 17 39 21
rect 24 8 28 12
<< pdcontact >>
rect 3 53 7 57
rect 13 51 17 55
rect 34 57 38 61
rect 44 51 48 55
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
<< psubstratepdiff >>
rect 0 2 64 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 64 2
rect 0 -3 64 -2
<< nsubstratendiff >>
rect 0 82 64 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 64 82
rect 0 77 64 78
<< labels >>
rlabel polycontact 22 29 22 29 6 a2n
rlabel metal1 4 32 4 32 6 z
rlabel metal1 12 28 12 28 6 b
rlabel metal1 20 36 20 36 6 b
rlabel metal1 20 52 20 52 6 z
rlabel metal1 12 52 12 52 6 z
rlabel metal1 32 6 32 6 6 vss
rlabel metal1 36 44 36 44 6 a1
rlabel metal1 28 52 28 52 6 a1
rlabel metal1 32 74 32 74 6 vdd
rlabel metal1 26 19 26 19 6 n1
rlabel ndcontact 46 27 46 27 6 a2n
rlabel metal1 32 29 32 29 6 a2n
rlabel pdcontact 45 53 45 53 6 a2n
rlabel polycontact 52 44 52 44 6 a2
rlabel metal1 60 40 60 40 6 a2
<< end >>
