magic
tech scmos
timestamp 1180600717
<< checkpaint >>
rect -22 -22 72 122
<< ab >>
rect 0 0 50 100
<< pwell >>
rect -4 -4 54 48
<< nwell >>
rect -4 48 54 104
<< polysilicon >>
rect 19 94 21 98
rect 27 94 29 98
rect 35 94 37 98
rect 19 53 21 56
rect 17 52 23 53
rect 17 49 18 52
rect 11 48 18 49
rect 22 48 23 52
rect 11 47 23 48
rect 11 25 13 47
rect 27 43 29 56
rect 35 53 37 56
rect 35 51 39 53
rect 27 42 33 43
rect 27 39 28 42
rect 23 38 28 39
rect 32 38 33 42
rect 23 37 33 38
rect 23 25 25 37
rect 37 33 39 51
rect 37 32 43 33
rect 37 29 38 32
rect 35 28 38 29
rect 42 28 43 32
rect 35 27 43 28
rect 35 24 37 27
rect 11 11 13 15
rect 23 11 25 15
rect 35 10 37 14
<< ndiffusion >>
rect 3 22 11 25
rect 3 18 4 22
rect 8 18 11 22
rect 3 15 11 18
rect 13 15 23 25
rect 25 24 30 25
rect 25 22 35 24
rect 25 18 28 22
rect 32 18 35 22
rect 25 15 35 18
rect 15 12 21 15
rect 15 8 16 12
rect 20 8 21 12
rect 27 14 35 15
rect 37 14 45 24
rect 39 12 45 14
rect 15 7 21 8
rect 39 8 40 12
rect 44 8 45 12
rect 39 7 45 8
<< pdiffusion >>
rect 14 85 19 94
rect 7 82 19 85
rect 7 78 8 82
rect 12 78 19 82
rect 7 72 19 78
rect 7 68 8 72
rect 12 68 19 72
rect 7 62 19 68
rect 7 58 8 62
rect 12 58 19 62
rect 7 56 19 58
rect 21 56 27 94
rect 29 56 35 94
rect 37 92 45 94
rect 37 88 40 92
rect 44 88 45 92
rect 37 56 45 88
rect 7 55 13 56
<< metal1 >>
rect -2 92 52 100
rect -2 88 40 92
rect 44 88 52 92
rect 8 82 12 83
rect 8 72 12 78
rect 8 62 12 68
rect 8 22 12 58
rect 18 52 22 83
rect 18 27 22 48
rect 28 42 32 83
rect 28 27 32 38
rect 38 32 42 83
rect 3 18 4 22
rect 8 18 28 22
rect 32 18 33 22
rect 38 17 42 28
rect -2 8 16 12
rect 20 8 40 12
rect 44 8 52 12
rect -2 0 52 8
<< ntransistor >>
rect 11 15 13 25
rect 23 15 25 25
rect 35 14 37 24
<< ptransistor >>
rect 19 56 21 94
rect 27 56 29 94
rect 35 56 37 94
<< polycontact >>
rect 18 48 22 52
rect 28 38 32 42
rect 38 28 42 32
<< ndcontact >>
rect 4 18 8 22
rect 28 18 32 22
rect 16 8 20 12
rect 40 8 44 12
<< pdcontact >>
rect 8 78 12 82
rect 8 68 12 72
rect 8 58 12 62
rect 40 88 44 92
<< labels >>
rlabel metal1 20 20 20 20 6 nq
rlabel metal1 10 50 10 50 6 nq
rlabel metal1 20 55 20 55 6 i1
rlabel metal1 25 6 25 6 6 vss
rlabel ndcontact 30 20 30 20 6 nq
rlabel metal1 30 55 30 55 6 i0
rlabel metal1 25 94 25 94 6 vdd
rlabel metal1 40 50 40 50 6 i2
<< end >>
