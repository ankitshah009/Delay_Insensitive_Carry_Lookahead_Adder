magic
tech scmos
timestamp 1180600734
<< checkpaint >>
rect -22 -22 132 122
<< ab >>
rect 0 0 110 100
<< pwell >>
rect -4 -4 114 48
<< nwell >>
rect -4 48 114 104
<< polysilicon >>
rect 11 85 13 89
rect 23 85 25 89
rect 35 85 37 89
rect 83 94 85 98
rect 95 94 97 98
rect 47 85 49 89
rect 71 76 73 80
rect 11 43 13 65
rect 23 43 25 65
rect 7 42 13 43
rect 7 38 8 42
rect 12 38 13 42
rect 7 37 13 38
rect 17 42 25 43
rect 17 38 18 42
rect 22 38 25 42
rect 17 37 25 38
rect 11 25 13 37
rect 23 25 25 37
rect 35 43 37 65
rect 47 43 49 65
rect 71 53 73 56
rect 71 52 79 53
rect 71 48 74 52
rect 78 48 79 52
rect 71 47 79 48
rect 35 42 43 43
rect 35 38 38 42
rect 42 38 43 42
rect 35 37 43 38
rect 47 42 53 43
rect 47 38 48 42
rect 52 38 53 42
rect 47 37 53 38
rect 35 25 37 37
rect 47 25 49 37
rect 71 25 73 47
rect 83 43 85 55
rect 95 43 97 55
rect 77 42 97 43
rect 77 38 78 42
rect 82 38 97 42
rect 77 37 97 38
rect 83 25 85 37
rect 95 25 97 37
rect 11 11 13 15
rect 23 11 25 15
rect 35 11 37 15
rect 47 11 49 15
rect 71 11 73 15
rect 83 2 85 6
rect 95 2 97 6
<< ndiffusion >>
rect 3 15 11 25
rect 13 15 23 25
rect 25 22 35 25
rect 25 18 28 22
rect 32 18 35 22
rect 25 15 35 18
rect 37 15 47 25
rect 49 15 57 25
rect 63 22 71 25
rect 63 18 64 22
rect 68 18 71 22
rect 63 15 71 18
rect 73 22 83 25
rect 73 18 76 22
rect 80 18 83 22
rect 73 15 83 18
rect 3 12 9 15
rect 3 8 4 12
rect 8 8 9 12
rect 51 12 57 15
rect 3 7 9 8
rect 51 8 52 12
rect 56 8 57 12
rect 75 12 83 15
rect 51 7 57 8
rect 75 8 76 12
rect 80 8 83 12
rect 75 6 83 8
rect 85 22 95 25
rect 85 18 88 22
rect 92 18 95 22
rect 85 6 95 18
rect 97 22 105 25
rect 97 18 100 22
rect 104 18 105 22
rect 97 12 105 18
rect 97 8 100 12
rect 104 8 105 12
rect 97 6 105 8
<< pdiffusion >>
rect 39 92 45 93
rect 39 88 40 92
rect 44 88 45 92
rect 75 92 83 94
rect 39 85 45 88
rect 75 88 76 92
rect 80 88 83 92
rect 3 82 11 85
rect 3 78 4 82
rect 8 78 11 82
rect 3 65 11 78
rect 13 72 23 85
rect 13 68 16 72
rect 20 68 23 72
rect 13 65 23 68
rect 25 82 35 85
rect 25 78 28 82
rect 32 78 35 82
rect 25 65 35 78
rect 37 65 47 85
rect 49 82 57 85
rect 49 78 52 82
rect 56 78 57 82
rect 75 82 83 88
rect 49 65 57 78
rect 75 78 76 82
rect 80 78 83 82
rect 75 76 83 78
rect 63 62 71 76
rect 63 58 64 62
rect 68 58 71 62
rect 63 56 71 58
rect 73 56 83 76
rect 78 55 83 56
rect 85 82 95 94
rect 85 78 88 82
rect 92 78 95 82
rect 85 72 95 78
rect 85 68 88 72
rect 92 68 95 72
rect 85 62 95 68
rect 85 58 88 62
rect 92 58 95 62
rect 85 55 95 58
rect 97 92 105 94
rect 97 88 100 92
rect 104 88 105 92
rect 97 82 105 88
rect 97 78 100 82
rect 104 78 105 82
rect 97 72 105 78
rect 97 68 100 72
rect 104 68 105 72
rect 97 62 105 68
rect 97 58 100 62
rect 104 58 105 62
rect 97 55 105 58
<< metal1 >>
rect -2 96 112 100
rect -2 92 4 96
rect 8 92 16 96
rect 20 92 28 96
rect 32 92 52 96
rect 56 92 64 96
rect 68 92 112 96
rect -2 88 40 92
rect 44 88 76 92
rect 80 88 100 92
rect 104 88 112 92
rect 76 82 80 88
rect 3 78 4 82
rect 8 78 28 82
rect 32 78 52 82
rect 56 78 57 82
rect 76 77 80 78
rect 88 82 92 83
rect 88 72 92 78
rect 15 68 16 72
rect 20 68 78 72
rect 8 42 12 63
rect 8 17 12 38
rect 18 42 22 63
rect 18 17 22 38
rect 28 22 32 68
rect 28 17 32 18
rect 38 42 42 63
rect 38 17 42 38
rect 48 42 52 63
rect 48 17 52 38
rect 64 62 68 63
rect 64 42 68 58
rect 74 52 78 68
rect 74 47 78 48
rect 88 62 92 68
rect 64 38 78 42
rect 82 38 83 42
rect 64 22 68 38
rect 64 17 68 18
rect 76 22 80 23
rect 76 12 80 18
rect 88 22 92 58
rect 100 82 104 88
rect 100 72 104 78
rect 100 62 104 68
rect 100 57 104 58
rect 88 17 92 18
rect 100 22 104 23
rect 100 12 104 18
rect -2 8 4 12
rect 8 8 52 12
rect 56 8 76 12
rect 80 8 100 12
rect 104 8 112 12
rect -2 4 16 8
rect 20 4 28 8
rect 32 4 40 8
rect 44 4 112 8
rect -2 0 112 4
<< ntransistor >>
rect 11 15 13 25
rect 23 15 25 25
rect 35 15 37 25
rect 47 15 49 25
rect 71 15 73 25
rect 83 6 85 25
rect 95 6 97 25
<< ptransistor >>
rect 11 65 13 85
rect 23 65 25 85
rect 35 65 37 85
rect 47 65 49 85
rect 71 56 73 76
rect 83 55 85 94
rect 95 55 97 94
<< polycontact >>
rect 8 38 12 42
rect 18 38 22 42
rect 74 48 78 52
rect 38 38 42 42
rect 48 38 52 42
rect 78 38 82 42
<< ndcontact >>
rect 28 18 32 22
rect 64 18 68 22
rect 76 18 80 22
rect 4 8 8 12
rect 52 8 56 12
rect 76 8 80 12
rect 88 18 92 22
rect 100 18 104 22
rect 100 8 104 12
<< pdcontact >>
rect 40 88 44 92
rect 76 88 80 92
rect 4 78 8 82
rect 16 68 20 72
rect 28 78 32 82
rect 52 78 56 82
rect 76 78 80 82
rect 64 58 68 62
rect 88 78 92 82
rect 88 68 92 72
rect 88 58 92 62
rect 100 88 104 92
rect 100 78 104 82
rect 100 68 104 72
rect 100 58 104 62
<< psubstratepcontact >>
rect 16 4 20 8
rect 28 4 32 8
rect 40 4 44 8
<< nsubstratencontact >>
rect 4 92 8 96
rect 16 92 20 96
rect 28 92 32 96
rect 52 92 56 96
rect 64 92 68 96
<< psubstratepdiff >>
rect 15 8 45 9
rect 15 4 16 8
rect 20 4 28 8
rect 32 4 40 8
rect 44 4 45 8
rect 15 3 45 4
<< nsubstratendiff >>
rect 3 96 33 97
rect 3 92 4 96
rect 8 92 16 96
rect 20 92 28 96
rect 32 92 33 96
rect 51 96 69 97
rect 3 91 33 92
rect 51 92 52 96
rect 56 92 64 96
rect 68 92 69 96
rect 51 91 69 92
<< labels >>
rlabel polycontact 10 40 10 40 6 i0
rlabel polycontact 40 40 40 40 6 i3
rlabel polycontact 20 40 20 40 6 i1
rlabel metal1 55 6 55 6 6 vss
rlabel polycontact 50 40 50 40 6 i2
rlabel nsubstratencontact 55 94 55 94 6 vdd
rlabel metal1 90 50 90 50 6 nq
<< end >>
