.subckt oai21bv0x05 a1 a2 b vdd vss z
*   SPICE3 file   created from oai21bv0x05.ext -      technology: scmos
m00 z      bn     vdd    vdd p w=8u   l=2.3636u ad=34.6667p pd=16u      as=59.5294p ps=23.0588u
m01 w1     a2     z      vdd p w=16u  l=2.3636u ad=40p      pd=21u      as=69.3333p ps=32u
m02 vdd    a1     w1     vdd p w=16u  l=2.3636u ad=119.059p pd=46.1176u as=40p      ps=21u
m03 bn     b      vdd    vdd p w=10u  l=2.3636u ad=62p      pd=34u      as=74.4118p ps=28.8235u
m04 n1     bn     z      vss n w=7u   l=2.3636u ad=35p      pd=19.3333u as=49p      ps=28u
m05 vss    a2     n1     vss n w=7u   l=2.3636u ad=72.8p    pd=32.2u    as=35p      ps=19.3333u
m06 vss    b      bn     vss n w=6u   l=2.3636u ad=62.4p    pd=27.6u    as=42p      ps=26u
m07 n1     a1     vss    vss n w=7u   l=2.3636u ad=35p      pd=19.3333u as=72.8p    ps=32.2u
C0  vss    vdd    0.003f
C1  b      a2     0.017f
C2  n1     bn     0.035f
C3  b      vdd    0.021f
C4  z      a2     0.033f
C5  w1     bn     0.007f
C6  vss    n1     0.194f
C7  a1     bn     0.265f
C8  z      vdd    0.160f
C9  a2     vdd    0.025f
C10 vss    a1     0.030f
C11 n1     z      0.065f
C12 b      a1     0.039f
C13 n1     a2     0.076f
C14 vss    bn     0.075f
C15 n1     vdd    0.008f
C16 z      a1     0.131f
C17 b      bn     0.096f
C18 z      bn     0.181f
C19 a1     a2     0.232f
C20 vss    b      0.019f
C21 a2     bn     0.209f
C22 a1     vdd    0.041f
C23 vss    z      0.027f
C24 bn     vdd    0.139f
C25 n1     a1     0.046f
C26 vss    a2     0.039f
C28 n1     vss    0.005f
C29 b      vss    0.031f
C30 z      vss    0.017f
C31 a1     vss    0.032f
C32 a2     vss    0.027f
C33 bn     vss    0.032f
.ends
