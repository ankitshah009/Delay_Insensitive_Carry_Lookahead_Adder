magic
tech scmos
timestamp 1179387083
<< checkpaint >>
rect -22 -25 78 105
<< ab >>
rect 0 0 56 80
<< pwell >>
rect -4 -7 60 36
<< nwell >>
rect -4 36 60 87
<< polysilicon >>
rect 13 70 15 74
rect 21 70 23 74
rect 31 70 33 74
rect 39 70 41 74
rect 13 40 15 43
rect 21 40 23 43
rect 9 39 15 40
rect 9 35 10 39
rect 14 35 15 39
rect 9 34 15 35
rect 19 39 25 40
rect 31 39 33 43
rect 39 40 41 43
rect 39 39 48 40
rect 19 35 20 39
rect 24 35 25 39
rect 19 34 25 35
rect 29 38 35 39
rect 29 34 30 38
rect 34 34 35 38
rect 39 35 43 39
rect 47 35 48 39
rect 39 34 48 35
rect 9 30 11 34
rect 19 30 21 34
rect 29 33 35 34
rect 29 27 31 33
rect 41 27 43 34
rect 9 11 11 16
rect 19 11 21 16
rect 29 11 31 16
rect 41 11 43 16
<< ndiffusion >>
rect 4 22 9 30
rect 2 21 9 22
rect 2 17 3 21
rect 7 17 9 21
rect 2 16 9 17
rect 11 29 19 30
rect 11 25 13 29
rect 17 25 19 29
rect 11 16 19 25
rect 21 27 26 30
rect 21 21 29 27
rect 21 17 23 21
rect 27 17 29 21
rect 21 16 29 17
rect 31 16 41 27
rect 43 22 48 27
rect 43 21 50 22
rect 43 17 45 21
rect 49 17 50 21
rect 43 16 50 17
rect 33 12 39 16
rect 33 8 34 12
rect 38 8 39 12
rect 33 7 39 8
<< pdiffusion >>
rect 5 69 13 70
rect 5 65 7 69
rect 11 65 13 69
rect 5 43 13 65
rect 15 43 21 70
rect 23 62 31 70
rect 23 58 25 62
rect 29 58 31 62
rect 23 43 31 58
rect 33 43 39 70
rect 41 69 48 70
rect 41 65 43 69
rect 47 65 48 69
rect 41 62 48 65
rect 41 58 43 62
rect 47 58 48 62
rect 41 43 48 58
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect -2 69 58 78
rect -2 68 7 69
rect 6 65 7 68
rect 11 68 43 69
rect 11 65 12 68
rect 42 65 43 68
rect 47 68 58 69
rect 47 65 48 68
rect 2 58 25 62
rect 29 58 30 62
rect 2 29 6 58
rect 34 54 38 63
rect 42 62 48 65
rect 42 58 43 62
rect 47 58 48 62
rect 10 50 23 54
rect 34 50 47 54
rect 10 39 14 50
rect 10 33 14 35
rect 18 42 39 46
rect 18 39 24 42
rect 18 35 20 39
rect 43 39 47 50
rect 18 33 24 35
rect 29 34 30 38
rect 34 34 39 38
rect 43 34 47 35
rect 33 30 39 34
rect 2 25 13 29
rect 17 25 18 29
rect 33 26 47 30
rect 2 17 3 21
rect 7 17 23 21
rect 27 17 45 21
rect 49 17 50 21
rect -2 8 34 12
rect 38 8 58 12
rect -2 2 58 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
<< ntransistor >>
rect 9 16 11 30
rect 19 16 21 30
rect 29 16 31 27
rect 41 16 43 27
<< ptransistor >>
rect 13 43 15 70
rect 21 43 23 70
rect 31 43 33 70
rect 39 43 41 70
<< polycontact >>
rect 10 35 14 39
rect 20 35 24 39
rect 30 34 34 38
rect 43 35 47 39
<< ndcontact >>
rect 3 17 7 21
rect 13 25 17 29
rect 23 17 27 21
rect 45 17 49 21
rect 34 8 38 12
<< pdcontact >>
rect 7 65 11 69
rect 25 58 29 62
rect 43 65 47 69
rect 43 58 47 62
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
<< psubstratepdiff >>
rect 0 2 56 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 56 2
rect 0 -3 56 -2
<< nsubstratendiff >>
rect 0 82 56 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 56 82
rect 0 77 56 78
<< labels >>
rlabel metal1 4 40 4 40 6 z
rlabel metal1 12 40 12 40 6 b1
rlabel metal1 12 60 12 60 6 z
rlabel metal1 28 6 28 6 6 vss
rlabel metal1 20 36 20 36 6 b2
rlabel metal1 28 44 28 44 6 b2
rlabel metal1 20 52 20 52 6 b1
rlabel metal1 20 60 20 60 6 z
rlabel metal1 28 74 28 74 6 vdd
rlabel metal1 44 28 44 28 6 a2
rlabel metal1 36 32 36 32 6 a2
rlabel metal1 36 44 36 44 6 b2
rlabel metal1 44 52 44 52 6 a1
rlabel metal1 36 60 36 60 6 a1
rlabel ndcontact 26 19 26 19 6 n3
<< end >>
