.subckt inv_x2 i nq vdd vss
*   SPICE3 file   created from inv_x2.ext -      technology: scmos
m00 nq     i      vdd    vdd p w=30u  l=2.3636u ad=240p     pd=76u      as=364p     ps=96u
m01 nq     i      vss    vss n w=20u  l=2.3636u ad=160p     pd=56u      as=264p     ps=76u
C0  vss    i      0.074f
C1  nq     vdd    0.046f
C2  vss    nq     0.046f
C3  nq     i      0.485f
C4  i      vdd    0.093f
C6  nq     vss    0.015f
C7  i      vss    0.029f
.ends
