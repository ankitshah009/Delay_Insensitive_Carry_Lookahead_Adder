magic
tech scmos
timestamp 1185039149
<< checkpaint >>
rect -22 -24 202 124
<< ab >>
rect 0 0 180 100
<< pwell >>
rect -2 -4 182 49
<< nwell >>
rect -2 49 182 104
<< polysilicon >>
rect 47 95 49 98
rect 59 95 61 98
rect 95 95 97 98
rect 107 95 109 98
rect 119 95 121 98
rect 131 95 133 98
rect 143 95 145 98
rect 155 95 157 98
rect 167 95 169 98
rect 11 85 13 88
rect 23 85 25 88
rect 71 85 73 88
rect 83 85 85 88
rect 47 73 49 75
rect 47 72 53 73
rect 47 68 48 72
rect 52 68 53 72
rect 47 67 53 68
rect 11 63 13 65
rect 11 62 19 63
rect 11 58 14 62
rect 18 58 19 62
rect 11 57 19 58
rect 3 52 9 53
rect 3 48 4 52
rect 8 51 9 52
rect 23 51 25 65
rect 59 63 61 75
rect 95 73 97 75
rect 95 72 103 73
rect 95 68 98 72
rect 102 68 103 72
rect 95 67 103 68
rect 71 63 73 65
rect 37 62 43 63
rect 37 58 38 62
rect 42 61 43 62
rect 57 62 63 63
rect 57 61 58 62
rect 42 59 58 61
rect 42 58 43 59
rect 37 57 43 58
rect 57 58 58 59
rect 62 58 63 62
rect 57 57 63 58
rect 67 62 73 63
rect 67 58 68 62
rect 72 58 73 62
rect 67 57 73 58
rect 67 52 73 53
rect 67 51 68 52
rect 8 49 68 51
rect 8 48 9 49
rect 3 47 9 48
rect 11 32 19 33
rect 11 28 14 32
rect 18 28 19 32
rect 11 27 19 28
rect 11 25 13 27
rect 23 25 25 49
rect 67 48 68 49
rect 72 51 73 52
rect 83 51 85 65
rect 107 63 109 75
rect 101 62 109 63
rect 101 58 102 62
rect 106 58 109 62
rect 101 57 109 58
rect 119 51 121 75
rect 131 73 133 75
rect 125 72 133 73
rect 125 68 126 72
rect 130 68 133 72
rect 125 67 133 68
rect 143 53 145 75
rect 143 52 151 53
rect 72 49 133 51
rect 72 48 73 49
rect 67 47 73 48
rect 29 42 35 43
rect 29 38 30 42
rect 34 41 35 42
rect 77 42 85 43
rect 77 41 78 42
rect 34 39 78 41
rect 34 38 35 39
rect 29 37 35 38
rect 77 38 78 39
rect 82 41 85 42
rect 119 42 127 43
rect 119 41 122 42
rect 82 39 122 41
rect 82 38 85 39
rect 77 37 85 38
rect 47 32 53 33
rect 47 28 48 32
rect 52 28 53 32
rect 47 27 53 28
rect 57 32 63 33
rect 57 28 58 32
rect 62 28 63 32
rect 57 27 63 28
rect 67 32 73 33
rect 67 28 68 32
rect 72 28 73 32
rect 67 27 73 28
rect 47 25 49 27
rect 59 25 61 27
rect 71 25 73 27
rect 83 25 85 37
rect 119 38 122 39
rect 126 38 127 42
rect 119 37 127 38
rect 101 32 109 33
rect 101 28 102 32
rect 106 28 109 32
rect 101 27 109 28
rect 95 22 103 23
rect 95 18 98 22
rect 102 18 103 22
rect 95 17 103 18
rect 95 15 97 17
rect 107 15 109 27
rect 119 25 121 37
rect 131 25 133 49
rect 143 48 146 52
rect 150 48 151 52
rect 143 47 151 48
rect 155 43 157 55
rect 167 43 169 55
rect 145 42 169 43
rect 145 38 146 42
rect 150 38 169 42
rect 145 37 169 38
rect 143 32 151 33
rect 143 28 146 32
rect 150 28 151 32
rect 143 27 151 28
rect 143 25 145 27
rect 155 25 157 37
rect 167 25 169 37
rect 11 12 13 15
rect 23 12 25 15
rect 47 12 49 15
rect 59 12 61 15
rect 71 12 73 15
rect 83 12 85 15
rect 119 12 121 15
rect 131 12 133 15
rect 143 12 145 15
rect 95 2 97 5
rect 107 2 109 5
rect 155 2 157 5
rect 167 2 169 5
<< ndiffusion >>
rect 3 22 11 25
rect 3 18 4 22
rect 8 18 11 22
rect 3 15 11 18
rect 13 15 23 25
rect 25 22 33 25
rect 25 18 28 22
rect 32 18 33 22
rect 25 15 33 18
rect 39 22 47 25
rect 39 18 40 22
rect 44 18 47 22
rect 39 15 47 18
rect 49 15 59 25
rect 61 15 71 25
rect 73 22 83 25
rect 73 18 76 22
rect 80 18 83 22
rect 73 15 83 18
rect 85 15 93 25
rect 111 22 119 25
rect 111 18 112 22
rect 116 18 119 22
rect 111 15 119 18
rect 121 22 131 25
rect 121 18 124 22
rect 128 18 131 22
rect 121 15 131 18
rect 133 15 143 25
rect 145 22 155 25
rect 145 18 148 22
rect 152 18 155 22
rect 145 15 155 18
rect 15 12 21 15
rect 51 12 57 15
rect 15 8 16 12
rect 20 8 21 12
rect 15 7 21 8
rect 51 8 52 12
rect 56 8 57 12
rect 51 7 57 8
rect 87 5 95 15
rect 97 12 107 15
rect 97 8 100 12
rect 104 8 107 12
rect 97 5 107 8
rect 109 5 117 15
rect 147 12 155 15
rect 147 8 148 12
rect 152 8 155 12
rect 147 5 155 8
rect 157 22 167 25
rect 157 18 160 22
rect 164 18 167 22
rect 157 5 167 18
rect 169 22 177 25
rect 169 18 172 22
rect 176 18 177 22
rect 169 12 177 18
rect 169 8 172 12
rect 176 8 177 12
rect 169 5 177 8
<< pdiffusion >>
rect 15 92 21 93
rect 15 88 16 92
rect 20 88 21 92
rect 15 85 21 88
rect 3 82 11 85
rect 3 78 4 82
rect 8 78 11 82
rect 3 72 11 78
rect 3 68 4 72
rect 8 68 11 72
rect 3 65 11 68
rect 13 65 23 85
rect 25 72 33 85
rect 39 82 47 95
rect 39 78 40 82
rect 44 78 47 82
rect 39 75 47 78
rect 49 92 59 95
rect 49 88 52 92
rect 56 88 59 92
rect 49 75 59 88
rect 61 85 69 95
rect 87 85 95 95
rect 61 75 71 85
rect 25 68 28 72
rect 32 68 33 72
rect 25 65 33 68
rect 63 65 71 75
rect 73 72 83 85
rect 73 68 76 72
rect 80 68 83 72
rect 73 65 83 68
rect 85 75 95 85
rect 97 92 107 95
rect 97 88 100 92
rect 104 88 107 92
rect 97 75 107 88
rect 109 82 119 95
rect 109 78 112 82
rect 116 78 119 82
rect 109 75 119 78
rect 121 82 131 95
rect 121 78 124 82
rect 128 78 131 82
rect 121 75 131 78
rect 133 75 143 95
rect 145 92 155 95
rect 145 88 148 92
rect 152 88 155 92
rect 145 82 155 88
rect 145 78 148 82
rect 152 78 155 82
rect 145 75 155 78
rect 85 65 93 75
rect 147 72 155 75
rect 147 68 148 72
rect 152 68 155 72
rect 147 62 155 68
rect 147 58 148 62
rect 152 58 155 62
rect 147 55 155 58
rect 157 82 167 95
rect 157 78 160 82
rect 164 78 167 82
rect 157 72 167 78
rect 157 68 160 72
rect 164 68 167 72
rect 157 62 167 68
rect 157 58 160 62
rect 164 58 167 62
rect 157 55 167 58
rect 169 92 177 95
rect 169 88 172 92
rect 176 88 177 92
rect 169 82 177 88
rect 169 78 172 82
rect 176 78 177 82
rect 169 72 177 78
rect 169 68 172 72
rect 176 68 177 72
rect 169 62 177 68
rect 169 58 172 62
rect 176 58 177 62
rect 169 55 177 58
<< metal1 >>
rect -2 92 182 101
rect -2 88 16 92
rect 20 88 52 92
rect 56 88 100 92
rect 104 88 148 92
rect 152 88 172 92
rect 176 88 182 92
rect -2 87 182 88
rect 3 82 9 83
rect 39 82 45 83
rect 58 82 62 83
rect 3 78 4 82
rect 8 78 9 82
rect 3 77 9 78
rect 4 73 8 77
rect 3 72 9 73
rect 3 68 4 72
rect 8 68 9 72
rect 3 67 9 68
rect 4 53 8 67
rect 17 63 23 82
rect 39 78 40 82
rect 44 78 45 82
rect 39 77 45 78
rect 49 78 62 82
rect 27 72 33 73
rect 27 68 28 72
rect 32 68 33 72
rect 27 67 33 68
rect 13 62 23 63
rect 13 58 14 62
rect 18 58 23 62
rect 13 57 23 58
rect 3 52 9 53
rect 3 48 4 52
rect 8 48 9 52
rect 3 47 9 48
rect 4 23 8 47
rect 17 33 23 57
rect 13 32 23 33
rect 13 28 14 32
rect 18 28 23 32
rect 13 27 23 28
rect 3 22 9 23
rect 3 18 4 22
rect 8 18 9 22
rect 17 18 23 27
rect 28 43 32 67
rect 39 63 43 77
rect 49 73 53 78
rect 58 77 62 78
rect 111 82 117 83
rect 111 78 112 82
rect 116 78 117 82
rect 111 77 117 78
rect 123 82 129 83
rect 147 82 153 87
rect 159 82 165 83
rect 123 78 124 82
rect 128 78 140 82
rect 123 77 129 78
rect 37 62 43 63
rect 37 58 38 62
rect 42 58 43 62
rect 37 57 43 58
rect 28 42 35 43
rect 28 38 30 42
rect 34 38 35 42
rect 28 37 35 38
rect 28 23 32 37
rect 39 23 43 57
rect 47 72 53 73
rect 47 68 48 72
rect 52 68 53 72
rect 47 32 53 68
rect 75 72 81 73
rect 97 72 103 73
rect 112 72 116 77
rect 125 72 131 73
rect 75 68 76 72
rect 80 68 92 72
rect 75 67 81 68
rect 57 62 63 63
rect 57 58 58 62
rect 62 58 63 62
rect 57 57 63 58
rect 67 62 73 63
rect 88 62 92 68
rect 97 68 98 72
rect 102 68 116 72
rect 97 67 103 68
rect 101 62 107 63
rect 67 58 68 62
rect 72 58 82 62
rect 67 57 73 58
rect 58 33 62 57
rect 67 52 73 53
rect 67 48 68 52
rect 72 48 73 52
rect 67 47 73 48
rect 68 33 72 47
rect 78 43 82 58
rect 88 58 102 62
rect 106 58 107 62
rect 77 42 83 43
rect 77 38 78 42
rect 82 38 83 42
rect 77 37 83 38
rect 47 28 48 32
rect 52 28 53 32
rect 47 27 53 28
rect 57 32 63 33
rect 57 28 58 32
rect 62 28 63 32
rect 57 27 63 28
rect 67 32 73 33
rect 67 28 68 32
rect 72 28 73 32
rect 67 27 73 28
rect 88 32 92 58
rect 101 57 107 58
rect 101 32 107 33
rect 88 28 102 32
rect 106 28 107 32
rect 27 22 33 23
rect 27 18 28 22
rect 32 18 33 22
rect 3 17 9 18
rect 27 17 33 18
rect 39 22 45 23
rect 39 18 40 22
rect 44 18 45 22
rect 49 22 53 27
rect 58 22 62 23
rect 49 18 62 22
rect 39 17 45 18
rect 58 17 62 18
rect 75 22 81 23
rect 88 22 92 28
rect 101 27 107 28
rect 112 23 116 68
rect 124 68 126 72
rect 130 68 131 72
rect 124 67 131 68
rect 124 43 128 67
rect 121 42 128 43
rect 121 38 122 42
rect 126 38 128 42
rect 136 42 140 78
rect 147 78 148 82
rect 152 78 153 82
rect 147 72 153 78
rect 147 68 148 72
rect 152 68 153 72
rect 147 62 153 68
rect 147 58 148 62
rect 152 58 153 62
rect 147 57 153 58
rect 157 78 160 82
rect 164 78 165 82
rect 157 77 165 78
rect 171 82 177 87
rect 171 78 172 82
rect 176 78 177 82
rect 157 73 163 77
rect 157 72 165 73
rect 157 68 160 72
rect 164 68 165 72
rect 157 67 165 68
rect 171 72 177 78
rect 171 68 172 72
rect 176 68 177 72
rect 157 63 163 67
rect 157 62 165 63
rect 157 58 160 62
rect 164 58 165 62
rect 157 57 165 58
rect 171 62 177 68
rect 171 58 172 62
rect 176 58 177 62
rect 171 57 177 58
rect 145 52 151 53
rect 157 52 163 57
rect 145 48 146 52
rect 150 48 164 52
rect 145 47 151 48
rect 145 42 151 43
rect 136 38 146 42
rect 150 38 151 42
rect 121 37 127 38
rect 75 18 76 22
rect 80 18 92 22
rect 97 22 103 23
rect 111 22 117 23
rect 97 18 98 22
rect 102 18 112 22
rect 116 18 117 22
rect 75 17 81 18
rect 97 17 103 18
rect 111 17 117 18
rect 123 22 129 23
rect 136 22 140 38
rect 145 37 151 38
rect 145 32 151 33
rect 157 32 163 48
rect 145 28 146 32
rect 150 28 164 32
rect 145 27 151 28
rect 157 23 163 28
rect 123 18 124 22
rect 128 18 140 22
rect 147 22 153 23
rect 147 18 148 22
rect 152 18 153 22
rect 157 22 165 23
rect 157 18 160 22
rect 164 18 165 22
rect 123 17 129 18
rect 147 13 153 18
rect 159 17 165 18
rect 171 22 177 23
rect 171 18 172 22
rect 176 18 177 22
rect 171 13 177 18
rect -2 12 182 13
rect -2 8 16 12
rect 20 8 52 12
rect 56 8 100 12
rect 104 8 148 12
rect 152 8 172 12
rect 176 8 182 12
rect -2 4 28 8
rect 32 4 40 8
rect 44 4 64 8
rect 68 4 76 8
rect 80 4 124 8
rect 128 4 136 8
rect 140 4 182 8
rect -2 -1 182 4
<< ntransistor >>
rect 11 15 13 25
rect 23 15 25 25
rect 47 15 49 25
rect 59 15 61 25
rect 71 15 73 25
rect 83 15 85 25
rect 119 15 121 25
rect 131 15 133 25
rect 143 15 145 25
rect 95 5 97 15
rect 107 5 109 15
rect 155 5 157 25
rect 167 5 169 25
<< ptransistor >>
rect 11 65 13 85
rect 23 65 25 85
rect 47 75 49 95
rect 59 75 61 95
rect 71 65 73 85
rect 83 65 85 85
rect 95 75 97 95
rect 107 75 109 95
rect 119 75 121 95
rect 131 75 133 95
rect 143 75 145 95
rect 155 55 157 95
rect 167 55 169 95
<< polycontact >>
rect 48 68 52 72
rect 14 58 18 62
rect 4 48 8 52
rect 98 68 102 72
rect 38 58 42 62
rect 58 58 62 62
rect 68 58 72 62
rect 14 28 18 32
rect 68 48 72 52
rect 102 58 106 62
rect 126 68 130 72
rect 30 38 34 42
rect 78 38 82 42
rect 48 28 52 32
rect 58 28 62 32
rect 68 28 72 32
rect 122 38 126 42
rect 102 28 106 32
rect 98 18 102 22
rect 146 48 150 52
rect 146 38 150 42
rect 146 28 150 32
<< ndcontact >>
rect 4 18 8 22
rect 28 18 32 22
rect 40 18 44 22
rect 76 18 80 22
rect 112 18 116 22
rect 124 18 128 22
rect 148 18 152 22
rect 16 8 20 12
rect 52 8 56 12
rect 100 8 104 12
rect 148 8 152 12
rect 160 18 164 22
rect 172 18 176 22
rect 172 8 176 12
<< pdcontact >>
rect 16 88 20 92
rect 4 78 8 82
rect 4 68 8 72
rect 40 78 44 82
rect 52 88 56 92
rect 28 68 32 72
rect 76 68 80 72
rect 100 88 104 92
rect 112 78 116 82
rect 124 78 128 82
rect 148 88 152 92
rect 148 78 152 82
rect 148 68 152 72
rect 148 58 152 62
rect 160 78 164 82
rect 160 68 164 72
rect 160 58 164 62
rect 172 88 176 92
rect 172 78 176 82
rect 172 68 176 72
rect 172 58 176 62
<< psubstratepcontact >>
rect 28 4 32 8
rect 40 4 44 8
rect 64 4 68 8
rect 76 4 80 8
rect 124 4 128 8
rect 136 4 140 8
<< psubstratepdiff >>
rect 27 8 45 9
rect 27 4 28 8
rect 32 4 40 8
rect 44 4 45 8
rect 63 8 81 9
rect 27 3 45 4
rect 63 4 64 8
rect 68 4 76 8
rect 80 4 81 8
rect 123 8 141 9
rect 63 3 81 4
rect 123 4 124 8
rect 128 4 136 8
rect 140 4 141 8
rect 123 3 141 4
<< labels >>
rlabel metal1 20 50 20 50 6 ck
rlabel metal1 20 50 20 50 6 ck
rlabel metal1 60 20 60 20 6 i
rlabel metal1 60 20 60 20 6 i
rlabel metal1 50 50 50 50 6 i
rlabel metal1 50 50 50 50 6 i
rlabel metal1 60 80 60 80 6 i
rlabel metal1 60 80 60 80 6 i
rlabel metal1 90 6 90 6 6 vss
rlabel metal1 90 6 90 6 6 vss
rlabel metal1 90 94 90 94 6 vdd
rlabel metal1 90 94 90 94 6 vdd
rlabel metal1 160 50 160 50 6 q
rlabel metal1 160 50 160 50 6 q
<< end >>
