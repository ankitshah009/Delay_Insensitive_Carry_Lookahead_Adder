magic
tech scmos
timestamp 1185039050
<< checkpaint >>
rect -22 -24 92 124
<< ab >>
rect 0 0 70 100
<< pwell >>
rect -2 -4 72 49
<< nwell >>
rect -2 49 72 104
<< polysilicon >>
rect 11 95 13 98
rect 23 95 25 98
rect 35 95 37 98
rect 47 95 49 98
rect 11 43 13 55
rect 23 43 25 55
rect 7 42 13 43
rect 7 38 8 42
rect 12 38 13 42
rect 7 37 13 38
rect 17 42 25 43
rect 17 38 18 42
rect 22 38 25 42
rect 17 37 25 38
rect 11 25 13 37
rect 23 25 25 37
rect 35 43 37 55
rect 47 43 49 55
rect 35 42 43 43
rect 35 38 38 42
rect 42 38 43 42
rect 35 37 43 38
rect 47 42 53 43
rect 47 38 48 42
rect 52 38 53 42
rect 47 37 53 38
rect 35 25 37 37
rect 47 25 49 37
rect 11 2 13 5
rect 23 2 25 5
rect 35 2 37 5
rect 47 2 49 5
<< ndiffusion >>
rect 3 12 11 25
rect 3 8 4 12
rect 8 8 11 12
rect 3 5 11 8
rect 13 5 23 25
rect 25 22 35 25
rect 25 18 28 22
rect 32 18 35 22
rect 25 5 35 18
rect 37 5 47 25
rect 49 12 57 25
rect 49 8 52 12
rect 56 8 57 12
rect 49 5 57 8
<< pdiffusion >>
rect 3 82 11 95
rect 3 78 4 82
rect 8 78 11 82
rect 3 55 11 78
rect 13 72 23 95
rect 13 68 16 72
rect 20 68 23 72
rect 13 55 23 68
rect 25 82 35 95
rect 25 78 28 82
rect 32 78 35 82
rect 25 55 35 78
rect 37 92 47 95
rect 37 88 40 92
rect 44 88 47 92
rect 37 55 47 88
rect 49 82 57 95
rect 49 78 52 82
rect 56 78 57 82
rect 49 73 57 78
rect 49 55 55 73
<< metal1 >>
rect -2 92 72 101
rect -2 88 40 92
rect 44 88 72 92
rect -2 87 72 88
rect 3 82 9 83
rect 27 82 33 83
rect 51 82 57 83
rect 3 78 4 82
rect 8 78 28 82
rect 32 78 52 82
rect 56 78 57 82
rect 3 77 9 78
rect 27 77 33 78
rect 51 77 57 78
rect 15 72 33 73
rect 15 68 16 72
rect 20 68 33 72
rect 15 67 33 68
rect 7 42 13 62
rect 7 38 8 42
rect 12 38 13 42
rect 7 18 13 38
rect 17 42 23 62
rect 17 38 18 42
rect 22 38 23 42
rect 17 18 23 38
rect 27 22 33 67
rect 27 18 28 22
rect 32 18 33 22
rect 37 42 43 72
rect 37 38 38 42
rect 42 38 43 42
rect 37 18 43 38
rect 47 42 53 72
rect 61 60 67 87
rect 61 56 62 60
rect 66 56 67 60
rect 61 55 67 56
rect 47 38 48 42
rect 52 38 53 42
rect 47 18 53 38
rect 27 17 33 18
rect -2 12 72 13
rect -2 8 4 12
rect 8 8 52 12
rect 56 8 72 12
rect -2 -1 72 8
<< ntransistor >>
rect 11 5 13 25
rect 23 5 25 25
rect 35 5 37 25
rect 47 5 49 25
<< ptransistor >>
rect 11 55 13 95
rect 23 55 25 95
rect 35 55 37 95
rect 47 55 49 95
<< polycontact >>
rect 8 38 12 42
rect 18 38 22 42
rect 38 38 42 42
rect 48 38 52 42
<< ndcontact >>
rect 4 8 8 12
rect 28 18 32 22
rect 52 8 56 12
<< pdcontact >>
rect 4 78 8 82
rect 16 68 20 72
rect 28 78 32 82
rect 40 88 44 92
rect 52 78 56 82
<< nsubstratencontact >>
rect 62 56 66 60
<< nsubstratendiff >>
rect 61 60 67 67
rect 61 56 62 60
rect 66 56 67 60
rect 61 55 67 56
<< labels >>
rlabel polycontact 10 40 10 40 6 i0
rlabel polycontact 10 40 10 40 6 i0
rlabel metal1 30 45 30 45 6 nq
rlabel polycontact 20 40 20 40 6 i1
rlabel metal1 30 45 30 45 6 nq
rlabel polycontact 20 40 20 40 6 i1
rlabel metal1 35 6 35 6 6 vss
rlabel metal1 35 6 35 6 6 vss
rlabel metal1 50 45 50 45 6 i2
rlabel metal1 40 45 40 45 6 i3
rlabel metal1 50 45 50 45 6 i2
rlabel metal1 40 45 40 45 6 i3
rlabel metal1 35 94 35 94 6 vdd
rlabel metal1 35 94 35 94 6 vdd
<< end >>
