.subckt oai21a2v0x1 a1 a2 b vdd vss z
*   SPICE3 file   created from oai21a2v0x1.ext -      technology: scmos
m00 z      b      vdd    vdd p w=15u  l=2.3636u ad=64.5349p pd=25.1163u as=79.6721p ps=29.0164u
m01 w1     w2     z      vdd p w=28u  l=2.3636u ad=70p      pd=33u      as=120.465p ps=46.8837u
m02 vdd    a1     w1     vdd p w=28u  l=2.3636u ad=148.721p pd=54.1639u as=70p      ps=33u
m03 w2     a2     vdd    vdd p w=18u  l=2.3636u ad=116p     pd=50u      as=95.6066p ps=34.8197u
m04 n1     b      z      vss n w=13u  l=2.3636u ad=60.3333p pd=27.3333u as=77p      ps=40u
m05 vss    w2     n1     vss n w=13u  l=2.3636u ad=62.0286p pd=27.4857u as=60.3333p ps=27.3333u
m06 n1     a1     vss    vss n w=13u  l=2.3636u ad=60.3333p pd=27.3333u as=62.0286p ps=27.4857u
m07 vss    a2     w2     vss n w=9u   l=2.3636u ad=42.9429p pd=19.0286u as=57p      ps=32u
C0  a2     vdd    0.024f
C1  z      w2     0.091f
C2  vss    n1     0.198f
C3  a1     b      0.055f
C4  z      vdd    0.179f
C5  w2     vdd    0.122f
C6  vss    a1     0.031f
C7  n1     z      0.040f
C8  a2     a1     0.017f
C9  n1     w2     0.041f
C10 vss    b      0.033f
C11 n1     vdd    0.004f
C12 z      a1     0.015f
C13 w1     w2     0.007f
C14 a2     b      0.016f
C15 z      b      0.203f
C16 a1     w2     0.318f
C17 w1     vdd    0.005f
C18 vss    a2     0.017f
C19 w2     b      0.227f
C20 a1     vdd    0.021f
C21 vss    z      0.042f
C22 b      vdd    0.018f
C23 n1     a1     0.063f
C24 vss    w2     0.057f
C25 vss    vdd    0.006f
C26 a2     w2     0.103f
C27 n1     b      0.083f
C29 a2     vss    0.030f
C30 z      vss    0.017f
C31 a1     vss    0.026f
C32 w2     vss    0.030f
C33 b      vss    0.032f
.ends
