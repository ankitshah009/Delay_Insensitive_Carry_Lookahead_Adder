.subckt nd2v0x4 a b vdd vss z
*   SPICE3 file   created from nd2v0x4.ext -      technology: scmos
m00 z      a      vdd    vdd p w=28u  l=2.3636u ad=176p     pd=50u      as=196p     ps=70u
m01 vdd    a      z      vdd p w=28u  l=2.3636u ad=196p     pd=70u      as=176p     ps=50u
m02 z      b      vdd    vdd p w=28u  l=2.3636u ad=176p     pd=50u      as=196p     ps=70u
m03 vdd    b      z      vdd p w=28u  l=2.3636u ad=196p     pd=70u      as=176p     ps=50u
m04 w1     a      vss    vss n w=20u  l=2.3636u ad=138p     pd=48u      as=140p     ps=54u
m05 vss    a      w1     vss n w=20u  l=2.3636u ad=140p     pd=54u      as=138p     ps=48u
m06 z      b      w1     vss n w=20u  l=2.3636u ad=136p     pd=42u      as=138p     ps=48u
m07 w1     b      z      vss n w=20u  l=2.3636u ad=138p     pd=48u      as=136p     ps=42u
C0  b      a      0.152f
C1  vss    vdd    0.007f
C2  z      vdd    0.156f
C3  w1     vss    0.195f
C4  w1     z      0.139f
C5  vss    b      0.204f
C6  w1     vdd    0.012f
C7  vss    a      0.073f
C8  b      z      0.213f
C9  z      a      0.137f
C10 b      vdd    0.062f
C11 a      vdd    0.071f
C12 w1     b      0.126f
C13 w1     a      0.109f
C14 vss    z      0.019f
C15 w1     vss    0.002f
C17 b      vss    0.090f
C18 z      vss    0.008f
C19 a      vss    0.095f
.ends
