magic
tech scmos
timestamp 1179387562
<< checkpaint >>
rect -22 -25 206 105
<< ab >>
rect 0 0 184 80
<< pwell >>
rect -4 -7 188 36
<< nwell >>
rect -4 36 188 87
<< polysilicon >>
rect 9 69 11 74
rect 19 69 21 74
rect 29 72 53 74
rect 29 69 31 72
rect 39 69 41 72
rect 51 55 53 72
rect 63 70 65 74
rect 73 70 75 74
rect 83 70 85 74
rect 93 70 95 74
rect 116 70 118 74
rect 123 70 125 74
rect 133 70 135 74
rect 151 70 153 74
rect 161 70 163 74
rect 48 54 54 55
rect 48 50 49 54
rect 53 50 54 54
rect 48 49 54 50
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 39 39 41 42
rect 63 41 65 44
rect 73 41 75 44
rect 9 38 22 39
rect 9 37 17 38
rect 16 34 17 37
rect 21 34 22 38
rect 29 37 41 39
rect 61 39 75 41
rect 83 39 85 42
rect 93 39 95 42
rect 116 39 118 42
rect 61 38 67 39
rect 16 33 22 34
rect 9 28 11 33
rect 16 31 28 33
rect 16 28 18 31
rect 26 28 28 31
rect 33 28 35 37
rect 61 35 62 38
rect 45 30 47 35
rect 55 34 62 35
rect 66 34 67 38
rect 80 38 108 39
rect 80 37 103 38
rect 80 35 82 37
rect 55 33 67 34
rect 55 30 57 33
rect 65 30 67 33
rect 75 33 82 35
rect 102 34 103 37
rect 107 34 108 38
rect 102 33 108 34
rect 112 38 118 39
rect 112 34 113 38
rect 117 34 118 38
rect 123 39 125 42
rect 133 39 135 42
rect 151 39 153 42
rect 161 39 163 42
rect 123 36 126 39
rect 133 38 153 39
rect 133 37 138 38
rect 112 33 118 34
rect 75 30 77 33
rect 86 31 92 32
rect 86 27 87 31
rect 91 27 92 31
rect 114 30 116 33
rect 124 30 126 36
rect 137 34 138 37
rect 142 37 153 38
rect 157 38 163 39
rect 142 34 148 37
rect 137 33 148 34
rect 157 34 158 38
rect 162 34 163 38
rect 157 33 163 34
rect 146 30 148 33
rect 85 25 97 27
rect 85 22 87 25
rect 95 22 97 25
rect 9 8 11 16
rect 16 12 18 16
rect 26 12 28 16
rect 33 8 35 16
rect 9 6 35 8
rect 45 8 47 16
rect 55 12 57 16
rect 65 12 67 16
rect 75 8 77 16
rect 133 21 139 22
rect 133 17 134 21
rect 138 17 139 21
rect 158 27 160 33
rect 133 16 139 17
rect 45 6 77 8
rect 85 6 87 10
rect 95 6 97 10
rect 114 11 116 16
rect 124 13 126 16
rect 133 13 135 16
rect 146 14 148 19
rect 124 11 135 13
rect 158 11 160 16
<< ndiffusion >>
rect 37 28 45 30
rect 4 22 9 28
rect 2 21 9 22
rect 2 17 3 21
rect 7 17 9 21
rect 2 16 9 17
rect 11 16 16 28
rect 18 27 26 28
rect 18 23 20 27
rect 24 23 26 27
rect 18 16 26 23
rect 28 16 33 28
rect 35 16 45 28
rect 47 29 55 30
rect 47 25 49 29
rect 53 25 55 29
rect 47 16 55 25
rect 57 21 65 30
rect 57 17 59 21
rect 63 17 65 21
rect 57 16 65 17
rect 67 29 75 30
rect 67 25 69 29
rect 73 25 75 29
rect 67 22 75 25
rect 67 18 69 22
rect 73 18 75 22
rect 67 16 75 18
rect 77 22 82 30
rect 109 23 114 30
rect 107 22 114 23
rect 77 21 85 22
rect 77 17 79 21
rect 83 17 85 21
rect 77 16 85 17
rect 37 12 43 16
rect 37 8 38 12
rect 42 8 43 12
rect 37 7 43 8
rect 80 10 85 16
rect 87 21 95 22
rect 87 17 89 21
rect 93 17 95 21
rect 87 10 95 17
rect 97 13 103 22
rect 107 18 108 22
rect 112 18 114 22
rect 107 17 114 18
rect 109 16 114 17
rect 116 29 124 30
rect 116 25 118 29
rect 122 25 124 29
rect 116 16 124 25
rect 126 29 133 30
rect 126 25 128 29
rect 132 25 133 29
rect 126 24 133 25
rect 139 29 146 30
rect 139 25 140 29
rect 144 25 146 29
rect 139 24 146 25
rect 126 16 131 24
rect 141 19 146 24
rect 148 27 156 30
rect 148 19 158 27
rect 97 12 105 13
rect 97 10 100 12
rect 99 8 100 10
rect 104 8 105 12
rect 150 16 158 19
rect 160 22 165 27
rect 160 21 167 22
rect 160 17 162 21
rect 166 17 167 21
rect 160 16 167 17
rect 150 12 156 16
rect 99 7 105 8
rect 150 8 151 12
rect 155 8 156 12
rect 150 7 156 8
<< pdiffusion >>
rect 4 63 9 69
rect 2 62 9 63
rect 2 58 3 62
rect 7 58 9 62
rect 2 55 9 58
rect 2 51 3 55
rect 7 51 9 55
rect 2 50 9 51
rect 4 42 9 50
rect 11 54 19 69
rect 11 50 13 54
rect 17 50 19 54
rect 11 47 19 50
rect 11 43 13 47
rect 17 43 19 47
rect 11 42 19 43
rect 21 62 29 69
rect 21 58 23 62
rect 27 58 29 62
rect 21 42 29 58
rect 31 47 39 69
rect 31 43 33 47
rect 37 43 39 47
rect 31 42 39 43
rect 41 63 46 69
rect 41 62 48 63
rect 41 58 43 62
rect 47 58 48 62
rect 41 57 48 58
rect 41 42 46 57
rect 56 69 63 70
rect 56 65 57 69
rect 61 65 63 69
rect 56 62 63 65
rect 56 58 57 62
rect 61 58 63 62
rect 56 44 63 58
rect 65 62 73 70
rect 65 58 67 62
rect 71 58 73 62
rect 65 55 73 58
rect 65 51 67 55
rect 71 51 73 55
rect 65 44 73 51
rect 75 69 83 70
rect 75 65 77 69
rect 81 65 83 69
rect 75 44 83 65
rect 78 42 83 44
rect 85 49 93 70
rect 85 45 87 49
rect 91 45 93 49
rect 85 42 93 45
rect 95 69 116 70
rect 95 65 97 69
rect 101 65 105 69
rect 109 65 116 69
rect 95 62 116 65
rect 95 58 105 62
rect 109 58 116 62
rect 95 42 116 58
rect 118 42 123 70
rect 125 63 133 70
rect 125 59 127 63
rect 131 59 133 63
rect 125 42 133 59
rect 135 64 140 70
rect 135 63 142 64
rect 135 59 137 63
rect 141 59 142 63
rect 135 58 142 59
rect 135 42 140 58
rect 146 54 151 70
rect 144 53 151 54
rect 144 49 145 53
rect 149 49 151 53
rect 144 48 151 49
rect 146 42 151 48
rect 153 69 161 70
rect 153 65 155 69
rect 159 65 161 69
rect 153 42 161 65
rect 163 55 168 70
rect 163 54 170 55
rect 163 50 165 54
rect 169 50 170 54
rect 163 47 170 50
rect 163 43 165 47
rect 169 43 170 47
rect 163 42 170 43
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect 118 78 122 82
rect 126 78 130 82
rect 134 78 138 82
rect 142 78 146 82
rect 150 78 154 82
rect 158 78 162 82
rect 166 78 170 82
rect 174 78 178 82
rect 182 78 186 82
rect -2 69 186 78
rect -2 68 57 69
rect 56 65 57 68
rect 61 68 77 69
rect 61 65 62 68
rect 56 62 62 65
rect 81 68 97 69
rect 77 64 81 65
rect 101 68 105 69
rect 97 64 101 65
rect 109 68 155 69
rect 154 65 155 68
rect 159 68 186 69
rect 159 65 160 68
rect 2 58 3 62
rect 7 58 23 62
rect 27 58 43 62
rect 47 58 48 62
rect 56 58 57 62
rect 61 58 62 62
rect 67 62 71 63
rect 105 62 109 65
rect 2 55 7 58
rect 2 51 3 55
rect 67 55 99 58
rect 105 57 109 58
rect 113 59 127 63
rect 131 59 132 63
rect 136 59 137 63
rect 141 62 142 63
rect 141 59 169 62
rect 2 50 7 51
rect 12 50 13 54
rect 17 50 49 54
rect 53 51 67 54
rect 71 54 99 55
rect 53 50 71 51
rect 2 30 6 50
rect 12 47 17 50
rect 87 49 91 50
rect 12 43 13 47
rect 12 42 17 43
rect 32 43 33 47
rect 37 43 38 47
rect 32 38 38 43
rect 48 45 87 46
rect 48 42 91 45
rect 48 38 52 42
rect 16 34 17 38
rect 21 34 52 38
rect 57 34 62 38
rect 66 34 87 38
rect 2 27 24 30
rect 2 26 20 27
rect 48 29 52 34
rect 81 32 87 34
rect 81 31 91 32
rect 48 25 49 29
rect 53 25 69 29
rect 73 25 74 29
rect 81 27 87 31
rect 81 26 91 27
rect 20 22 24 23
rect 69 22 74 25
rect 3 21 7 22
rect 20 21 64 22
rect 20 18 59 21
rect 58 17 59 18
rect 63 17 64 21
rect 73 18 74 22
rect 95 21 99 54
rect 113 53 117 59
rect 136 58 169 59
rect 103 49 117 53
rect 121 49 145 53
rect 149 49 150 53
rect 103 38 107 49
rect 121 38 125 49
rect 129 42 142 46
rect 138 38 142 42
rect 154 39 158 55
rect 165 54 169 58
rect 165 47 169 50
rect 112 34 113 38
rect 117 34 131 38
rect 103 29 107 34
rect 127 29 131 34
rect 138 33 142 34
rect 146 38 162 39
rect 146 34 158 38
rect 146 33 162 34
rect 103 25 118 29
rect 122 25 123 29
rect 127 25 128 29
rect 132 25 140 29
rect 144 25 145 29
rect 154 25 158 33
rect 69 17 74 18
rect 78 17 79 21
rect 83 17 84 21
rect 88 17 89 21
rect 93 17 99 21
rect 107 18 108 22
rect 112 21 113 22
rect 165 21 169 43
rect 112 18 134 21
rect 107 17 134 18
rect 138 17 162 21
rect 166 17 169 21
rect 3 12 7 17
rect 78 12 84 17
rect -2 8 38 12
rect 42 8 100 12
rect 104 8 151 12
rect 155 8 186 12
rect -2 2 186 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 122 2
rect 126 -2 130 2
rect 134 -2 138 2
rect 142 -2 146 2
rect 150 -2 154 2
rect 158 -2 162 2
rect 166 -2 170 2
rect 174 -2 178 2
rect 182 -2 186 2
<< ntransistor >>
rect 9 16 11 28
rect 16 16 18 28
rect 26 16 28 28
rect 33 16 35 28
rect 45 16 47 30
rect 55 16 57 30
rect 65 16 67 30
rect 75 16 77 30
rect 85 10 87 22
rect 95 10 97 22
rect 114 16 116 30
rect 124 16 126 30
rect 146 19 148 30
rect 158 16 160 27
<< ptransistor >>
rect 9 42 11 69
rect 19 42 21 69
rect 29 42 31 69
rect 39 42 41 69
rect 63 44 65 70
rect 73 44 75 70
rect 83 42 85 70
rect 93 42 95 70
rect 116 42 118 70
rect 123 42 125 70
rect 133 42 135 70
rect 151 42 153 70
rect 161 42 163 70
<< polycontact >>
rect 49 50 53 54
rect 17 34 21 38
rect 62 34 66 38
rect 103 34 107 38
rect 113 34 117 38
rect 87 27 91 31
rect 138 34 142 38
rect 158 34 162 38
rect 134 17 138 21
<< ndcontact >>
rect 3 17 7 21
rect 20 23 24 27
rect 49 25 53 29
rect 59 17 63 21
rect 69 25 73 29
rect 69 18 73 22
rect 79 17 83 21
rect 38 8 42 12
rect 89 17 93 21
rect 108 18 112 22
rect 118 25 122 29
rect 128 25 132 29
rect 140 25 144 29
rect 100 8 104 12
rect 162 17 166 21
rect 151 8 155 12
<< pdcontact >>
rect 3 58 7 62
rect 3 51 7 55
rect 13 50 17 54
rect 13 43 17 47
rect 23 58 27 62
rect 33 43 37 47
rect 43 58 47 62
rect 57 65 61 69
rect 57 58 61 62
rect 67 58 71 62
rect 67 51 71 55
rect 77 65 81 69
rect 87 45 91 49
rect 97 65 101 69
rect 105 65 109 69
rect 105 58 109 62
rect 127 59 131 63
rect 137 59 141 63
rect 145 49 149 53
rect 155 65 159 69
rect 165 50 169 54
rect 165 43 169 47
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
rect 90 -2 94 2
rect 98 -2 102 2
rect 106 -2 110 2
rect 114 -2 118 2
rect 122 -2 126 2
rect 130 -2 134 2
rect 138 -2 142 2
rect 146 -2 150 2
rect 154 -2 158 2
rect 162 -2 166 2
rect 170 -2 174 2
rect 178 -2 182 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
rect 90 78 94 82
rect 98 78 102 82
rect 106 78 110 82
rect 114 78 118 82
rect 122 78 126 82
rect 130 78 134 82
rect 138 78 142 82
rect 146 78 150 82
rect 154 78 158 82
rect 162 78 166 82
rect 170 78 174 82
rect 178 78 182 82
<< psubstratepdiff >>
rect 0 2 184 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 122 2
rect 126 -2 130 2
rect 134 -2 138 2
rect 142 -2 146 2
rect 150 -2 154 2
rect 158 -2 162 2
rect 166 -2 170 2
rect 174 -2 178 2
rect 182 -2 184 2
rect 0 -3 184 -2
<< nsubstratendiff >>
rect 0 82 184 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect 118 78 122 82
rect 126 78 130 82
rect 134 78 138 82
rect 142 78 146 82
rect 150 78 154 82
rect 158 78 162 82
rect 166 78 170 82
rect 174 78 178 82
rect 182 78 184 82
rect 0 77 184 78
<< labels >>
rlabel ptransistor 20 52 20 52 6 zn
rlabel polysilicon 52 61 52 61 6 cn
rlabel ntransistor 115 25 115 25 6 bn
rlabel polycontact 105 36 105 36 6 iz
rlabel polycontact 136 19 136 19 6 an
rlabel metal1 12 28 12 28 6 z
rlabel metal1 20 28 20 28 6 z
rlabel metal1 4 44 4 44 6 z
rlabel metal1 14 48 14 48 6 cn
rlabel metal1 20 60 20 60 6 z
rlabel metal1 12 60 12 60 6 z
rlabel metal1 28 20 28 20 6 z
rlabel metal1 52 20 52 20 6 z
rlabel metal1 44 20 44 20 6 z
rlabel metal1 36 20 36 20 6 z
rlabel metal1 35 40 35 40 6 zn
rlabel metal1 28 60 28 60 6 z
rlabel pdcontact 44 60 44 60 6 z
rlabel metal1 36 60 36 60 6 z
rlabel ndcontact 60 20 60 20 6 z
rlabel metal1 71 23 71 23 6 zn
rlabel metal1 61 27 61 27 6 zn
rlabel metal1 60 36 60 36 6 c
rlabel metal1 76 36 76 36 6 c
rlabel metal1 84 32 84 32 6 c
rlabel metal1 68 36 68 36 6 c
rlabel metal1 69 44 69 44 6 zn
rlabel metal1 41 52 41 52 6 cn
rlabel metal1 92 6 92 6 6 vss
rlabel metal1 93 19 93 19 6 cn
rlabel metal1 105 39 105 39 6 iz
rlabel metal1 83 56 83 56 6 cn
rlabel metal1 92 74 92 74 6 vdd
rlabel metal1 136 27 136 27 6 bn
rlabel metal1 113 27 113 27 6 iz
rlabel metal1 148 36 148 36 6 a
rlabel polycontact 140 36 140 36 6 b
rlabel metal1 132 44 132 44 6 b
rlabel metal1 123 43 123 43 6 bn
rlabel metal1 135 51 135 51 6 bn
rlabel metal1 122 61 122 61 6 iz
rlabel metal1 138 19 138 19 6 an
rlabel metal1 156 28 156 28 6 a
rlabel metal1 156 40 156 40 6 a
rlabel metal1 167 39 167 39 6 an
rlabel metal1 152 60 152 60 6 an
<< end >>
