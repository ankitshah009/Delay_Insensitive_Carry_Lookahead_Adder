magic
tech scmos
timestamp 1179385271
<< checkpaint >>
rect -22 -25 62 105
<< ab >>
rect 0 0 40 80
<< pwell >>
rect -4 -7 44 36
<< nwell >>
rect -4 36 44 87
<< polysilicon >>
rect 9 69 11 74
rect 19 69 21 74
rect 29 69 31 74
rect 9 39 11 42
rect 19 39 21 42
rect 9 38 15 39
rect 9 34 10 38
rect 14 34 15 38
rect 9 33 15 34
rect 19 38 25 39
rect 19 34 20 38
rect 24 34 25 38
rect 19 33 25 34
rect 10 22 12 33
rect 20 22 22 33
rect 29 31 31 42
rect 29 30 35 31
rect 29 28 30 30
rect 27 26 30 28
rect 34 26 35 30
rect 27 25 35 26
rect 27 22 29 25
rect 10 10 12 15
rect 20 6 22 10
rect 27 6 29 10
<< ndiffusion >>
rect 2 15 10 22
rect 12 21 20 22
rect 12 17 14 21
rect 18 17 20 21
rect 12 15 20 17
rect 2 12 8 15
rect 2 8 3 12
rect 7 8 8 12
rect 15 10 20 15
rect 22 10 27 22
rect 29 12 38 22
rect 29 10 32 12
rect 2 7 8 8
rect 31 8 32 10
rect 36 8 38 12
rect 31 7 38 8
<< pdiffusion >>
rect 4 63 9 69
rect 2 62 9 63
rect 2 58 3 62
rect 7 58 9 62
rect 2 55 9 58
rect 2 51 3 55
rect 7 51 9 55
rect 2 50 9 51
rect 4 42 9 50
rect 11 62 19 69
rect 11 58 13 62
rect 17 58 19 62
rect 11 55 19 58
rect 11 51 13 55
rect 17 51 19 55
rect 11 42 19 51
rect 21 68 29 69
rect 21 64 23 68
rect 27 64 29 68
rect 21 61 29 64
rect 21 57 23 61
rect 27 57 29 61
rect 21 42 29 57
rect 31 63 36 69
rect 31 62 38 63
rect 31 58 33 62
rect 37 58 38 62
rect 31 55 38 58
rect 31 51 33 55
rect 37 51 38 55
rect 31 50 38 51
rect 31 42 36 50
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect -2 68 42 78
rect 22 64 23 68
rect 27 64 28 68
rect 2 62 8 63
rect 2 58 3 62
rect 7 58 8 62
rect 2 55 8 58
rect 2 51 3 55
rect 7 51 8 55
rect 13 62 17 63
rect 13 55 17 58
rect 22 61 28 64
rect 22 57 23 61
rect 27 57 28 61
rect 33 62 37 63
rect 33 55 37 58
rect 17 51 33 54
rect 2 22 6 51
rect 13 50 37 51
rect 10 42 23 47
rect 10 38 14 42
rect 34 38 38 47
rect 19 34 20 38
rect 24 34 38 38
rect 10 33 14 34
rect 25 26 30 30
rect 2 21 23 22
rect 2 17 14 21
rect 18 17 23 21
rect 34 17 38 30
rect -2 8 3 12
rect 7 8 32 12
rect 36 8 42 12
rect -2 2 42 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
<< ntransistor >>
rect 10 15 12 22
rect 20 10 22 22
rect 27 10 29 22
<< ptransistor >>
rect 9 42 11 69
rect 19 42 21 69
rect 29 42 31 69
<< polycontact >>
rect 10 34 14 38
rect 20 34 24 38
rect 30 26 34 30
<< ndcontact >>
rect 14 17 18 21
rect 3 8 7 12
rect 32 8 36 12
<< pdcontact >>
rect 3 58 7 62
rect 3 51 7 55
rect 13 58 17 62
rect 13 51 17 55
rect 23 64 27 68
rect 23 57 27 61
rect 33 58 37 62
rect 33 51 37 55
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
<< psubstratepdiff >>
rect 0 2 40 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 40 2
rect 0 -3 40 -2
<< nsubstratendiff >>
rect 0 82 40 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 40 82
rect 0 77 40 78
<< labels >>
rlabel metal1 4 40 4 40 6 z
rlabel metal1 12 20 12 20 6 z
rlabel metal1 12 40 12 40 6 b
rlabel metal1 15 56 15 56 6 n1
rlabel metal1 20 6 20 6 6 vss
rlabel metal1 20 20 20 20 6 z
rlabel metal1 28 36 28 36 6 a2
rlabel metal1 28 28 28 28 6 a1
rlabel metal1 20 44 20 44 6 b
rlabel metal1 20 74 20 74 6 vdd
rlabel metal1 36 20 36 20 6 a1
rlabel metal1 36 44 36 44 6 a2
rlabel metal1 35 56 35 56 6 n1
<< end >>
