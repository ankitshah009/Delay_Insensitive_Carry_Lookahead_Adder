.subckt xor2v0x05 a b vdd vss z
*   SPICE3 file   created from xor2v0x05.ext -      technology: scmos
m00 vdd    b      bn     vdd p w=21u  l=2.3636u ad=145.765p pd=40.7647u as=124p     ps=56u
m01 an     a      vdd    vdd p w=13u  l=2.3636u ad=52p      pd=21u      as=90.2353p ps=25.2353u
m02 z      bn     an     vdd p w=13u  l=2.3636u ad=55.0588p pd=22.1765u as=52p      ps=21u
m03 bn     an     z      vdd p w=21u  l=2.3636u ad=124p     pd=56u      as=88.9412p ps=35.8235u
m04 vss    b      bn     vss n w=7u   l=2.3636u ad=55.3913p pd=24.3478u as=49p      ps=28u
m05 an     a      vss    vss n w=7u   l=2.3636u ad=28p      pd=15u      as=55.3913p ps=24.3478u
m06 z      b      an     vss n w=7u   l=2.3636u ad=28.875p  pd=14.875u  as=28p      ps=15u
m07 w1     bn     z      vss n w=9u   l=2.3636u ad=22.5p    pd=14u      as=37.125p  ps=19.125u
m08 vss    an     w1     vss n w=9u   l=2.3636u ad=71.2174p pd=31.3043u as=22.5p    ps=14u
C0  vss    an     0.088f
C1  z      a      0.013f
C2  a      an     0.075f
C3  z      bn     0.164f
C4  vss    b      0.016f
C5  a      b      0.071f
C6  an     bn     0.165f
C7  z      vdd    0.032f
C8  bn     b      0.114f
C9  an     vdd    0.029f
C10 w1     z      0.011f
C11 b      vdd    0.113f
C12 vss    a      0.069f
C13 z      an     0.287f
C14 vss    bn     0.040f
C15 a      bn     0.142f
C16 z      b      0.004f
C17 an     b      0.026f
C18 a      vdd    0.017f
C19 bn     vdd    0.320f
C20 vss    z      0.148f
C22 z      vss    0.013f
C23 a      vss    0.024f
C24 an     vss    0.032f
C25 bn     vss    0.034f
C26 b      vss    0.052f
.ends
