magic
tech scmos
timestamp 1179385108
<< checkpaint >>
rect -22 -25 78 105
<< ab >>
rect 0 0 56 80
<< pwell >>
rect -4 -7 60 36
<< nwell >>
rect -4 36 60 87
<< polysilicon >>
rect 9 70 11 74
rect 19 67 21 72
rect 29 67 31 72
rect 41 67 43 72
rect 19 47 21 58
rect 29 55 31 58
rect 29 54 37 55
rect 29 50 32 54
rect 36 50 37 54
rect 29 49 37 50
rect 19 46 25 47
rect 19 42 20 46
rect 24 42 25 46
rect 9 39 11 42
rect 19 41 25 42
rect 9 38 15 39
rect 9 34 10 38
rect 14 34 15 38
rect 9 33 15 34
rect 9 30 11 33
rect 22 26 24 41
rect 29 26 31 49
rect 41 35 43 58
rect 40 34 46 35
rect 40 31 41 34
rect 36 30 41 31
rect 45 30 46 34
rect 36 29 46 30
rect 36 26 38 29
rect 9 12 11 16
rect 22 12 24 17
rect 29 12 31 17
rect 36 12 38 17
<< ndiffusion >>
rect 4 23 9 30
rect 2 22 9 23
rect 2 18 3 22
rect 7 18 9 22
rect 2 16 9 18
rect 11 26 20 30
rect 11 17 22 26
rect 24 17 29 26
rect 31 17 36 26
rect 38 23 43 26
rect 38 22 45 23
rect 38 18 40 22
rect 44 18 45 22
rect 38 17 45 18
rect 11 16 20 17
rect 13 12 20 16
rect 13 8 14 12
rect 18 8 20 12
rect 13 7 20 8
<< pdiffusion >>
rect 33 72 39 73
rect 4 55 9 70
rect 2 54 9 55
rect 2 50 3 54
rect 7 50 9 54
rect 2 47 9 50
rect 2 43 3 47
rect 7 43 9 47
rect 2 42 9 43
rect 11 67 16 70
rect 33 68 34 72
rect 38 68 39 72
rect 33 67 39 68
rect 11 66 19 67
rect 11 62 13 66
rect 17 62 19 66
rect 11 58 19 62
rect 21 63 29 67
rect 21 59 23 63
rect 27 59 29 63
rect 21 58 29 59
rect 31 58 41 67
rect 43 64 48 67
rect 43 63 50 64
rect 43 59 45 63
rect 49 59 50 63
rect 43 58 50 59
rect 11 42 17 58
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect -2 72 58 78
rect -2 68 34 72
rect 38 68 58 72
rect 13 66 17 68
rect 2 54 7 63
rect 13 61 17 62
rect 22 59 23 63
rect 27 59 45 63
rect 49 59 50 63
rect 22 54 26 59
rect 2 50 3 54
rect 2 47 7 50
rect 2 43 3 47
rect 2 42 7 43
rect 10 50 26 54
rect 31 50 32 54
rect 36 50 47 54
rect 2 22 6 42
rect 10 38 14 50
rect 17 42 20 46
rect 24 42 31 46
rect 41 42 47 50
rect 25 34 31 42
rect 41 34 47 38
rect 10 30 14 34
rect 45 30 47 34
rect 10 26 22 30
rect 25 26 47 30
rect 18 22 22 26
rect 2 18 3 22
rect 7 18 15 22
rect 18 18 40 22
rect 44 18 45 22
rect -2 8 14 12
rect 18 8 58 12
rect -2 2 58 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
<< ntransistor >>
rect 9 16 11 30
rect 22 17 24 26
rect 29 17 31 26
rect 36 17 38 26
<< ptransistor >>
rect 9 42 11 70
rect 19 58 21 67
rect 29 58 31 67
rect 41 58 43 67
<< polycontact >>
rect 32 50 36 54
rect 20 42 24 46
rect 10 34 14 38
rect 41 30 45 34
<< ndcontact >>
rect 3 18 7 22
rect 40 18 44 22
rect 14 8 18 12
<< pdcontact >>
rect 3 50 7 54
rect 3 43 7 47
rect 34 68 38 72
rect 13 62 17 66
rect 23 59 27 63
rect 45 59 49 63
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
<< psubstratepdiff >>
rect 0 2 56 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 56 2
rect 0 -3 56 -2
<< nsubstratendiff >>
rect 0 82 56 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 56 82
rect 0 77 56 78
<< labels >>
rlabel polycontact 12 36 12 36 6 zn
rlabel pdcontact 4 44 4 44 6 z
rlabel metal1 12 20 12 20 6 z
rlabel metal1 20 44 20 44 6 a
rlabel metal1 12 40 12 40 6 zn
rlabel metal1 28 6 28 6 6 vss
rlabel metal1 28 28 28 28 6 c
rlabel metal1 36 28 36 28 6 c
rlabel metal1 28 40 28 40 6 a
rlabel metal1 36 52 36 52 6 b
rlabel metal1 28 74 28 74 6 vdd
rlabel metal1 31 20 31 20 6 zn
rlabel polycontact 44 32 44 32 6 c
rlabel metal1 44 48 44 48 6 b
rlabel metal1 36 61 36 61 6 zn
<< end >>
