magic
tech scmos
timestamp 1185039076
<< checkpaint >>
rect -22 -24 152 124
<< ab >>
rect 0 0 130 100
<< pwell >>
rect -2 -4 132 49
<< nwell >>
rect -2 49 132 104
<< polysilicon >>
rect 23 95 25 98
rect 35 95 37 98
rect 11 79 13 82
rect 47 85 49 88
rect 59 85 61 88
rect 71 85 73 88
rect 83 85 85 88
rect 97 85 99 88
rect 107 85 109 88
rect 117 85 119 88
rect 11 43 13 55
rect 23 53 25 55
rect 35 53 37 55
rect 17 52 37 53
rect 17 48 18 52
rect 22 51 37 52
rect 22 48 23 51
rect 17 47 23 48
rect 47 43 49 63
rect 59 43 61 63
rect 71 43 73 63
rect 83 43 85 61
rect 11 42 43 43
rect 11 41 38 42
rect 11 29 13 41
rect 37 38 38 41
rect 42 38 43 42
rect 37 37 43 38
rect 47 42 53 43
rect 47 38 48 42
rect 52 38 53 42
rect 47 37 53 38
rect 57 42 63 43
rect 57 38 58 42
rect 62 38 63 42
rect 57 37 63 38
rect 67 42 73 43
rect 67 38 68 42
rect 72 38 73 42
rect 67 37 73 38
rect 77 42 85 43
rect 77 38 78 42
rect 82 38 85 42
rect 97 53 99 55
rect 107 53 109 55
rect 97 52 103 53
rect 97 48 98 52
rect 102 48 103 52
rect 97 47 103 48
rect 107 52 113 53
rect 107 48 108 52
rect 112 48 113 52
rect 107 47 113 48
rect 97 39 99 47
rect 107 39 109 47
rect 77 37 85 38
rect 93 37 99 39
rect 105 37 109 39
rect 117 43 119 55
rect 117 42 123 43
rect 117 38 118 42
rect 122 38 123 42
rect 117 37 123 38
rect 17 36 23 37
rect 17 32 18 36
rect 22 33 23 36
rect 49 33 51 37
rect 59 33 61 37
rect 69 33 71 37
rect 22 32 37 33
rect 17 31 37 32
rect 23 29 25 31
rect 35 29 37 31
rect 11 12 13 15
rect 81 29 83 37
rect 93 25 95 37
rect 105 25 107 37
rect 117 25 119 37
rect 49 14 51 17
rect 59 14 61 17
rect 69 14 71 17
rect 81 14 83 17
rect 93 14 95 17
rect 23 6 25 9
rect 35 6 37 9
rect 105 14 107 17
rect 117 14 119 17
<< ndiffusion >>
rect 41 29 49 33
rect 3 26 11 29
rect 3 22 4 26
rect 8 22 11 26
rect 3 15 11 22
rect 13 26 23 29
rect 13 22 16 26
rect 20 22 23 26
rect 13 16 23 22
rect 13 15 16 16
rect 15 12 16 15
rect 20 12 23 16
rect 15 9 23 12
rect 25 22 35 29
rect 25 18 28 22
rect 32 18 35 22
rect 25 9 35 18
rect 37 17 49 29
rect 51 17 59 33
rect 61 17 69 33
rect 71 29 75 33
rect 71 22 81 29
rect 71 18 74 22
rect 78 18 81 22
rect 71 17 81 18
rect 83 25 90 29
rect 83 22 93 25
rect 83 18 86 22
rect 90 18 93 22
rect 83 17 93 18
rect 95 17 105 25
rect 107 22 117 25
rect 107 18 110 22
rect 114 18 117 22
rect 107 17 117 18
rect 119 22 127 25
rect 119 18 122 22
rect 126 18 127 22
rect 119 17 127 18
rect 37 12 47 17
rect 37 9 42 12
rect 41 8 42 9
rect 46 8 47 12
rect 97 12 103 17
rect 41 7 47 8
rect 97 8 98 12
rect 102 8 103 12
rect 97 7 103 8
<< pdiffusion >>
rect 15 92 23 95
rect 15 88 16 92
rect 20 88 23 92
rect 15 82 23 88
rect 15 79 16 82
rect 3 72 11 79
rect 3 68 4 72
rect 8 68 11 72
rect 3 62 11 68
rect 3 58 4 62
rect 8 58 11 62
rect 3 55 11 58
rect 13 78 16 79
rect 20 78 23 82
rect 13 72 23 78
rect 13 68 16 72
rect 20 68 23 72
rect 13 62 23 68
rect 13 58 16 62
rect 20 58 23 62
rect 13 55 23 58
rect 25 82 35 95
rect 25 78 28 82
rect 32 78 35 82
rect 25 72 35 78
rect 25 68 28 72
rect 32 68 35 72
rect 25 62 35 68
rect 25 58 28 62
rect 32 58 35 62
rect 25 55 35 58
rect 37 85 44 95
rect 63 92 69 93
rect 63 88 64 92
rect 68 88 69 92
rect 63 85 69 88
rect 37 82 47 85
rect 37 78 40 82
rect 44 78 47 82
rect 37 63 47 78
rect 49 82 59 85
rect 49 78 52 82
rect 56 78 59 82
rect 49 63 59 78
rect 61 63 71 85
rect 73 82 83 85
rect 73 78 76 82
rect 80 78 83 82
rect 73 63 83 78
rect 37 55 44 63
rect 76 61 83 63
rect 85 72 97 85
rect 85 68 88 72
rect 92 68 97 72
rect 85 62 97 68
rect 85 61 88 62
rect 87 58 88 61
rect 92 58 97 62
rect 87 55 97 58
rect 99 55 107 85
rect 109 55 117 85
rect 119 82 127 85
rect 119 78 122 82
rect 126 78 127 82
rect 119 55 127 78
<< metal1 >>
rect -2 96 132 101
rect -2 92 4 96
rect 8 92 76 96
rect 80 92 88 96
rect 92 92 100 96
rect 104 92 112 96
rect 116 92 132 96
rect -2 88 16 92
rect 20 88 64 92
rect 68 88 132 92
rect -2 87 132 88
rect 15 82 21 87
rect 15 78 16 82
rect 20 78 21 82
rect 3 72 9 73
rect 3 68 4 72
rect 8 68 9 72
rect 3 67 9 68
rect 15 72 21 78
rect 15 68 16 72
rect 20 68 21 72
rect 4 63 8 67
rect 3 62 9 63
rect 3 58 4 62
rect 8 58 9 62
rect 3 57 9 58
rect 15 62 21 68
rect 15 58 16 62
rect 20 58 21 62
rect 15 57 21 58
rect 27 82 33 83
rect 27 78 28 82
rect 32 78 33 82
rect 27 72 33 78
rect 39 82 45 87
rect 39 78 40 82
rect 44 78 45 82
rect 39 77 45 78
rect 51 82 57 83
rect 75 82 81 83
rect 121 82 127 83
rect 51 78 52 82
rect 56 78 76 82
rect 80 78 122 82
rect 126 78 127 82
rect 51 77 57 78
rect 75 77 81 78
rect 121 77 127 78
rect 87 72 93 73
rect 27 68 28 72
rect 32 68 33 72
rect 27 62 33 68
rect 27 58 28 62
rect 32 58 33 62
rect 4 52 8 57
rect 17 52 23 53
rect 4 48 18 52
rect 22 48 23 52
rect 4 36 8 48
rect 17 47 23 48
rect 17 36 23 37
rect 4 32 18 36
rect 22 32 23 36
rect 4 27 8 32
rect 17 31 23 32
rect 3 26 9 27
rect 3 22 4 26
rect 8 22 9 26
rect 3 21 9 22
rect 15 26 21 27
rect 15 22 16 26
rect 20 22 21 26
rect 15 16 21 22
rect 27 22 33 58
rect 37 42 43 43
rect 37 38 38 42
rect 42 38 43 42
rect 37 37 43 38
rect 47 42 53 72
rect 47 38 48 42
rect 52 38 53 42
rect 27 18 28 22
rect 32 18 33 22
rect 38 22 42 37
rect 47 28 53 38
rect 57 42 63 72
rect 57 38 58 42
rect 62 38 63 42
rect 57 28 63 38
rect 67 42 73 72
rect 67 38 68 42
rect 72 38 73 42
rect 67 37 73 38
rect 77 42 83 72
rect 87 68 88 72
rect 92 68 93 72
rect 87 67 93 68
rect 88 63 92 67
rect 87 62 93 63
rect 87 58 88 62
rect 92 58 93 62
rect 87 57 93 58
rect 77 38 78 42
rect 82 38 83 42
rect 77 37 83 38
rect 88 32 92 57
rect 74 28 92 32
rect 97 52 103 72
rect 97 48 98 52
rect 102 48 103 52
rect 97 28 103 48
rect 107 52 113 72
rect 107 48 108 52
rect 112 48 113 52
rect 107 28 113 48
rect 117 42 123 72
rect 117 38 118 42
rect 122 38 123 42
rect 117 28 123 38
rect 74 23 78 28
rect 73 22 79 23
rect 38 18 74 22
rect 78 18 79 22
rect 27 17 33 18
rect 73 17 79 18
rect 85 22 91 23
rect 109 22 115 23
rect 85 18 86 22
rect 90 18 110 22
rect 114 18 115 22
rect 85 17 91 18
rect 109 17 115 18
rect 121 22 127 23
rect 121 18 122 22
rect 126 18 127 22
rect 15 13 16 16
rect -2 12 16 13
rect 20 13 21 16
rect 121 13 127 18
rect 20 12 132 13
rect -2 8 42 12
rect 46 10 98 12
rect 46 8 54 10
rect -2 6 54 8
rect 58 6 64 10
rect 68 6 74 10
rect 78 6 85 10
rect 89 8 98 10
rect 102 10 132 12
rect 102 8 112 10
rect 89 6 112 8
rect 116 6 120 10
rect 124 6 132 10
rect -2 -1 132 6
<< ntransistor >>
rect 11 15 13 29
rect 23 9 25 29
rect 35 9 37 29
rect 49 17 51 33
rect 59 17 61 33
rect 69 17 71 33
rect 81 17 83 29
rect 93 17 95 25
rect 105 17 107 25
rect 117 17 119 25
<< ptransistor >>
rect 11 55 13 79
rect 23 55 25 95
rect 35 55 37 95
rect 47 63 49 85
rect 59 63 61 85
rect 71 63 73 85
rect 83 61 85 85
rect 97 55 99 85
rect 107 55 109 85
rect 117 55 119 85
<< polycontact >>
rect 18 48 22 52
rect 38 38 42 42
rect 48 38 52 42
rect 58 38 62 42
rect 68 38 72 42
rect 78 38 82 42
rect 98 48 102 52
rect 108 48 112 52
rect 118 38 122 42
rect 18 32 22 36
<< ndcontact >>
rect 4 22 8 26
rect 16 22 20 26
rect 16 12 20 16
rect 28 18 32 22
rect 74 18 78 22
rect 86 18 90 22
rect 110 18 114 22
rect 122 18 126 22
rect 42 8 46 12
rect 98 8 102 12
<< pdcontact >>
rect 16 88 20 92
rect 4 68 8 72
rect 4 58 8 62
rect 16 78 20 82
rect 16 68 20 72
rect 16 58 20 62
rect 28 78 32 82
rect 28 68 32 72
rect 28 58 32 62
rect 64 88 68 92
rect 40 78 44 82
rect 52 78 56 82
rect 76 78 80 82
rect 88 68 92 72
rect 88 58 92 62
rect 122 78 126 82
<< psubstratepcontact >>
rect 54 6 58 10
rect 64 6 68 10
rect 74 6 78 10
rect 85 6 89 10
rect 112 6 116 10
rect 120 6 124 10
<< nsubstratencontact >>
rect 4 92 8 96
rect 76 92 80 96
rect 88 92 92 96
rect 100 92 104 96
rect 112 92 116 96
<< psubstratepdiff >>
rect 53 10 90 11
rect 53 6 54 10
rect 58 6 64 10
rect 68 6 74 10
rect 78 6 85 10
rect 89 6 90 10
rect 111 10 125 11
rect 53 5 90 6
rect 111 6 112 10
rect 116 6 120 10
rect 124 6 125 10
rect 111 5 125 6
<< nsubstratendiff >>
rect 3 96 9 97
rect 3 92 4 96
rect 8 92 9 96
rect 75 96 117 97
rect 3 85 9 92
rect 75 92 76 96
rect 80 92 88 96
rect 92 92 100 96
rect 104 92 112 96
rect 116 92 117 96
rect 75 91 117 92
<< labels >>
rlabel metal1 30 50 30 50 6 nq
rlabel metal1 30 50 30 50 6 nq
rlabel metal1 65 6 65 6 6 vss
rlabel metal1 65 6 65 6 6 vss
rlabel metal1 50 50 50 50 6 i0
rlabel metal1 50 50 50 50 6 i0
rlabel metal1 60 50 60 50 6 i1
rlabel metal1 70 55 70 55 6 i2
rlabel metal1 70 55 70 55 6 i2
rlabel metal1 60 50 60 50 6 i1
rlabel metal1 65 94 65 94 6 vdd
rlabel metal1 65 94 65 94 6 vdd
rlabel metal1 80 55 80 55 6 i6
rlabel metal1 80 55 80 55 6 i6
rlabel polycontact 100 50 100 50 6 i3
rlabel polycontact 100 50 100 50 6 i3
rlabel metal1 120 50 120 50 6 i5
rlabel polycontact 110 50 110 50 6 i4
rlabel metal1 120 50 120 50 6 i5
rlabel polycontact 110 50 110 50 6 i4
<< end >>
