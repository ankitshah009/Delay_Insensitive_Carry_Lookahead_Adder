.subckt xnr2v0x1 a b vdd vss z
*   SPICE3 file   created from xnr2v0x1.ext -      technology: scmos
m00 vdd    b      bn     vdd p w=18u  l=2.3636u ad=119.531p pd=38.25u   as=116p     ps=50u
m01 an     a      vdd    vdd p w=18u  l=2.3636u ad=72p      pd=26u      as=119.531p ps=38.25u
m02 z      b      an     vdd p w=18u  l=2.3636u ad=75.913p  pd=28.1739u as=72p      ps=26u
m03 w1     bn     z      vdd p w=28u  l=2.3636u ad=70p      pd=33u      as=118.087p ps=43.8261u
m04 vdd    an     w1     vdd p w=28u  l=2.3636u ad=185.938p pd=59.5u    as=70p      ps=33u
m05 vss    b      bn     vss n w=9u   l=2.3636u ad=36p      pd=17u      as=57p      ps=32u
m06 an     a      vss    vss n w=9u   l=2.3636u ad=36p      pd=17u      as=36p      ps=17u
m07 z      bn     an     vss n w=9u   l=2.3636u ad=36p      pd=17u      as=36p      ps=17u
m08 bn     an     z      vss n w=9u   l=2.3636u ad=57p      pd=32u      as=36p      ps=17u
C0  vss    vdd    0.003f
C1  an     bn     0.181f
C2  z      a      0.016f
C3  an     b      0.135f
C4  bn     a      0.086f
C5  z      vdd    0.132f
C6  a      b      0.160f
C7  bn     vdd    0.021f
C8  vss    z      0.099f
C9  b      vdd    0.086f
C10 vss    bn     0.192f
C11 z      bn     0.182f
C12 vss    b      0.016f
C13 w1     vdd    0.005f
C14 an     a      0.147f
C15 z      b      0.023f
C16 bn     b      0.186f
C17 an     vdd    0.048f
C18 a      vdd    0.014f
C19 w1     z      0.010f
C20 vss    an     0.069f
C21 vss    a      0.062f
C22 z      an     0.350f
C24 z      vss    0.019f
C25 an     vss    0.031f
C26 bn     vss    0.072f
C27 a      vss    0.024f
C28 b      vss    0.039f
.ends
