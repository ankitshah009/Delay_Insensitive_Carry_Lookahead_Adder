.subckt cgi2bv0x1 a b c vdd vss z
*   SPICE3 file   created from cgi2bv0x1.ext -      technology: scmos
m00 vdd    a      n1     vdd p w=27u  l=2.3636u ad=108p     pd=35u      as=125.667p ps=46u
m01 w1     a      vdd    vdd p w=27u  l=2.3636u ad=67.5p    pd=32u      as=108p     ps=35u
m02 z      bn     w1     vdd p w=27u  l=2.3636u ad=108p     pd=35u      as=67.5p    ps=32u
m03 n1     c      z      vdd p w=27u  l=2.3636u ad=125.667p pd=46u      as=108p     ps=35u
m04 vdd    bn     n1     vdd p w=27u  l=2.3636u ad=108p     pd=35u      as=125.667p ps=46u
m05 bn     b      vdd    vdd p w=27u  l=2.3636u ad=161p     pd=68u      as=108p     ps=35u
m06 vss    a      n3     vss n w=12u  l=2.3636u ad=73.5p    pd=27u      as=56p      ps=26u
m07 w2     a      vss    vss n w=12u  l=2.3636u ad=30p      pd=17u      as=73.5p    ps=27u
m08 z      bn     w2     vss n w=12u  l=2.3636u ad=48p      pd=20u      as=30p      ps=17u
m09 n3     c      z      vss n w=12u  l=2.3636u ad=56p      pd=26u      as=48p      ps=20u
m10 vss    bn     n3     vss n w=12u  l=2.3636u ad=73.5p    pd=27u      as=56p      ps=26u
m11 bn     b      vss    vss n w=12u  l=2.3636u ad=72p      pd=38u      as=73.5p    ps=27u
C0  bn     a      0.119f
C1  c      vdd    0.018f
C2  n3     c      0.097f
C3  z      n1     0.191f
C4  vss    b      0.019f
C5  a      vdd    0.022f
C6  z      c      0.116f
C7  vss    bn     0.125f
C8  n3     a      0.041f
C9  w2     n3     0.006f
C10 n1     c      0.025f
C11 vss    vdd    0.004f
C12 z      a      0.098f
C13 n3     vss    0.337f
C14 w2     z      0.008f
C15 w1     vdd    0.004f
C16 b      bn     0.403f
C17 n1     a      0.042f
C18 vss    z      0.068f
C19 c      a      0.043f
C20 b      vdd    0.024f
C21 z      w1     0.007f
C22 vss    n1     0.018f
C23 bn     vdd    0.152f
C24 w1     n1     0.023f
C25 vss    c      0.024f
C26 n3     bn     0.005f
C27 z      b      0.014f
C28 z      bn     0.065f
C29 n3     vdd    0.005f
C30 vss    a      0.020f
C31 z      vdd    0.062f
C32 b      c      0.035f
C33 n1     bn     0.017f
C34 n3     z      0.177f
C35 b      a      0.015f
C36 c      bn     0.239f
C37 n1     vdd    0.403f
C38 n3     n1     0.038f
C39 n3     vss    0.003f
C41 z      vss    0.003f
C42 b      vss    0.021f
C43 c      vss    0.021f
C44 bn     vss    0.041f
C45 a      vss    0.042f
.ends
