magic
tech scmos
timestamp 1180639975
<< checkpaint >>
rect -24 -26 114 126
<< ab >>
rect 0 0 90 100
<< pwell >>
rect -4 -6 94 49
<< nwell >>
rect -4 49 94 106
<< polysilicon >>
rect 11 93 13 98
rect 41 93 43 98
rect 53 93 55 98
rect 65 93 67 98
rect 77 93 79 98
rect 11 52 13 55
rect 11 51 32 52
rect 11 50 27 51
rect 25 47 27 50
rect 31 47 32 51
rect 25 46 32 47
rect 25 36 27 46
rect 41 43 43 55
rect 53 52 55 55
rect 65 52 67 55
rect 53 49 57 52
rect 65 51 73 52
rect 65 49 68 51
rect 55 43 57 49
rect 67 47 68 49
rect 72 47 73 51
rect 67 46 73 47
rect 41 42 51 43
rect 41 41 46 42
rect 45 38 46 41
rect 50 38 51 42
rect 45 37 51 38
rect 55 42 63 43
rect 55 38 58 42
rect 62 38 63 42
rect 55 37 63 38
rect 47 34 49 37
rect 55 34 57 37
rect 67 34 69 46
rect 77 43 79 55
rect 77 42 83 43
rect 77 40 78 42
rect 75 38 78 40
rect 82 38 83 42
rect 75 37 83 38
rect 75 34 77 37
rect 25 12 27 17
rect 47 12 49 17
rect 55 12 57 17
rect 67 12 69 17
rect 75 12 77 17
<< ndiffusion >>
rect 17 35 25 36
rect 17 31 18 35
rect 22 31 25 35
rect 17 27 25 31
rect 17 23 18 27
rect 22 23 25 27
rect 17 22 25 23
rect 20 17 25 22
rect 27 34 41 36
rect 27 32 47 34
rect 27 28 30 32
rect 34 28 47 32
rect 27 22 47 28
rect 27 18 30 22
rect 34 18 47 22
rect 27 17 47 18
rect 49 17 55 34
rect 57 22 67 34
rect 57 18 60 22
rect 64 18 67 22
rect 57 17 67 18
rect 69 17 75 34
rect 77 22 86 34
rect 77 18 80 22
rect 84 18 86 22
rect 77 17 86 18
<< pdiffusion >>
rect 3 92 11 93
rect 3 88 4 92
rect 8 88 11 92
rect 3 82 11 88
rect 3 78 4 82
rect 8 78 11 82
rect 3 72 11 78
rect 3 68 4 72
rect 8 68 11 72
rect 3 55 11 68
rect 13 71 18 93
rect 36 83 41 93
rect 33 82 41 83
rect 33 78 34 82
rect 38 78 41 82
rect 33 77 41 78
rect 13 70 21 71
rect 13 66 16 70
rect 20 66 21 70
rect 13 62 21 66
rect 13 58 16 62
rect 20 58 21 62
rect 13 57 21 58
rect 13 55 18 57
rect 36 55 41 77
rect 43 72 53 93
rect 43 68 46 72
rect 50 68 53 72
rect 43 55 53 68
rect 55 82 65 93
rect 55 78 58 82
rect 62 78 65 82
rect 55 55 65 78
rect 67 92 77 93
rect 67 88 70 92
rect 74 88 77 92
rect 67 55 77 88
rect 79 82 84 93
rect 79 81 87 82
rect 79 77 82 81
rect 86 77 87 81
rect 79 73 87 77
rect 79 69 82 73
rect 86 69 87 73
rect 79 68 87 69
rect 79 55 84 68
<< metal1 >>
rect -2 92 92 100
rect -2 88 4 92
rect 8 88 70 92
rect 74 88 92 92
rect 4 82 8 88
rect 33 78 34 82
rect 38 78 58 82
rect 62 81 86 82
rect 62 78 82 81
rect 4 72 8 78
rect 82 73 86 77
rect 4 67 8 68
rect 16 70 22 73
rect 20 66 22 70
rect 16 62 22 66
rect 7 58 16 62
rect 20 58 22 62
rect 18 35 22 58
rect 38 68 46 72
rect 50 68 51 72
rect 38 51 42 68
rect 58 62 62 73
rect 47 58 62 62
rect 26 47 27 51
rect 31 47 42 51
rect 18 27 22 31
rect 18 17 22 23
rect 30 32 34 33
rect 30 22 34 28
rect 38 22 42 47
rect 48 43 52 53
rect 46 42 52 43
rect 50 38 52 42
rect 46 37 52 38
rect 58 42 62 58
rect 58 37 62 38
rect 68 62 72 73
rect 82 68 86 69
rect 68 58 83 62
rect 68 51 72 58
rect 68 37 72 47
rect 78 42 82 53
rect 48 32 52 37
rect 78 32 82 38
rect 48 27 63 32
rect 67 27 82 32
rect 80 22 84 23
rect 38 18 60 22
rect 64 18 65 22
rect 30 12 34 18
rect 80 12 84 18
rect -2 0 92 12
<< ntransistor >>
rect 25 17 27 36
rect 47 17 49 34
rect 55 17 57 34
rect 67 17 69 34
rect 75 17 77 34
<< ptransistor >>
rect 11 55 13 93
rect 41 55 43 93
rect 53 55 55 93
rect 65 55 67 93
rect 77 55 79 93
<< polycontact >>
rect 27 47 31 51
rect 68 47 72 51
rect 46 38 50 42
rect 58 38 62 42
rect 78 38 82 42
<< ndcontact >>
rect 18 31 22 35
rect 18 23 22 27
rect 30 28 34 32
rect 30 18 34 22
rect 60 18 64 22
rect 80 18 84 22
<< pdcontact >>
rect 4 88 8 92
rect 4 78 8 82
rect 4 68 8 72
rect 34 78 38 82
rect 16 66 20 70
rect 16 58 20 62
rect 46 68 50 72
rect 58 78 62 82
rect 70 88 74 92
rect 82 77 86 81
rect 82 69 86 73
<< psubstratepcontact >>
rect 8 4 12 8
rect 18 4 22 8
<< nsubstratencontact >>
rect 25 92 29 96
<< psubstratepdiff >>
rect 7 8 23 9
rect 7 4 8 8
rect 12 4 18 8
rect 22 4 23 8
rect 7 3 23 4
<< nsubstratendiff >>
rect 24 96 30 97
rect 24 92 25 96
rect 29 92 30 96
rect 24 91 30 92
<< labels >>
rlabel polycontact 28 49 28 49 6 zn
rlabel metal1 10 60 10 60 6 z
rlabel metal1 10 60 10 60 6 z
rlabel metal1 20 45 20 45 6 z
rlabel metal1 20 45 20 45 6 z
rlabel metal1 45 6 45 6 6 vss
rlabel metal1 45 6 45 6 6 vss
rlabel metal1 50 40 50 40 6 b1
rlabel metal1 50 40 50 40 6 b1
rlabel metal1 34 49 34 49 6 zn
rlabel metal1 50 60 50 60 6 b2
rlabel metal1 50 60 50 60 6 b2
rlabel metal1 44 70 44 70 6 zn
rlabel metal1 45 94 45 94 6 vdd
rlabel metal1 45 94 45 94 6 vdd
rlabel metal1 51 20 51 20 6 zn
rlabel metal1 70 30 70 30 6 a1
rlabel metal1 60 30 60 30 6 b1
rlabel metal1 60 30 60 30 6 b1
rlabel metal1 70 30 70 30 6 a1
rlabel metal1 60 55 60 55 6 b2
rlabel metal1 70 55 70 55 6 a2
rlabel metal1 70 55 70 55 6 a2
rlabel metal1 60 55 60 55 6 b2
rlabel polycontact 80 40 80 40 6 a1
rlabel polycontact 80 40 80 40 6 a1
rlabel metal1 80 60 80 60 6 a2
rlabel metal1 80 60 80 60 6 a2
rlabel metal1 84 75 84 75 6 n3
rlabel pdcontact 59 80 59 80 6 n3
<< end >>
