magic
tech scmos
timestamp 1179385135
<< checkpaint >>
rect -22 -25 86 105
<< ab >>
rect 0 0 64 80
<< pwell >>
rect -4 -7 68 36
<< nwell >>
rect -4 36 68 87
<< polysilicon >>
rect 20 65 22 70
rect 30 65 32 70
rect 42 65 44 70
rect 52 65 54 70
rect 9 61 11 65
rect 9 39 11 43
rect 20 39 22 52
rect 30 49 32 52
rect 30 48 37 49
rect 30 44 32 48
rect 36 44 37 48
rect 30 43 37 44
rect 42 47 44 52
rect 42 46 48 47
rect 9 38 15 39
rect 9 34 10 38
rect 14 34 15 38
rect 9 33 15 34
rect 20 38 26 39
rect 20 34 21 38
rect 25 34 26 38
rect 20 33 26 34
rect 9 28 11 33
rect 24 28 26 33
rect 31 28 33 43
rect 42 42 43 46
rect 47 42 48 46
rect 42 41 48 42
rect 42 39 44 41
rect 38 37 44 39
rect 52 39 54 52
rect 52 38 58 39
rect 38 28 40 37
rect 52 34 53 38
rect 57 34 58 38
rect 52 33 58 34
rect 45 31 58 33
rect 45 28 47 31
rect 9 15 11 19
rect 24 7 26 12
rect 31 7 33 12
rect 38 7 40 12
rect 45 7 47 12
<< ndiffusion >>
rect 4 25 9 28
rect 2 24 9 25
rect 2 20 3 24
rect 7 20 9 24
rect 2 19 9 20
rect 11 19 24 28
rect 13 12 24 19
rect 26 12 31 28
rect 33 12 38 28
rect 40 12 45 28
rect 47 22 52 28
rect 47 21 54 22
rect 47 17 49 21
rect 53 17 54 21
rect 47 16 54 17
rect 47 12 52 16
rect 13 8 15 12
rect 19 8 22 12
rect 13 7 22 8
<< pdiffusion >>
rect 34 72 40 73
rect 34 68 35 72
rect 39 68 40 72
rect 34 65 40 68
rect 13 63 20 65
rect 13 61 14 63
rect 4 56 9 61
rect 2 55 9 56
rect 2 51 3 55
rect 7 51 9 55
rect 2 48 9 51
rect 2 44 3 48
rect 7 44 9 48
rect 2 43 9 44
rect 11 59 14 61
rect 18 59 20 63
rect 11 52 20 59
rect 22 63 30 65
rect 22 59 24 63
rect 28 59 30 63
rect 22 52 30 59
rect 32 52 42 65
rect 44 63 52 65
rect 44 59 46 63
rect 50 59 52 63
rect 44 52 52 59
rect 54 64 61 65
rect 54 60 56 64
rect 60 60 61 64
rect 54 57 61 60
rect 54 53 56 57
rect 60 53 61 57
rect 54 52 61 53
rect 11 43 18 52
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect -2 72 66 78
rect -2 68 35 72
rect 39 68 66 72
rect 14 63 18 68
rect 56 64 60 68
rect 2 55 7 63
rect 14 58 18 59
rect 22 59 24 63
rect 28 59 46 63
rect 50 59 51 63
rect 2 51 3 55
rect 22 54 26 59
rect 56 57 60 60
rect 2 48 7 51
rect 2 44 3 48
rect 2 43 7 44
rect 12 50 26 54
rect 2 25 6 43
rect 12 39 16 50
rect 34 48 38 55
rect 25 44 32 46
rect 36 44 38 48
rect 25 42 38 44
rect 42 46 46 55
rect 56 52 60 53
rect 42 42 43 46
rect 47 42 55 46
rect 10 38 16 39
rect 14 34 16 38
rect 20 34 21 38
rect 25 34 31 38
rect 41 34 53 38
rect 57 34 62 38
rect 10 33 16 34
rect 12 30 16 33
rect 27 30 31 34
rect 12 26 23 30
rect 27 26 47 30
rect 2 24 7 25
rect 2 20 3 24
rect 7 20 15 22
rect 2 17 15 20
rect 19 21 23 26
rect 19 17 49 21
rect 53 17 54 21
rect 58 17 62 34
rect -2 8 15 12
rect 19 8 66 12
rect -2 2 66 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
<< ntransistor >>
rect 9 19 11 28
rect 24 12 26 28
rect 31 12 33 28
rect 38 12 40 28
rect 45 12 47 28
<< ptransistor >>
rect 9 43 11 61
rect 20 52 22 65
rect 30 52 32 65
rect 42 52 44 65
rect 52 52 54 65
<< polycontact >>
rect 32 44 36 48
rect 10 34 14 38
rect 21 34 25 38
rect 43 42 47 46
rect 53 34 57 38
<< ndcontact >>
rect 3 20 7 24
rect 49 17 53 21
rect 15 8 19 12
<< pdcontact >>
rect 35 68 39 72
rect 3 51 7 55
rect 3 44 7 48
rect 14 59 18 63
rect 24 59 28 63
rect 46 59 50 63
rect 56 60 60 64
rect 56 53 60 57
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
<< psubstratepdiff >>
rect 0 2 64 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 64 2
rect 0 -3 64 -2
<< nsubstratendiff >>
rect 0 82 64 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 64 82
rect 0 77 64 78
<< labels >>
rlabel polycontact 12 36 12 36 6 zn
rlabel metal1 4 40 4 40 6 z
rlabel metal1 12 20 12 20 6 z
rlabel metal1 14 40 14 40 6 zn
rlabel metal1 32 6 32 6 6 vss
rlabel metal1 36 28 36 28 6 a
rlabel metal1 28 36 28 36 6 a
rlabel metal1 28 44 28 44 6 b
rlabel metal1 36 52 36 52 6 b
rlabel metal1 32 74 32 74 6 vdd
rlabel metal1 44 28 44 28 6 a
rlabel metal1 44 36 44 36 6 d
rlabel metal1 44 52 44 52 6 c
rlabel metal1 36 61 36 61 6 zn
rlabel metal1 36 19 36 19 6 zn
rlabel metal1 60 24 60 24 6 d
rlabel metal1 52 36 52 36 6 d
rlabel metal1 52 44 52 44 6 c
<< end >>
