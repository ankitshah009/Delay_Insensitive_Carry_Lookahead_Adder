magic
tech scmos
timestamp 1179386880
<< checkpaint >>
rect -22 -22 86 94
<< ab >>
rect 0 0 64 72
<< pwell >>
rect -4 -4 68 32
<< nwell >>
rect -4 32 68 76
<< polysilicon >>
rect 11 66 13 70
rect 18 66 20 70
rect 25 66 27 70
rect 35 66 37 70
rect 42 66 44 70
rect 49 66 51 70
rect 11 27 13 38
rect 18 35 20 38
rect 25 35 27 38
rect 35 35 37 38
rect 18 32 21 35
rect 25 33 37 35
rect 19 27 21 32
rect 35 27 37 33
rect 9 26 15 27
rect 9 22 10 26
rect 14 22 15 26
rect 9 21 15 22
rect 19 26 25 27
rect 19 22 20 26
rect 24 22 25 26
rect 19 21 25 22
rect 31 26 37 27
rect 31 22 32 26
rect 36 22 37 26
rect 42 29 44 38
rect 49 35 51 38
rect 49 34 58 35
rect 49 33 53 34
rect 52 30 53 33
rect 57 30 58 34
rect 52 29 58 30
rect 42 28 48 29
rect 42 24 43 28
rect 47 24 48 28
rect 42 23 48 24
rect 31 21 37 22
rect 9 18 11 21
rect 21 18 23 21
rect 31 18 33 21
rect 9 3 11 8
rect 21 3 23 8
rect 31 3 33 8
<< ndiffusion >>
rect 2 17 9 18
rect 2 13 3 17
rect 7 13 9 17
rect 2 12 9 13
rect 4 8 9 12
rect 11 8 21 18
rect 23 17 31 18
rect 23 13 25 17
rect 29 13 31 17
rect 23 8 31 13
rect 33 8 42 18
rect 13 4 14 8
rect 18 4 19 8
rect 13 3 19 4
rect 35 4 36 8
rect 40 4 42 8
rect 35 3 42 4
<< pdiffusion >>
rect 4 65 11 66
rect 4 61 5 65
rect 9 61 11 65
rect 4 58 11 61
rect 4 54 5 58
rect 9 54 11 58
rect 4 38 11 54
rect 13 38 18 66
rect 20 38 25 66
rect 27 58 35 66
rect 27 54 29 58
rect 33 54 35 58
rect 27 51 35 54
rect 27 47 29 51
rect 33 47 35 51
rect 27 38 35 47
rect 37 38 42 66
rect 44 38 49 66
rect 51 65 58 66
rect 51 61 53 65
rect 57 61 58 65
rect 51 58 58 61
rect 51 54 53 58
rect 57 54 58 58
rect 51 38 58 54
<< metal1 >>
rect -2 65 66 72
rect -2 64 5 65
rect 4 61 5 64
rect 9 64 53 65
rect 9 61 10 64
rect 4 58 10 61
rect 52 61 53 64
rect 57 64 66 65
rect 57 61 58 64
rect 4 54 5 58
rect 9 54 10 58
rect 29 58 33 59
rect 52 58 58 61
rect 52 54 53 58
rect 57 54 58 58
rect 29 51 33 54
rect 2 47 29 50
rect 33 47 39 50
rect 2 46 39 47
rect 2 17 6 46
rect 10 38 55 42
rect 10 26 14 38
rect 51 34 55 38
rect 10 21 14 22
rect 18 30 47 34
rect 51 30 53 34
rect 57 30 58 34
rect 18 26 24 30
rect 43 28 47 30
rect 18 22 20 26
rect 31 22 32 26
rect 36 22 39 26
rect 47 24 55 26
rect 43 22 55 24
rect 18 21 24 22
rect 34 18 39 22
rect 2 13 3 17
rect 7 13 25 17
rect 29 13 30 17
rect 34 13 47 18
rect -2 4 14 8
rect 18 4 36 8
rect 40 4 52 8
rect 56 4 66 8
rect -2 0 66 4
<< ntransistor >>
rect 9 8 11 18
rect 21 8 23 18
rect 31 8 33 18
<< ptransistor >>
rect 11 38 13 66
rect 18 38 20 66
rect 25 38 27 66
rect 35 38 37 66
rect 42 38 44 66
rect 49 38 51 66
<< polycontact >>
rect 10 22 14 26
rect 20 22 24 26
rect 32 22 36 26
rect 53 30 57 34
rect 43 24 47 28
<< ndcontact >>
rect 3 13 7 17
rect 25 13 29 17
rect 14 4 18 8
rect 36 4 40 8
<< pdcontact >>
rect 5 61 9 65
rect 5 54 9 58
rect 29 54 33 58
rect 29 47 33 51
rect 53 61 57 65
rect 53 54 57 58
<< psubstratepcontact >>
rect 52 4 56 8
<< psubstratepdiff >>
rect 51 8 57 24
rect 51 4 52 8
rect 56 4 57 8
rect 51 3 57 4
<< labels >>
rlabel metal1 4 28 4 28 6 z
rlabel metal1 20 24 20 24 6 b
rlabel metal1 12 28 12 28 6 a
rlabel metal1 20 40 20 40 6 a
rlabel metal1 12 48 12 48 6 z
rlabel metal1 20 48 20 48 6 z
rlabel metal1 32 4 32 4 6 vss
rlabel metal1 36 20 36 20 6 c
rlabel metal1 36 32 36 32 6 b
rlabel metal1 28 32 28 32 6 b
rlabel metal1 28 40 28 40 6 a
rlabel metal1 36 40 36 40 6 a
rlabel metal1 28 48 28 48 6 z
rlabel metal1 36 48 36 48 6 z
rlabel metal1 32 68 32 68 6 vdd
rlabel metal1 44 16 44 16 6 c
rlabel metal1 44 32 44 32 6 b
rlabel metal1 44 40 44 40 6 a
rlabel metal1 52 24 52 24 6 b
rlabel metal1 52 40 52 40 6 a
<< end >>
