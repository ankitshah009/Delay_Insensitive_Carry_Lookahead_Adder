magic
tech scmos
timestamp 1179386058
<< checkpaint >>
rect -22 -25 46 105
<< ab >>
rect 0 0 24 80
<< pwell >>
rect -4 -7 28 36
<< nwell >>
rect -4 36 28 87
<< polysilicon >>
rect 13 60 15 65
rect 13 39 15 45
rect 9 38 15 39
rect 9 34 10 38
rect 14 34 15 38
rect 9 33 15 34
rect 9 29 11 33
rect 9 17 11 22
<< ndiffusion >>
rect 2 28 9 29
rect 2 24 3 28
rect 7 24 9 28
rect 2 22 9 24
rect 11 22 19 29
rect 13 18 14 22
rect 18 18 19 22
rect 13 17 19 18
<< pdiffusion >>
rect 5 62 11 63
rect 5 58 6 62
rect 10 60 11 62
rect 10 58 13 60
rect 5 45 13 58
rect 15 55 20 60
rect 15 54 22 55
rect 15 50 17 54
rect 21 50 22 54
rect 15 49 22 50
rect 15 45 20 49
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect -2 68 26 78
rect 5 62 11 68
rect 5 58 6 62
rect 10 58 11 62
rect 2 50 17 54
rect 21 50 22 54
rect 2 29 6 50
rect 10 38 22 39
rect 14 34 22 38
rect 10 33 22 34
rect 2 28 7 29
rect 2 24 3 28
rect 18 25 22 33
rect 2 23 7 24
rect 13 18 14 22
rect 18 18 19 22
rect 13 12 19 18
rect -2 2 26 12
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
<< ntransistor >>
rect 9 22 11 29
<< ptransistor >>
rect 13 45 15 60
<< polycontact >>
rect 10 34 14 38
<< ndcontact >>
rect 3 24 7 28
rect 14 18 18 22
<< pdcontact >>
rect 6 58 10 62
rect 17 50 21 54
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
<< psubstratepdiff >>
rect 0 2 24 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 24 2
rect 0 -3 24 -2
<< nsubstratendiff >>
rect 0 82 24 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 24 82
rect 0 77 24 78
<< labels >>
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 6 12 6 6 vss
rlabel polycontact 12 36 12 36 6 a
rlabel metal1 12 52 12 52 6 z
rlabel metal1 12 74 12 74 6 vdd
rlabel metal1 20 32 20 32 6 a
<< end >>
