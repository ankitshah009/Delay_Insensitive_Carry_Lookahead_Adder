.subckt bf1v1x2 a vdd vss z
*   SPICE3 file   created from bf1v1x2.ext -      technology: scmos
m00 vdd    an     z      vdd p w=28u  l=2.3636u ad=160.533p pd=47.2889u as=166p     ps=70u
m01 an     a      vdd    vdd p w=17u  l=2.3636u ad=97p      pd=48u      as=97.4667p ps=28.7111u
m02 vss    an     z      vss n w=19u  l=2.3636u ad=110.2p   pd=36.7333u as=121p     ps=52u
m03 an     a      vss    vss n w=11u  l=2.3636u ad=67p      pd=36u      as=63.8p    ps=21.2667u
C0  vss    a      0.017f
C1  vss    an     0.104f
C2  a      z      0.027f
C3  z      an     0.287f
C4  a      vdd    0.014f
C5  an     vdd    0.091f
C6  vss    z      0.053f
C7  a      an     0.262f
C8  z      vdd    0.096f
C10 a      vss    0.021f
C11 z      vss    0.008f
C12 an     vss    0.016f
.ends
