magic
tech scmos
timestamp 1179386514
<< checkpaint >>
rect -22 -25 70 105
<< ab >>
rect 0 0 48 80
<< pwell >>
rect -4 -7 52 36
<< nwell >>
rect -4 36 52 87
<< polysilicon >>
rect 30 67 32 72
rect 37 67 39 72
rect 9 60 11 65
rect 19 60 21 65
rect 9 49 11 52
rect 9 48 15 49
rect 9 44 10 48
rect 14 44 15 48
rect 9 43 15 44
rect 9 30 11 43
rect 19 39 21 52
rect 30 49 32 52
rect 25 48 32 49
rect 25 44 26 48
rect 30 44 32 48
rect 25 43 32 44
rect 16 38 23 39
rect 16 34 18 38
rect 22 34 23 38
rect 16 33 23 34
rect 16 30 18 33
rect 27 30 29 43
rect 37 39 39 52
rect 37 38 46 39
rect 37 34 41 38
rect 45 34 46 38
rect 37 33 46 34
rect 37 30 39 33
rect 9 18 11 23
rect 16 18 18 23
rect 27 19 29 24
rect 37 19 39 24
<< ndiffusion >>
rect 2 28 9 30
rect 2 24 3 28
rect 7 24 9 28
rect 2 23 9 24
rect 11 23 16 30
rect 18 29 27 30
rect 18 25 20 29
rect 24 25 27 29
rect 18 24 27 25
rect 29 29 37 30
rect 29 25 31 29
rect 35 25 37 29
rect 29 24 37 25
rect 39 24 46 30
rect 18 23 25 24
rect 41 13 46 24
rect 40 12 46 13
rect 40 8 41 12
rect 45 8 46 12
rect 40 7 46 8
<< pdiffusion >>
rect 2 72 8 73
rect 2 68 3 72
rect 7 68 8 72
rect 2 67 8 68
rect 2 60 7 67
rect 23 62 30 67
rect 23 60 24 62
rect 2 52 9 60
rect 11 57 19 60
rect 11 53 13 57
rect 17 53 19 57
rect 11 52 19 53
rect 21 58 24 60
rect 28 58 30 62
rect 21 52 30 58
rect 32 52 37 67
rect 39 58 44 67
rect 39 57 46 58
rect 39 53 41 57
rect 45 53 46 57
rect 39 52 46 53
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect -2 72 50 78
rect -2 68 3 72
rect 7 68 50 72
rect 23 62 29 68
rect 23 58 24 62
rect 28 58 29 62
rect 2 53 13 57
rect 17 53 18 57
rect 34 55 38 63
rect 2 28 6 53
rect 26 49 38 55
rect 41 57 45 58
rect 10 48 14 49
rect 26 48 30 49
rect 14 44 22 47
rect 10 41 22 44
rect 41 46 45 53
rect 26 41 30 44
rect 34 42 45 46
rect 10 33 14 41
rect 34 38 38 42
rect 17 34 18 38
rect 22 34 38 38
rect 41 38 46 39
rect 45 34 46 38
rect 20 29 24 30
rect 2 24 3 28
rect 7 24 14 28
rect 10 17 14 24
rect 30 29 36 34
rect 41 33 46 34
rect 30 25 31 29
rect 35 25 36 29
rect 20 12 24 25
rect 42 22 46 33
rect 33 17 46 22
rect -2 8 41 12
rect 45 8 50 12
rect -2 2 50 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
<< ntransistor >>
rect 9 23 11 30
rect 16 23 18 30
rect 27 24 29 30
rect 37 24 39 30
<< ptransistor >>
rect 9 52 11 60
rect 19 52 21 60
rect 30 52 32 67
rect 37 52 39 67
<< polycontact >>
rect 10 44 14 48
rect 26 44 30 48
rect 18 34 22 38
rect 41 34 45 38
<< ndcontact >>
rect 3 24 7 28
rect 20 25 24 29
rect 31 25 35 29
rect 41 8 45 12
<< pdcontact >>
rect 3 68 7 72
rect 13 53 17 57
rect 24 58 28 62
rect 41 53 45 57
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
<< psubstratepdiff >>
rect 0 2 48 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 48 2
rect 0 -3 48 -2
<< nsubstratendiff >>
rect 0 82 48 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 48 82
rect 0 77 48 78
<< labels >>
rlabel polysilicon 20 49 20 49 6 nd
rlabel metal1 4 40 4 40 6 z
rlabel metal1 12 20 12 20 6 z
rlabel metal1 20 44 20 44 6 c
rlabel metal1 12 40 12 40 6 c
rlabel metal1 24 6 24 6 6 vss
rlabel metal1 33 31 33 31 6 nd
rlabel metal1 28 48 28 48 6 a
rlabel metal1 24 74 24 74 6 vdd
rlabel metal1 36 20 36 20 6 b
rlabel metal1 27 36 27 36 6 nd
rlabel metal1 44 28 44 28 6 b
rlabel metal1 43 50 43 50 6 nd
rlabel metal1 36 56 36 56 6 a
<< end >>
