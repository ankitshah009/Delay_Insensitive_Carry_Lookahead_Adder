magic
tech scmos
timestamp 1179384997
<< checkpaint >>
rect -22 -25 102 105
<< ab >>
rect 0 0 80 80
<< pwell >>
rect -4 -7 84 36
<< nwell >>
rect -4 36 84 87
<< polysilicon >>
rect 9 69 11 74
rect 19 69 21 74
rect 29 69 31 74
rect 39 58 41 63
rect 49 58 51 63
rect 59 58 61 63
rect 69 58 71 63
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 39 39 41 42
rect 49 39 51 42
rect 59 39 61 42
rect 9 38 32 39
rect 9 37 26 38
rect 20 34 26 37
rect 30 34 32 38
rect 20 33 32 34
rect 39 38 45 39
rect 39 34 40 38
rect 44 34 45 38
rect 39 33 45 34
rect 49 38 61 39
rect 49 34 56 38
rect 60 34 61 38
rect 69 37 71 42
rect 49 33 61 34
rect 20 30 22 33
rect 30 30 32 33
rect 42 30 44 33
rect 49 30 51 33
rect 59 30 61 33
rect 66 35 71 37
rect 66 30 68 35
rect 20 6 22 10
rect 30 6 32 10
rect 42 8 44 17
rect 49 12 51 17
rect 59 12 61 17
rect 66 8 68 17
rect 42 6 68 8
<< ndiffusion >>
rect 13 22 20 30
rect 13 18 14 22
rect 18 18 20 22
rect 13 15 20 18
rect 13 11 14 15
rect 18 11 20 15
rect 13 10 20 11
rect 22 29 30 30
rect 22 25 24 29
rect 28 25 30 29
rect 22 22 30 25
rect 22 18 24 22
rect 28 18 30 22
rect 22 10 30 18
rect 32 17 42 30
rect 44 17 49 30
rect 51 22 59 30
rect 51 18 53 22
rect 57 18 59 22
rect 51 17 59 18
rect 61 17 66 30
rect 68 29 75 30
rect 68 25 70 29
rect 74 25 75 29
rect 68 22 75 25
rect 68 18 70 22
rect 74 18 75 22
rect 68 17 75 18
rect 32 15 39 17
rect 32 11 34 15
rect 38 11 39 15
rect 32 10 39 11
<< pdiffusion >>
rect 4 55 9 69
rect 2 54 9 55
rect 2 50 3 54
rect 7 50 9 54
rect 2 47 9 50
rect 2 43 3 47
rect 7 43 9 47
rect 2 42 9 43
rect 11 68 19 69
rect 11 64 13 68
rect 17 64 19 68
rect 11 61 19 64
rect 11 57 13 61
rect 17 57 19 61
rect 11 42 19 57
rect 21 54 29 69
rect 21 50 23 54
rect 27 50 29 54
rect 21 47 29 50
rect 21 43 23 47
rect 27 43 29 47
rect 21 42 29 43
rect 31 58 37 69
rect 31 57 39 58
rect 31 53 33 57
rect 37 53 39 57
rect 31 42 39 53
rect 41 54 49 58
rect 41 50 43 54
rect 47 50 49 54
rect 41 47 49 50
rect 41 43 43 47
rect 47 43 49 47
rect 41 42 49 43
rect 51 57 59 58
rect 51 53 53 57
rect 57 53 59 57
rect 51 42 59 53
rect 61 55 69 58
rect 61 51 63 55
rect 67 51 69 55
rect 61 48 69 51
rect 61 44 63 48
rect 67 44 69 48
rect 61 42 69 44
rect 71 57 78 58
rect 71 53 73 57
rect 77 53 78 57
rect 71 42 78 53
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect -2 68 82 78
rect 13 61 17 64
rect 13 56 17 57
rect 33 57 37 68
rect 2 54 7 55
rect 2 50 3 54
rect 2 47 7 50
rect 2 43 3 47
rect 23 54 27 55
rect 53 57 57 68
rect 33 52 37 53
rect 43 54 47 55
rect 23 47 27 50
rect 73 57 77 68
rect 53 52 57 53
rect 63 55 67 56
rect 43 47 47 50
rect 73 52 77 53
rect 63 48 67 51
rect 7 43 23 46
rect 2 42 27 43
rect 31 43 43 47
rect 47 44 63 47
rect 47 43 67 44
rect 9 30 14 42
rect 31 38 35 43
rect 74 38 78 47
rect 25 34 26 38
rect 30 34 35 38
rect 39 34 40 38
rect 44 34 47 38
rect 55 34 56 38
rect 60 34 78 38
rect 9 29 28 30
rect 9 26 24 29
rect 24 22 28 25
rect 13 18 14 22
rect 18 18 19 22
rect 13 15 19 18
rect 31 22 35 34
rect 41 30 47 34
rect 41 26 55 30
rect 70 29 74 30
rect 70 22 74 25
rect 31 18 53 22
rect 57 18 58 22
rect 24 17 28 18
rect 13 12 14 15
rect -2 11 14 12
rect 18 12 19 15
rect 33 12 34 15
rect 18 11 34 12
rect 38 12 39 15
rect 70 12 74 18
rect 38 11 82 12
rect -2 2 82 11
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
<< ntransistor >>
rect 20 10 22 30
rect 30 10 32 30
rect 42 17 44 30
rect 49 17 51 30
rect 59 17 61 30
rect 66 17 68 30
<< ptransistor >>
rect 9 42 11 69
rect 19 42 21 69
rect 29 42 31 69
rect 39 42 41 58
rect 49 42 51 58
rect 59 42 61 58
rect 69 42 71 58
<< polycontact >>
rect 26 34 30 38
rect 40 34 44 38
rect 56 34 60 38
<< ndcontact >>
rect 14 18 18 22
rect 14 11 18 15
rect 24 25 28 29
rect 24 18 28 22
rect 53 18 57 22
rect 70 25 74 29
rect 70 18 74 22
rect 34 11 38 15
<< pdcontact >>
rect 3 50 7 54
rect 3 43 7 47
rect 13 64 17 68
rect 13 57 17 61
rect 23 50 27 54
rect 23 43 27 47
rect 33 53 37 57
rect 43 50 47 54
rect 43 43 47 47
rect 53 53 57 57
rect 63 51 67 55
rect 63 44 67 48
rect 73 53 77 57
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
<< psubstratepdiff >>
rect 0 2 80 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 80 2
rect 0 -3 80 -2
<< nsubstratendiff >>
rect 0 82 80 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 80 82
rect 0 77 80 78
<< labels >>
rlabel polysilicon 26 36 26 36 6 zn
rlabel pdcontact 4 52 4 52 6 z
rlabel metal1 20 28 20 28 6 z
rlabel metal1 12 36 12 36 6 z
rlabel metal1 20 44 20 44 6 z
rlabel metal1 40 6 40 6 6 vss
rlabel metal1 44 32 44 32 6 a
rlabel metal1 30 36 30 36 6 zn
rlabel metal1 45 49 45 49 6 zn
rlabel metal1 40 74 40 74 6 vdd
rlabel metal1 52 28 52 28 6 a
rlabel metal1 44 20 44 20 6 zn
rlabel metal1 60 36 60 36 6 b
rlabel metal1 68 36 68 36 6 b
rlabel metal1 49 45 49 45 6 zn
rlabel metal1 76 44 76 44 6 b
rlabel metal1 65 49 65 49 6 zn
<< end >>
