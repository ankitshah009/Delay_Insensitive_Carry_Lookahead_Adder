magic
tech scmos
timestamp 1179386727
<< checkpaint >>
rect -22 -25 54 105
<< ab >>
rect 0 0 32 80
<< pwell >>
rect -4 -7 36 36
<< nwell >>
rect -4 36 36 87
<< polysilicon >>
rect 12 70 14 74
rect 19 70 21 74
rect 12 47 14 50
rect 9 46 15 47
rect 9 42 10 46
rect 14 42 15 46
rect 9 41 15 42
rect 10 29 12 41
rect 19 38 21 50
rect 19 37 25 38
rect 19 33 20 37
rect 24 33 25 37
rect 19 32 25 33
rect 20 29 22 32
rect 10 18 12 23
rect 20 18 22 23
<< ndiffusion >>
rect 2 28 10 29
rect 2 24 3 28
rect 7 24 10 28
rect 2 23 10 24
rect 12 28 20 29
rect 12 24 14 28
rect 18 24 20 28
rect 12 23 20 24
rect 22 28 30 29
rect 22 24 25 28
rect 29 24 30 28
rect 22 23 30 24
<< pdiffusion >>
rect 7 64 12 70
rect 5 63 12 64
rect 5 59 6 63
rect 10 59 12 63
rect 5 58 12 59
rect 7 50 12 58
rect 14 50 19 70
rect 21 69 30 70
rect 21 65 25 69
rect 29 65 30 69
rect 21 62 30 65
rect 21 58 25 62
rect 29 58 30 62
rect 21 50 30 58
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect -2 69 34 78
rect -2 68 25 69
rect 29 68 34 69
rect 2 37 6 63
rect 10 59 11 63
rect 25 62 29 65
rect 25 57 29 58
rect 18 50 22 55
rect 10 46 22 50
rect 10 41 14 42
rect 26 39 30 47
rect 18 37 30 39
rect 2 33 14 37
rect 18 33 20 37
rect 24 33 30 37
rect 3 28 7 29
rect 10 24 14 33
rect 25 28 29 29
rect 18 24 19 28
rect 3 12 7 24
rect 25 12 29 24
rect -2 2 34 12
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
<< ntransistor >>
rect 10 23 12 29
rect 20 23 22 29
<< ptransistor >>
rect 12 50 14 70
rect 19 50 21 70
<< polycontact >>
rect 10 42 14 46
rect 20 33 24 37
<< ndcontact >>
rect 3 24 7 28
rect 14 24 18 28
rect 25 24 29 28
<< pdcontact >>
rect 6 59 10 63
rect 25 65 29 69
rect 25 58 29 62
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
<< psubstratepdiff >>
rect 0 2 32 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 32 2
rect 0 -3 32 -2
<< nsubstratendiff >>
rect 0 82 32 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 32 82
rect 0 77 32 78
<< labels >>
rlabel metal1 4 48 4 48 6 z
rlabel metal1 12 28 12 28 6 z
rlabel polycontact 12 44 12 44 6 b
rlabel metal1 16 6 16 6 6 vss
rlabel metal1 20 36 20 36 6 a
rlabel metal1 20 52 20 52 6 b
rlabel metal1 16 74 16 74 6 vdd
rlabel metal1 28 40 28 40 6 a
<< end >>
