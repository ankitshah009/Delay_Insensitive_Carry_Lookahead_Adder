magic
tech scmos
timestamp 1185094803
<< checkpaint >>
rect -22 -22 72 122
<< ab >>
rect 0 0 50 100
<< pwell >>
rect -4 -4 54 48
<< nwell >>
rect -4 48 54 104
<< polysilicon >>
rect 27 83 29 88
rect 35 83 37 88
rect 15 76 17 81
rect 15 53 17 56
rect 13 52 23 53
rect 13 48 18 52
rect 22 48 23 52
rect 13 47 23 48
rect 13 34 15 47
rect 27 43 29 56
rect 35 53 37 56
rect 35 52 43 53
rect 35 50 38 52
rect 37 48 38 50
rect 42 48 43 52
rect 37 47 43 48
rect 27 42 33 43
rect 27 40 28 42
rect 25 38 28 40
rect 32 38 33 42
rect 25 37 33 38
rect 25 34 27 37
rect 37 34 39 47
rect 13 19 15 24
rect 25 22 27 27
rect 37 22 39 27
<< ndiffusion >>
rect 5 33 13 34
rect 5 29 6 33
rect 10 29 13 33
rect 5 28 13 29
rect 8 24 13 28
rect 15 27 25 34
rect 27 32 37 34
rect 27 28 30 32
rect 34 28 37 32
rect 27 27 37 28
rect 39 32 47 34
rect 39 28 42 32
rect 46 28 47 32
rect 39 27 47 28
rect 15 24 23 27
rect 17 12 23 24
rect 17 8 18 12
rect 22 8 23 12
rect 17 7 23 8
<< pdiffusion >>
rect 19 82 27 83
rect 19 78 20 82
rect 24 78 27 82
rect 19 76 27 78
rect 10 70 15 76
rect 7 69 15 70
rect 7 65 8 69
rect 12 65 15 69
rect 7 61 15 65
rect 7 57 8 61
rect 12 57 15 61
rect 7 56 15 57
rect 17 56 27 76
rect 29 56 35 83
rect 37 82 45 83
rect 37 78 40 82
rect 44 78 45 82
rect 37 74 45 78
rect 37 70 40 74
rect 44 70 45 74
rect 37 69 45 70
rect 37 56 42 69
<< metal1 >>
rect -2 96 52 100
rect -2 92 32 96
rect 36 92 42 96
rect 46 92 52 96
rect -2 88 52 92
rect 20 82 24 88
rect 20 77 24 78
rect 40 82 44 83
rect 40 74 44 78
rect 8 69 12 73
rect 8 61 12 65
rect 8 34 12 57
rect 6 33 12 34
rect 10 29 12 33
rect 6 28 12 29
rect 18 70 40 72
rect 18 68 44 70
rect 18 52 22 68
rect 27 58 42 63
rect 18 32 22 48
rect 28 42 32 53
rect 38 52 42 58
rect 38 47 42 48
rect 32 38 43 42
rect 28 37 43 38
rect 42 32 46 33
rect 18 28 30 32
rect 34 28 35 32
rect 8 22 12 28
rect 8 17 23 22
rect 42 12 46 28
rect -2 8 18 12
rect 22 8 52 12
rect -2 4 32 8
rect 36 4 42 8
rect 46 4 52 8
rect -2 0 52 4
<< ntransistor >>
rect 13 24 15 34
rect 25 27 27 34
rect 37 27 39 34
<< ptransistor >>
rect 15 56 17 76
rect 27 56 29 83
rect 35 56 37 83
<< polycontact >>
rect 18 48 22 52
rect 38 48 42 52
rect 28 38 32 42
<< ndcontact >>
rect 6 29 10 33
rect 30 28 34 32
rect 42 28 46 32
rect 18 8 22 12
<< pdcontact >>
rect 20 78 24 82
rect 8 65 12 69
rect 8 57 12 61
rect 40 78 44 82
rect 40 70 44 74
<< psubstratepcontact >>
rect 32 4 36 8
rect 42 4 46 8
<< nsubstratencontact >>
rect 32 92 36 96
rect 42 92 46 96
<< psubstratepdiff >>
rect 31 8 47 9
rect 31 4 32 8
rect 36 4 42 8
rect 46 4 47 8
rect 31 3 47 4
<< nsubstratendiff >>
rect 31 96 47 97
rect 31 92 32 96
rect 36 92 42 96
rect 46 92 47 96
rect 31 91 47 92
<< labels >>
rlabel metal1 20 20 20 20 6 z
rlabel metal1 10 45 10 45 6 z
rlabel polycontact 20 50 20 50 6 zn
rlabel metal1 25 6 25 6 6 vss
rlabel metal1 26 30 26 30 6 zn
rlabel metal1 30 45 30 45 6 a
rlabel metal1 30 60 30 60 6 b
rlabel metal1 25 94 25 94 6 vdd
rlabel metal1 40 40 40 40 6 a
rlabel metal1 40 55 40 55 6 b
rlabel metal1 42 75 42 75 6 zn
<< end >>
