.subckt nd2v5x05 a b vdd vss z
*   SPICE3 file   created from nd2v5x05.ext -      technology: scmos
m00 z      b      vdd    vdd p w=12u  l=2.3636u ad=48p      pd=20u      as=147p     ps=57u
m01 vdd    a      z      vdd p w=12u  l=2.3636u ad=147p     pd=57u      as=48p      ps=20u
m02 w1     b      z      vss n w=8u   l=2.3636u ad=20p      pd=13u      as=52p      ps=30u
m03 vss    a      w1     vss n w=8u   l=2.3636u ad=107p     pd=44u      as=20p      ps=13u
C0  z      a      0.052f
C1  vss    vdd    0.006f
C2  a      b      0.081f
C3  z      vdd    0.037f
C4  b      vdd    0.139f
C5  vss    z      0.026f
C6  vss    b      0.007f
C7  z      b      0.073f
C8  a      vdd    0.019f
C9  vss    a      0.092f
C11 z      vss    0.006f
C12 a      vss    0.020f
C13 b      vss    0.022f
.ends
