.subckt mxi2v2x2 a0 a1 s vdd vss z
*   SPICE3 file   created from mxi2v2x2.ext -      technology: scmos
m00 a0n    s      z      vdd p w=20u  l=2.3636u ad=80p      pd=28u      as=106p     ps=42.5u
m01 vdd    a0     a0n    vdd p w=20u  l=2.3636u ad=90p      pd=32.9167u as=80p      ps=28u
m02 a0n    a0     vdd    vdd p w=20u  l=2.3636u ad=80p      pd=28u      as=90p      ps=32.9167u
m03 z      s      a0n    vdd p w=20u  l=2.3636u ad=106p     pd=42.5u    as=80p      ps=28u
m04 a1n    sn     z      vdd p w=20u  l=2.3636u ad=95p      pd=29.5u    as=106p     ps=42.5u
m05 vdd    a1     a1n    vdd p w=20u  l=2.3636u ad=90p      pd=32.9167u as=95p      ps=29.5u
m06 a1n    a1     vdd    vdd p w=20u  l=2.3636u ad=95p      pd=29.5u    as=90p      ps=32.9167u
m07 z      sn     a1n    vdd p w=20u  l=2.3636u ad=106p     pd=42.5u    as=95p      ps=29.5u
m08 vdd    s      sn     vdd p w=16u  l=2.3636u ad=72p      pd=26.3333u as=92p      ps=46u
m09 a0n    a0     vss    vss n w=20u  l=2.3636u ad=100p     pd=30u      as=197.2p   ps=68u
m10 z      sn     a0n    vss n w=20u  l=2.3636u ad=119p     pd=54u      as=100p     ps=30u
m11 a1n    a1     vss    vss n w=20u  l=2.3636u ad=80p      pd=28u      as=197.2p   ps=68u
m12 z      s      a1n    vss n w=20u  l=2.3636u ad=119p     pd=54u      as=80p      ps=28u
m13 vss    s      sn     vss n w=10u  l=2.3636u ad=98.6p    pd=34u      as=62p      ps=34u
C0  a0n    vdd    0.063f
C1  z      s      0.067f
C2  a1     a0     0.025f
C3  vss    a1n    0.050f
C4  a1     vdd    0.020f
C5  sn     s      0.243f
C6  vss    z      0.311f
C7  a1n    a0n    0.021f
C8  a0     vdd    0.004f
C9  a0n    z      0.529f
C10 a1n    a1     0.162f
C11 vss    sn     0.065f
C12 a0n    sn     0.039f
C13 z      a1     0.152f
C14 vss    s      0.103f
C15 a1     sn     0.166f
C16 a1n    vdd    0.074f
C17 z      a0     0.060f
C18 a1     s      0.080f
C19 z      vdd    0.244f
C20 sn     a0     0.034f
C21 vss    a0n    0.112f
C22 sn     vdd    0.274f
C23 a0     s      0.083f
C24 a1n    z      0.348f
C25 vss    a1     0.039f
C26 s      vdd    0.052f
C27 vss    a0     0.122f
C28 a0n    a1     0.021f
C29 a1n    sn     0.423f
C30 z      sn     0.682f
C31 a0n    a0     0.124f
C32 a1n    s      0.023f
C33 vss    vdd    0.005f
C35 a1n    vss    0.005f
C36 a0n    vss    0.005f
C37 z      vss    0.017f
C38 a1     vss    0.029f
C39 sn     vss    0.041f
C40 a0     vss    0.043f
C41 s      vss    0.098f
.ends
