magic
tech scmos
timestamp 1182081810
<< checkpaint >>
rect -25 -26 121 114
<< ab >>
rect 0 0 96 88
<< pwell >>
rect -7 -8 103 40
<< nwell >>
rect -7 40 103 96
<< polysilicon >>
rect 5 80 14 86
rect 18 80 27 86
rect 37 80 46 86
rect 50 80 59 86
rect 69 85 78 86
rect 69 81 73 85
rect 77 81 78 85
rect 69 80 78 81
rect 82 85 91 86
rect 82 81 83 85
rect 87 81 91 85
rect 82 80 91 81
rect 9 77 11 80
rect 21 77 23 80
rect 41 77 43 80
rect 53 77 55 80
rect 73 77 75 80
rect 85 77 87 80
rect 9 48 11 51
rect 21 48 23 51
rect 41 48 43 51
rect 53 48 55 51
rect 73 48 75 51
rect 85 48 87 51
rect 2 47 11 48
rect 2 43 6 47
rect 10 43 11 47
rect 2 42 11 43
rect 15 47 30 48
rect 15 43 22 47
rect 26 43 30 47
rect 15 42 30 43
rect 34 47 43 48
rect 34 43 38 47
rect 42 43 43 47
rect 34 42 43 43
rect 47 47 62 48
rect 47 43 48 47
rect 52 43 62 47
rect 47 42 62 43
rect 66 47 75 48
rect 66 43 70 47
rect 74 43 75 47
rect 66 42 75 43
rect 79 42 94 48
rect 2 32 17 38
rect 21 32 30 38
rect 34 37 49 38
rect 34 33 35 37
rect 39 33 49 37
rect 34 32 49 33
rect 53 37 62 38
rect 53 33 54 37
rect 58 33 62 37
rect 53 32 62 33
rect 66 37 81 38
rect 66 33 70 37
rect 74 33 81 37
rect 66 32 81 33
rect 85 32 94 38
rect 9 29 11 32
rect 21 29 23 32
rect 41 29 43 32
rect 53 29 55 32
rect 73 29 75 32
rect 85 29 87 32
rect 9 8 11 11
rect 21 8 23 11
rect 41 8 43 11
rect 53 8 55 11
rect 73 8 75 11
rect 85 8 87 11
rect 5 7 14 8
rect 5 3 6 7
rect 10 3 14 7
rect 5 2 14 3
rect 18 7 27 8
rect 18 3 22 7
rect 26 3 27 7
rect 18 2 27 3
rect 37 2 46 8
rect 50 2 59 8
rect 69 2 78 8
rect 82 7 91 8
rect 82 3 83 7
rect 87 3 91 7
rect 82 2 91 3
<< ndiffusion >>
rect 2 11 9 29
rect 11 11 21 29
rect 23 11 30 29
rect 34 25 41 29
rect 34 21 35 25
rect 39 21 41 25
rect 34 18 41 21
rect 34 14 35 18
rect 39 14 41 18
rect 34 11 41 14
rect 43 17 53 29
rect 43 13 46 17
rect 50 13 53 17
rect 43 11 53 13
rect 55 26 62 29
rect 55 22 57 26
rect 61 22 62 26
rect 55 19 62 22
rect 55 15 57 19
rect 61 15 62 19
rect 55 11 62 15
rect 66 26 73 29
rect 66 22 67 26
rect 71 22 73 26
rect 66 19 73 22
rect 66 15 67 19
rect 71 15 73 19
rect 66 11 73 15
rect 75 17 85 29
rect 75 13 78 17
rect 82 13 85 17
rect 75 11 85 13
rect 87 11 94 29
<< pdiffusion >>
rect 2 75 9 77
rect 2 71 3 75
rect 7 71 9 75
rect 2 68 9 71
rect 2 64 3 68
rect 7 64 9 68
rect 2 51 9 64
rect 11 66 21 77
rect 11 62 14 66
rect 18 62 21 66
rect 11 59 21 62
rect 11 55 14 59
rect 18 55 21 59
rect 11 51 21 55
rect 23 75 30 77
rect 23 71 25 75
rect 29 71 30 75
rect 23 68 30 71
rect 23 64 25 68
rect 29 64 30 68
rect 23 51 30 64
rect 34 66 41 77
rect 34 62 35 66
rect 39 62 41 66
rect 34 59 41 62
rect 34 55 35 59
rect 39 55 41 59
rect 34 51 41 55
rect 43 74 53 77
rect 43 70 46 74
rect 50 70 53 74
rect 43 67 53 70
rect 43 63 46 67
rect 50 63 53 67
rect 43 51 53 63
rect 55 66 62 77
rect 55 62 57 66
rect 61 62 62 66
rect 55 59 62 62
rect 55 55 57 59
rect 61 55 62 59
rect 55 51 62 55
rect 66 75 73 77
rect 66 71 67 75
rect 71 71 73 75
rect 66 68 73 71
rect 66 64 67 68
rect 71 64 73 68
rect 66 51 73 64
rect 75 66 85 77
rect 75 62 78 66
rect 82 62 85 66
rect 75 58 85 62
rect 75 54 78 58
rect 82 54 85 58
rect 75 51 85 54
rect 87 74 94 77
rect 87 70 89 74
rect 93 70 94 74
rect 87 67 94 70
rect 87 63 89 67
rect 93 63 94 67
rect 87 51 94 63
<< metal1 >>
rect -2 86 2 90
rect 30 86 34 90
rect 2 82 30 85
rect -2 81 34 82
rect 62 86 66 90
rect 94 86 98 90
rect 62 81 66 82
rect 72 81 73 85
rect 77 81 83 85
rect 87 81 88 85
rect 94 81 98 82
rect 3 75 7 81
rect 3 68 7 71
rect 25 75 29 81
rect 25 68 29 71
rect 3 63 7 64
rect 14 66 18 67
rect 46 74 67 75
rect 50 71 67 74
rect 71 74 93 75
rect 71 71 89 74
rect 46 67 50 70
rect 67 68 71 71
rect 25 63 29 64
rect 35 66 39 67
rect 14 59 18 62
rect 46 62 50 63
rect 57 66 61 67
rect 89 67 93 70
rect 67 63 71 64
rect 78 66 82 67
rect 35 59 39 62
rect 18 55 35 58
rect 57 59 61 62
rect 89 62 93 63
rect 39 55 57 58
rect 14 54 61 55
rect 6 50 10 51
rect 6 47 27 50
rect 46 47 50 51
rect 70 47 74 59
rect 10 46 22 47
rect 6 37 10 43
rect 21 43 22 46
rect 26 43 27 47
rect 37 43 38 47
rect 42 43 48 47
rect 52 43 59 47
rect 21 34 27 43
rect 35 37 39 38
rect 21 33 35 34
rect 21 30 39 33
rect 53 37 59 43
rect 53 33 54 37
rect 58 33 59 37
rect 53 30 59 33
rect 70 37 74 43
rect 70 32 74 33
rect 78 58 82 62
rect 78 26 82 54
rect 35 25 57 26
rect 39 22 57 25
rect 61 22 67 26
rect 71 22 82 26
rect 39 21 42 22
rect 35 18 42 21
rect 57 19 61 22
rect 39 14 42 18
rect 35 13 42 14
rect 46 17 50 18
rect 57 14 61 15
rect 67 19 71 22
rect 67 13 71 15
rect 78 17 82 18
rect 46 7 50 13
rect 78 7 82 13
rect -2 6 6 7
rect 2 3 6 6
rect 10 3 22 7
rect 26 6 83 7
rect 26 3 30 6
rect -2 -2 2 2
rect 34 3 62 6
rect 30 -2 34 2
rect 66 3 83 6
rect 87 6 98 7
rect 87 3 94 6
rect 62 -2 66 2
rect 94 -2 98 2
<< metal2 >>
rect -2 86 98 90
rect 2 82 30 86
rect 34 82 62 86
rect 66 82 94 86
rect -2 80 98 82
rect -2 6 98 8
rect 2 2 30 6
rect 34 2 62 6
rect 66 2 94 6
rect -2 -2 98 2
<< ntransistor >>
rect 9 11 11 29
rect 21 11 23 29
rect 41 11 43 29
rect 53 11 55 29
rect 73 11 75 29
rect 85 11 87 29
<< ptransistor >>
rect 9 51 11 77
rect 21 51 23 77
rect 41 51 43 77
rect 53 51 55 77
rect 73 51 75 77
rect 85 51 87 77
<< polycontact >>
rect 73 81 77 85
rect 83 81 87 85
rect 6 43 10 47
rect 22 43 26 47
rect 38 43 42 47
rect 48 43 52 47
rect 70 43 74 47
rect 35 33 39 37
rect 54 33 58 37
rect 70 33 74 37
rect 6 3 10 7
rect 22 3 26 7
rect 83 3 87 7
<< ndcontact >>
rect 35 21 39 25
rect 35 14 39 18
rect 46 13 50 17
rect 57 22 61 26
rect 57 15 61 19
rect 67 22 71 26
rect 67 15 71 19
rect 78 13 82 17
<< pdcontact >>
rect 3 71 7 75
rect 3 64 7 68
rect 14 62 18 66
rect 14 55 18 59
rect 25 71 29 75
rect 25 64 29 68
rect 35 62 39 66
rect 35 55 39 59
rect 46 70 50 74
rect 46 63 50 67
rect 57 62 61 66
rect 57 55 61 59
rect 67 71 71 75
rect 67 64 71 68
rect 78 62 82 66
rect 78 54 82 58
rect 89 70 93 74
rect 89 63 93 67
<< m2contact >>
rect -2 82 2 86
rect 30 82 34 86
rect 62 82 66 86
rect 94 82 98 86
rect -2 2 2 6
rect 30 2 34 6
rect 62 2 66 6
rect 94 2 98 6
<< psubstratepcontact >>
rect -2 2 2 6
rect 30 2 34 6
rect 62 2 66 6
rect 94 2 98 6
<< nsubstratencontact >>
rect -2 82 2 86
rect 30 82 34 86
rect 62 82 66 86
rect 94 82 98 86
<< psubstratepdiff >>
rect -3 6 3 7
rect -3 2 -2 6
rect 2 2 3 6
rect 29 6 35 7
rect 29 2 30 6
rect 34 2 35 6
rect 61 6 67 7
rect 61 2 62 6
rect 66 2 67 6
rect 93 6 99 7
rect 93 2 94 6
rect 98 2 99 6
rect -3 0 3 2
rect 29 0 35 2
rect 61 0 67 2
rect 93 0 99 2
<< nsubstratendiff >>
rect -3 86 3 88
rect 29 86 35 88
rect 61 86 67 88
rect 93 86 99 88
rect -3 82 -2 86
rect 2 82 3 86
rect -3 81 3 82
rect 29 82 30 86
rect 34 82 35 86
rect 29 81 35 82
rect 61 82 62 86
rect 66 82 67 86
rect 61 81 67 82
rect 93 82 94 86
rect 98 82 99 86
rect 93 81 99 82
<< labels >>
rlabel polycontact 8 44 8 44 6 a
rlabel metal1 32 32 32 32 6 a
rlabel metal1 16 48 16 48 6 a
rlabel metal1 24 40 24 40 6 a
rlabel metal1 40 20 40 20 6 z
rlabel metal1 56 24 56 24 6 z
rlabel metal1 48 24 48 24 6 z
rlabel polycontact 56 36 56 36 6 b
rlabel metal1 48 48 48 48 6 b
rlabel metal1 72 24 72 24 6 z
rlabel metal1 64 24 64 24 6 z
rlabel metal1 72 48 72 48 6 c
rlabel metal1 80 48 80 48 6 z
rlabel metal2 48 4 48 4 6 vss
rlabel metal2 48 84 48 84 6 vdd
<< end >>
