magic
tech scmos
timestamp 1179385678
<< checkpaint >>
rect -22 -22 222 94
<< ab >>
rect 0 0 200 72
<< pwell >>
rect -4 -4 204 32
<< nwell >>
rect -4 32 204 76
<< polysilicon >>
rect 21 66 23 70
rect 31 66 33 70
rect 41 66 43 70
rect 51 66 53 70
rect 61 66 63 70
rect 71 66 73 70
rect 81 66 83 70
rect 91 66 93 70
rect 101 66 103 70
rect 108 66 110 70
rect 121 66 123 70
rect 128 66 130 70
rect 138 66 140 70
rect 145 66 147 70
rect 157 66 159 70
rect 167 66 169 70
rect 177 66 179 70
rect 10 46 12 51
rect 10 35 12 38
rect 21 35 23 38
rect 31 35 33 38
rect 10 34 33 35
rect 10 30 11 34
rect 15 30 18 34
rect 22 33 33 34
rect 22 30 23 33
rect 10 29 23 30
rect 21 26 23 29
rect 31 26 33 33
rect 41 35 43 38
rect 51 35 53 38
rect 41 34 54 35
rect 41 30 42 34
rect 46 30 49 34
rect 53 31 54 34
rect 61 31 63 38
rect 53 30 63 31
rect 41 29 63 30
rect 41 26 43 29
rect 51 26 53 29
rect 61 26 63 29
rect 71 35 73 38
rect 81 35 83 38
rect 91 35 93 38
rect 101 35 103 38
rect 71 34 93 35
rect 71 30 72 34
rect 76 33 93 34
rect 76 30 83 33
rect 71 29 83 30
rect 71 26 73 29
rect 81 26 83 29
rect 91 26 93 33
rect 97 34 103 35
rect 97 30 98 34
rect 102 30 103 34
rect 97 29 103 30
rect 101 26 103 29
rect 108 35 110 38
rect 121 35 123 38
rect 108 34 123 35
rect 108 30 114 34
rect 118 30 123 34
rect 108 29 123 30
rect 108 26 110 29
rect 121 26 123 29
rect 128 35 130 38
rect 138 35 140 38
rect 128 34 140 35
rect 128 30 129 34
rect 133 30 140 34
rect 128 29 140 30
rect 128 26 130 29
rect 138 26 140 29
rect 145 35 147 38
rect 157 35 159 38
rect 167 35 169 38
rect 177 35 179 38
rect 145 34 179 35
rect 145 30 146 34
rect 150 33 179 34
rect 150 30 160 33
rect 145 29 160 30
rect 145 26 147 29
rect 158 26 160 29
rect 168 26 170 33
rect 21 5 23 10
rect 31 5 33 10
rect 41 7 43 12
rect 51 7 53 12
rect 61 4 63 12
rect 71 8 73 12
rect 81 8 83 12
rect 91 8 93 12
rect 101 4 103 12
rect 108 7 110 12
rect 61 2 103 4
rect 121 7 123 12
rect 128 7 130 12
rect 138 7 140 12
rect 145 7 147 12
rect 158 2 160 6
rect 168 2 170 6
<< ndiffusion >>
rect 14 24 21 26
rect 14 20 15 24
rect 19 20 21 24
rect 14 17 21 20
rect 14 13 15 17
rect 19 13 21 17
rect 14 10 21 13
rect 23 25 31 26
rect 23 21 25 25
rect 29 21 31 25
rect 23 18 31 21
rect 23 14 25 18
rect 29 14 31 18
rect 23 10 31 14
rect 33 24 41 26
rect 33 20 35 24
rect 39 20 41 24
rect 33 17 41 20
rect 33 13 35 17
rect 39 13 41 17
rect 33 12 41 13
rect 43 25 51 26
rect 43 21 45 25
rect 49 21 51 25
rect 43 18 51 21
rect 43 14 45 18
rect 49 14 51 18
rect 43 12 51 14
rect 53 17 61 26
rect 53 13 55 17
rect 59 13 61 17
rect 53 12 61 13
rect 63 25 71 26
rect 63 21 65 25
rect 69 21 71 25
rect 63 18 71 21
rect 63 14 65 18
rect 69 14 71 18
rect 63 12 71 14
rect 73 25 81 26
rect 73 21 75 25
rect 79 21 81 25
rect 73 12 81 21
rect 83 18 91 26
rect 83 14 85 18
rect 89 14 91 18
rect 83 12 91 14
rect 93 25 101 26
rect 93 21 95 25
rect 99 21 101 25
rect 93 12 101 21
rect 103 12 108 26
rect 110 12 121 26
rect 123 12 128 26
rect 130 25 138 26
rect 130 21 132 25
rect 136 21 138 25
rect 130 12 138 21
rect 140 12 145 26
rect 147 12 158 26
rect 33 10 39 12
rect 112 8 119 12
rect 112 4 113 8
rect 117 4 119 8
rect 149 11 158 12
rect 149 7 150 11
rect 154 7 158 11
rect 149 6 158 7
rect 160 25 168 26
rect 160 21 162 25
rect 166 21 168 25
rect 160 18 168 21
rect 160 14 162 18
rect 166 14 168 18
rect 160 6 168 14
rect 170 19 178 26
rect 170 15 172 19
rect 176 15 178 19
rect 170 11 178 15
rect 170 7 172 11
rect 176 7 178 11
rect 170 6 178 7
rect 112 3 119 4
<< pdiffusion >>
rect 14 65 21 66
rect 14 61 15 65
rect 19 61 21 65
rect 14 58 21 61
rect 14 54 15 58
rect 19 54 21 58
rect 14 51 21 54
rect 14 47 15 51
rect 19 47 21 51
rect 14 46 21 47
rect 5 44 10 46
rect 3 43 10 44
rect 3 39 4 43
rect 8 39 10 43
rect 3 38 10 39
rect 12 38 21 46
rect 23 50 31 66
rect 23 46 25 50
rect 29 46 31 50
rect 23 43 31 46
rect 23 39 25 43
rect 29 39 31 43
rect 23 38 31 39
rect 33 65 41 66
rect 33 61 35 65
rect 39 61 41 65
rect 33 58 41 61
rect 33 54 35 58
rect 39 54 41 58
rect 33 51 41 54
rect 33 47 35 51
rect 39 47 41 51
rect 33 38 41 47
rect 43 58 51 66
rect 43 54 45 58
rect 49 54 51 58
rect 43 51 51 54
rect 43 47 45 51
rect 49 47 51 51
rect 43 38 51 47
rect 53 65 61 66
rect 53 61 55 65
rect 59 61 61 65
rect 53 58 61 61
rect 53 54 55 58
rect 59 54 61 58
rect 53 38 61 54
rect 63 58 71 66
rect 63 54 65 58
rect 69 54 71 58
rect 63 51 71 54
rect 63 47 65 51
rect 69 47 71 51
rect 63 38 71 47
rect 73 50 81 66
rect 73 46 75 50
rect 79 46 81 50
rect 73 43 81 46
rect 73 39 75 43
rect 79 39 81 43
rect 73 38 81 39
rect 83 58 91 66
rect 83 54 85 58
rect 89 54 91 58
rect 83 51 91 54
rect 83 47 85 51
rect 89 47 91 51
rect 83 38 91 47
rect 93 50 101 66
rect 93 46 95 50
rect 99 46 101 50
rect 93 43 101 46
rect 93 39 95 43
rect 99 39 101 43
rect 93 38 101 39
rect 103 38 108 66
rect 110 65 121 66
rect 110 61 113 65
rect 117 61 121 65
rect 110 38 121 61
rect 123 38 128 66
rect 130 50 138 66
rect 130 46 132 50
rect 136 46 138 50
rect 130 38 138 46
rect 140 38 145 66
rect 147 65 157 66
rect 147 61 150 65
rect 154 61 157 65
rect 147 38 157 61
rect 159 58 167 66
rect 159 54 161 58
rect 165 54 167 58
rect 159 51 167 54
rect 159 47 161 51
rect 165 47 167 51
rect 159 38 167 47
rect 169 65 177 66
rect 169 61 171 65
rect 175 61 177 65
rect 169 58 177 61
rect 169 54 171 58
rect 175 54 177 58
rect 169 38 177 54
rect 179 51 184 66
rect 179 50 186 51
rect 179 46 181 50
rect 185 46 186 50
rect 179 43 186 46
rect 179 39 181 43
rect 185 39 186 43
rect 179 38 186 39
<< metal1 >>
rect -2 68 202 72
rect -2 64 4 68
rect 8 65 189 68
rect 8 64 15 65
rect 4 60 8 64
rect 4 55 8 56
rect 19 64 35 65
rect 15 58 19 61
rect 15 51 19 54
rect 39 64 55 65
rect 35 58 39 61
rect 59 64 113 65
rect 112 61 113 64
rect 117 64 150 65
rect 117 61 118 64
rect 149 61 150 64
rect 154 64 171 65
rect 154 61 155 64
rect 170 61 171 64
rect 175 64 189 65
rect 193 64 202 68
rect 175 61 176 64
rect 35 51 39 54
rect 15 46 19 47
rect 25 50 29 51
rect 35 46 39 47
rect 45 58 49 59
rect 45 51 49 54
rect 55 58 59 61
rect 170 58 176 61
rect 55 53 59 54
rect 64 54 65 58
rect 69 54 85 58
rect 89 54 161 58
rect 165 54 166 58
rect 170 54 171 58
rect 175 54 176 58
rect 189 60 193 64
rect 189 55 193 56
rect 64 51 69 54
rect 85 51 89 54
rect 64 50 65 51
rect 49 47 65 50
rect 45 46 69 47
rect 74 50 79 51
rect 74 46 75 50
rect 161 51 166 54
rect 85 46 89 47
rect 94 46 95 50
rect 99 46 132 50
rect 136 46 158 50
rect 165 50 166 51
rect 165 47 181 50
rect 161 46 181 47
rect 185 46 186 50
rect 25 43 29 46
rect 74 43 79 46
rect 94 43 99 46
rect 3 39 4 43
rect 8 39 25 43
rect 2 34 22 35
rect 2 30 11 34
rect 15 30 18 34
rect 2 29 22 30
rect 25 34 29 39
rect 66 35 70 43
rect 74 39 75 43
rect 79 39 95 43
rect 82 38 99 39
rect 113 38 150 42
rect 66 34 78 35
rect 25 30 42 34
rect 46 30 49 34
rect 53 30 54 34
rect 66 30 72 34
rect 76 30 78 34
rect 2 21 6 29
rect 25 25 29 30
rect 66 29 78 30
rect 45 25 69 26
rect 82 25 86 38
rect 113 34 119 38
rect 146 34 150 38
rect 97 30 98 34
rect 102 30 108 34
rect 113 30 114 34
rect 118 30 119 34
rect 123 30 129 34
rect 133 30 134 34
rect 104 26 108 30
rect 123 26 127 30
rect 146 29 150 30
rect 15 24 19 25
rect 15 17 19 20
rect 4 16 8 17
rect 4 8 8 12
rect 25 18 29 21
rect 25 13 29 14
rect 35 24 39 25
rect 35 17 39 20
rect 49 22 65 25
rect 45 18 49 21
rect 64 21 65 22
rect 74 21 75 25
rect 79 21 95 25
rect 99 21 100 25
rect 104 22 127 26
rect 154 25 158 46
rect 180 43 186 46
rect 180 39 181 43
rect 185 39 186 43
rect 131 21 132 25
rect 136 21 158 25
rect 162 25 167 26
rect 166 21 167 25
rect 64 18 69 21
rect 162 18 167 21
rect 45 13 49 14
rect 55 17 59 18
rect 64 14 65 18
rect 69 14 85 18
rect 89 14 162 18
rect 166 14 167 18
rect 172 19 176 20
rect 15 8 19 13
rect 35 8 39 13
rect 55 8 59 13
rect 172 11 176 15
rect 149 8 150 11
rect -2 4 4 8
rect 8 4 113 8
rect 117 7 150 8
rect 154 8 155 11
rect 154 7 172 8
rect 186 16 190 17
rect 186 8 190 12
rect 176 7 186 8
rect 117 4 186 7
rect 190 4 202 8
rect -2 0 202 4
<< ntransistor >>
rect 21 10 23 26
rect 31 10 33 26
rect 41 12 43 26
rect 51 12 53 26
rect 61 12 63 26
rect 71 12 73 26
rect 81 12 83 26
rect 91 12 93 26
rect 101 12 103 26
rect 108 12 110 26
rect 121 12 123 26
rect 128 12 130 26
rect 138 12 140 26
rect 145 12 147 26
rect 158 6 160 26
rect 168 6 170 26
<< ptransistor >>
rect 10 38 12 46
rect 21 38 23 66
rect 31 38 33 66
rect 41 38 43 66
rect 51 38 53 66
rect 61 38 63 66
rect 71 38 73 66
rect 81 38 83 66
rect 91 38 93 66
rect 101 38 103 66
rect 108 38 110 66
rect 121 38 123 66
rect 128 38 130 66
rect 138 38 140 66
rect 145 38 147 66
rect 157 38 159 66
rect 167 38 169 66
rect 177 38 179 66
<< polycontact >>
rect 11 30 15 34
rect 18 30 22 34
rect 42 30 46 34
rect 49 30 53 34
rect 72 30 76 34
rect 98 30 102 34
rect 114 30 118 34
rect 129 30 133 34
rect 146 30 150 34
<< ndcontact >>
rect 15 20 19 24
rect 15 13 19 17
rect 25 21 29 25
rect 25 14 29 18
rect 35 20 39 24
rect 35 13 39 17
rect 45 21 49 25
rect 45 14 49 18
rect 55 13 59 17
rect 65 21 69 25
rect 65 14 69 18
rect 75 21 79 25
rect 85 14 89 18
rect 95 21 99 25
rect 132 21 136 25
rect 113 4 117 8
rect 150 7 154 11
rect 162 21 166 25
rect 162 14 166 18
rect 172 15 176 19
rect 172 7 176 11
<< pdcontact >>
rect 15 61 19 65
rect 15 54 19 58
rect 15 47 19 51
rect 4 39 8 43
rect 25 46 29 50
rect 25 39 29 43
rect 35 61 39 65
rect 35 54 39 58
rect 35 47 39 51
rect 45 54 49 58
rect 45 47 49 51
rect 55 61 59 65
rect 55 54 59 58
rect 65 54 69 58
rect 65 47 69 51
rect 75 46 79 50
rect 75 39 79 43
rect 85 54 89 58
rect 85 47 89 51
rect 95 46 99 50
rect 95 39 99 43
rect 113 61 117 65
rect 132 46 136 50
rect 150 61 154 65
rect 161 54 165 58
rect 161 47 165 51
rect 171 61 175 65
rect 171 54 175 58
rect 181 46 185 50
rect 181 39 185 43
<< psubstratepcontact >>
rect 4 12 8 16
rect 4 4 8 8
rect 186 12 190 16
rect 186 4 190 8
<< nsubstratencontact >>
rect 4 64 8 68
rect 4 56 8 60
rect 189 64 193 68
rect 189 56 193 60
<< psubstratepdiff >>
rect 3 16 9 24
rect 3 12 4 16
rect 8 12 9 16
rect 3 8 9 12
rect 3 4 4 8
rect 8 4 9 8
rect 3 3 9 4
rect 185 16 191 24
rect 185 12 186 16
rect 190 12 191 16
rect 185 8 191 12
rect 185 4 186 8
rect 190 4 191 8
rect 185 3 191 4
<< nsubstratendiff >>
rect 3 68 9 69
rect 3 64 4 68
rect 8 64 9 68
rect 188 68 194 69
rect 3 60 9 64
rect 3 56 4 60
rect 8 56 9 60
rect 3 55 9 56
rect 188 64 189 68
rect 193 64 194 68
rect 188 60 194 64
rect 188 56 189 60
rect 193 56 194 60
rect 188 55 194 56
<< labels >>
rlabel polysilicon 47 32 47 32 6 bn
rlabel polycontact 100 32 100 32 6 bn
rlabel polysilicon 134 32 134 32 6 bn
rlabel polycontact 20 32 20 32 6 b
rlabel polycontact 12 32 12 32 6 b
rlabel metal1 4 28 4 28 6 b
rlabel metal1 16 41 16 41 6 bn
rlabel metal1 47 19 47 19 6 n3
rlabel metal1 66 20 66 20 6 n3
rlabel metal1 76 32 76 32 6 c
rlabel metal1 39 32 39 32 6 bn
rlabel metal1 68 36 68 36 6 c
rlabel pdcontact 76 48 76 48 6 z
rlabel metal1 66 52 66 52 6 n1
rlabel metal1 47 52 47 52 6 n1
rlabel metal1 100 4 100 4 6 vss
rlabel metal1 84 32 84 32 6 z
rlabel metal1 102 32 102 32 6 bn
rlabel metal1 92 40 92 40 6 z
rlabel metal1 116 36 116 36 6 a
rlabel metal1 108 48 108 48 6 z
rlabel metal1 100 48 100 48 6 z
rlabel metal1 116 48 116 48 6 z
rlabel metal1 87 52 87 52 6 n1
rlabel metal1 100 68 100 68 6 vdd
rlabel metal1 156 32 156 32 6 z
rlabel polycontact 148 32 148 32 6 a
rlabel metal1 128 32 128 32 6 bn
rlabel metal1 124 40 124 40 6 a
rlabel metal1 140 40 140 40 6 a
rlabel metal1 132 40 132 40 6 a
rlabel metal1 124 48 124 48 6 z
rlabel metal1 132 48 132 48 6 z
rlabel metal1 148 48 148 48 6 z
rlabel metal1 140 48 140 48 6 z
rlabel metal1 164 20 164 20 6 n3
rlabel metal1 115 16 115 16 6 n3
rlabel metal1 183 44 183 44 6 n1
rlabel metal1 163 52 163 52 6 n1
rlabel metal1 115 56 115 56 6 n1
<< end >>
