magic
tech scmos
timestamp 1185039022
<< checkpaint >>
rect -22 -24 142 124
<< ab >>
rect 0 0 120 100
<< pwell >>
rect -2 -4 122 49
<< nwell >>
rect -2 49 122 104
<< polysilicon >>
rect 27 95 29 98
rect 39 95 41 98
rect 51 95 53 98
rect 59 95 61 98
rect 71 95 73 98
rect 83 95 85 98
rect 91 95 93 98
rect 15 69 17 72
rect 15 53 17 55
rect 7 52 17 53
rect 7 48 8 52
rect 12 48 17 52
rect 7 47 17 48
rect 15 37 17 47
rect 27 53 29 75
rect 39 73 41 75
rect 33 72 41 73
rect 33 68 34 72
rect 38 68 41 72
rect 33 67 41 68
rect 27 52 33 53
rect 27 48 28 52
rect 32 48 33 52
rect 27 47 33 48
rect 15 26 17 29
rect 27 23 29 47
rect 39 41 41 67
rect 51 63 53 75
rect 47 62 53 63
rect 47 58 48 62
rect 52 58 53 62
rect 47 57 53 58
rect 47 52 53 53
rect 47 48 48 52
rect 52 51 53 52
rect 59 51 61 75
rect 71 73 73 75
rect 83 73 85 75
rect 52 49 61 51
rect 52 48 53 49
rect 47 47 53 48
rect 39 39 53 41
rect 33 32 41 33
rect 33 28 34 32
rect 38 28 41 32
rect 33 27 41 28
rect 39 23 41 27
rect 51 23 53 39
rect 59 23 61 49
rect 69 71 73 73
rect 79 71 85 73
rect 69 33 71 71
rect 79 53 81 71
rect 91 63 93 75
rect 103 69 105 72
rect 85 62 93 63
rect 85 58 86 62
rect 90 58 93 62
rect 85 57 93 58
rect 75 52 81 53
rect 75 48 76 52
rect 80 51 81 52
rect 103 51 105 55
rect 80 49 105 51
rect 80 48 81 49
rect 75 47 81 48
rect 79 39 81 47
rect 65 32 71 33
rect 65 28 66 32
rect 70 28 71 32
rect 65 27 71 28
rect 75 37 81 39
rect 85 42 93 43
rect 85 38 86 42
rect 90 38 93 42
rect 85 37 93 38
rect 103 37 105 49
rect 75 23 77 37
rect 81 32 87 33
rect 81 28 82 32
rect 86 28 87 32
rect 81 27 87 28
rect 71 21 77 23
rect 71 19 73 21
rect 83 19 85 27
rect 91 19 93 37
rect 103 26 105 29
rect 27 8 29 11
rect 39 8 41 11
rect 51 8 53 11
rect 59 8 61 11
rect 71 4 73 7
rect 83 4 85 7
rect 91 4 93 7
<< ndiffusion >>
rect 7 29 15 37
rect 17 34 25 37
rect 17 30 20 34
rect 24 30 25 34
rect 17 29 25 30
rect 7 22 13 29
rect 43 32 49 33
rect 43 28 44 32
rect 48 28 49 32
rect 43 23 49 28
rect 7 18 8 22
rect 12 18 13 22
rect 7 17 13 18
rect 19 22 27 23
rect 19 18 20 22
rect 24 18 27 22
rect 19 11 27 18
rect 29 11 39 23
rect 41 11 51 23
rect 53 11 59 23
rect 61 22 69 23
rect 61 18 64 22
rect 68 19 69 22
rect 95 34 103 37
rect 95 30 96 34
rect 100 30 103 34
rect 95 29 103 30
rect 105 29 113 37
rect 95 22 101 23
rect 95 19 96 22
rect 68 18 71 19
rect 61 11 71 18
rect 63 7 71 11
rect 73 12 83 19
rect 73 8 76 12
rect 80 8 83 12
rect 73 7 83 8
rect 85 7 91 19
rect 93 18 96 19
rect 100 18 101 22
rect 93 7 101 18
rect 107 12 113 29
rect 107 8 108 12
rect 112 8 113 12
rect 107 7 113 8
<< pdiffusion >>
rect 7 82 13 83
rect 7 78 8 82
rect 12 78 13 82
rect 7 69 13 78
rect 19 82 27 95
rect 19 78 20 82
rect 24 78 27 82
rect 19 75 27 78
rect 29 75 39 95
rect 41 75 51 95
rect 53 75 59 95
rect 61 82 71 95
rect 61 78 64 82
rect 68 78 71 82
rect 61 75 71 78
rect 73 92 83 95
rect 73 88 76 92
rect 80 88 83 92
rect 73 75 83 88
rect 85 75 91 95
rect 93 82 101 95
rect 93 78 96 82
rect 100 78 101 82
rect 93 75 101 78
rect 107 82 113 83
rect 107 78 108 82
rect 112 78 113 82
rect 7 55 15 69
rect 17 62 25 69
rect 17 58 20 62
rect 24 58 25 62
rect 17 55 25 58
rect 43 72 49 75
rect 43 68 44 72
rect 48 68 49 72
rect 43 67 49 68
rect 107 69 113 78
rect 95 62 103 69
rect 95 58 96 62
rect 100 58 103 62
rect 95 55 103 58
rect 105 55 113 69
<< metal1 >>
rect -2 92 122 101
rect -2 88 76 92
rect 80 88 122 92
rect -2 87 122 88
rect 7 82 13 87
rect 7 78 8 82
rect 12 78 13 82
rect 7 77 13 78
rect 19 82 69 83
rect 19 78 20 82
rect 24 78 64 82
rect 68 78 69 82
rect 19 77 69 78
rect 95 82 101 83
rect 95 78 96 82
rect 100 78 101 82
rect 95 73 101 78
rect 107 82 113 87
rect 107 78 108 82
rect 112 78 113 82
rect 107 77 113 78
rect 8 72 39 73
rect 7 68 34 72
rect 38 68 39 72
rect 7 67 39 68
rect 43 72 112 73
rect 43 68 44 72
rect 48 68 113 72
rect 43 67 113 68
rect 7 52 13 67
rect 18 62 53 63
rect 7 48 8 52
rect 12 48 13 52
rect 7 28 13 48
rect 17 58 20 62
rect 24 58 48 62
rect 52 58 53 62
rect 17 57 53 58
rect 17 35 23 57
rect 27 52 33 53
rect 27 48 28 52
rect 32 48 33 52
rect 27 40 33 48
rect 38 52 53 53
rect 38 48 48 52
rect 52 48 53 52
rect 38 47 53 48
rect 57 43 63 67
rect 78 62 91 63
rect 44 42 63 43
rect 43 38 63 42
rect 67 53 73 62
rect 78 58 86 62
rect 90 58 91 62
rect 78 57 91 58
rect 95 62 101 63
rect 95 58 96 62
rect 100 58 103 62
rect 95 57 103 58
rect 85 53 91 57
rect 67 52 81 53
rect 67 48 76 52
rect 80 48 81 52
rect 67 47 81 48
rect 85 47 92 53
rect 67 38 73 47
rect 85 43 91 47
rect 78 42 91 43
rect 78 38 86 42
rect 90 38 91 42
rect 43 37 62 38
rect 78 37 91 38
rect 17 34 25 35
rect 17 30 20 34
rect 24 33 25 34
rect 24 32 39 33
rect 24 30 34 32
rect 17 28 34 30
rect 38 28 39 32
rect 18 27 39 28
rect 43 32 49 37
rect 97 35 103 57
rect 95 34 103 35
rect 95 33 96 34
rect 43 28 44 32
rect 48 28 49 32
rect 43 27 49 28
rect 65 32 96 33
rect 65 28 66 32
rect 70 28 82 32
rect 86 30 96 32
rect 100 30 103 34
rect 86 28 103 30
rect 65 27 102 28
rect 107 23 113 67
rect 7 22 13 23
rect 7 18 8 22
rect 12 18 13 22
rect 7 13 13 18
rect 19 22 69 23
rect 19 18 20 22
rect 24 18 64 22
rect 68 18 69 22
rect 19 17 69 18
rect 95 22 113 23
rect 95 18 96 22
rect 100 18 113 22
rect 95 17 112 18
rect -2 12 122 13
rect -2 8 76 12
rect 80 8 108 12
rect 112 8 122 12
rect -2 -1 122 8
<< ntransistor >>
rect 15 29 17 37
rect 27 11 29 23
rect 39 11 41 23
rect 51 11 53 23
rect 59 11 61 23
rect 103 29 105 37
rect 71 7 73 19
rect 83 7 85 19
rect 91 7 93 19
<< ptransistor >>
rect 27 75 29 95
rect 39 75 41 95
rect 51 75 53 95
rect 59 75 61 95
rect 71 75 73 95
rect 83 75 85 95
rect 91 75 93 95
rect 15 55 17 69
rect 103 55 105 69
<< polycontact >>
rect 8 48 12 52
rect 34 68 38 72
rect 28 48 32 52
rect 48 58 52 62
rect 48 48 52 52
rect 34 28 38 32
rect 86 58 90 62
rect 76 48 80 52
rect 66 28 70 32
rect 86 38 90 42
rect 82 28 86 32
<< ndcontact >>
rect 20 30 24 34
rect 44 28 48 32
rect 8 18 12 22
rect 20 18 24 22
rect 64 18 68 22
rect 96 30 100 34
rect 76 8 80 12
rect 96 18 100 22
rect 108 8 112 12
<< pdcontact >>
rect 8 78 12 82
rect 20 78 24 82
rect 64 78 68 82
rect 76 88 80 92
rect 96 78 100 82
rect 108 78 112 82
rect 20 58 24 62
rect 44 68 48 72
rect 96 58 100 62
<< labels >>
rlabel polycontact 10 50 10 50 6 cmd1
rlabel polycontact 10 50 10 50 6 cmd1
rlabel polycontact 30 50 30 50 6 i2
rlabel polycontact 30 50 30 50 6 i2
rlabel metal1 60 6 60 6 6 vss
rlabel metal1 60 6 60 6 6 vss
rlabel polycontact 50 50 50 50 6 i1
rlabel polycontact 50 50 50 50 6 i1
rlabel metal1 70 50 70 50 6 cmd0
rlabel metal1 70 50 70 50 6 cmd0
rlabel metal1 60 94 60 94 6 vdd
rlabel metal1 60 94 60 94 6 vdd
rlabel metal1 80 40 80 40 6 i0
rlabel metal1 80 40 80 40 6 i0
rlabel metal1 90 50 90 50 6 i0
rlabel metal1 90 50 90 50 6 i0
rlabel metal1 80 60 80 60 6 i0
rlabel metal1 80 60 80 60 6 i0
rlabel metal1 110 45 110 45 6 nq
rlabel metal1 110 45 110 45 6 nq
<< end >>
