magic
tech scmos
timestamp 1179385042
<< checkpaint >>
rect -22 -25 78 105
<< ab >>
rect 0 0 56 80
<< pwell >>
rect -4 -7 60 36
<< nwell >>
rect -4 36 60 87
<< polysilicon >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 61 31 66
rect 39 61 41 65
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 46
rect 39 43 41 46
rect 39 42 47 43
rect 9 38 22 39
rect 9 34 17 38
rect 21 34 22 38
rect 9 33 22 34
rect 28 38 34 39
rect 28 34 29 38
rect 33 34 34 38
rect 28 33 34 34
rect 10 30 12 33
rect 20 30 22 33
rect 32 30 34 33
rect 39 38 42 42
rect 46 38 47 42
rect 39 37 47 38
rect 39 30 41 37
rect 10 11 12 16
rect 20 11 22 16
rect 32 13 34 18
rect 39 13 41 18
<< ndiffusion >>
rect 2 16 10 30
rect 12 22 20 30
rect 12 18 14 22
rect 18 18 20 22
rect 12 16 20 18
rect 22 18 32 30
rect 34 18 39 30
rect 41 24 46 30
rect 41 23 48 24
rect 41 19 43 23
rect 47 19 48 23
rect 41 18 48 19
rect 22 16 30 18
rect 2 12 8 16
rect 2 8 3 12
rect 7 8 8 12
rect 24 12 30 16
rect 2 7 8 8
rect 24 8 25 12
rect 29 8 30 12
rect 24 7 30 8
<< pdiffusion >>
rect 2 69 9 70
rect 2 65 3 69
rect 7 65 9 69
rect 2 62 9 65
rect 2 58 3 62
rect 7 58 9 62
rect 2 42 9 58
rect 11 62 19 70
rect 11 58 13 62
rect 17 58 19 62
rect 11 55 19 58
rect 11 51 13 55
rect 17 51 19 55
rect 11 42 19 51
rect 21 61 27 70
rect 21 60 29 61
rect 21 56 23 60
rect 27 56 29 60
rect 21 46 29 56
rect 31 60 39 61
rect 31 56 33 60
rect 37 56 39 60
rect 31 53 39 56
rect 31 49 33 53
rect 37 49 39 53
rect 31 46 39 49
rect 41 60 48 61
rect 41 56 43 60
rect 47 56 48 60
rect 41 53 48 56
rect 41 49 43 53
rect 47 49 48 53
rect 41 46 48 49
rect 21 42 27 46
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect -2 69 58 78
rect -2 68 3 69
rect 2 65 3 68
rect 7 68 58 69
rect 7 65 8 68
rect 2 62 8 65
rect 2 58 3 62
rect 7 58 8 62
rect 13 62 17 63
rect 13 55 17 58
rect 22 60 28 68
rect 42 60 48 68
rect 22 56 23 60
rect 27 56 28 60
rect 32 56 33 60
rect 37 56 38 60
rect 2 51 13 54
rect 32 53 38 56
rect 2 50 17 51
rect 2 22 6 50
rect 23 49 33 53
rect 37 49 38 53
rect 42 56 43 60
rect 47 56 48 60
rect 42 53 48 56
rect 42 49 43 53
rect 47 49 48 53
rect 23 46 27 49
rect 17 42 27 46
rect 33 42 46 46
rect 17 38 21 42
rect 25 34 29 38
rect 33 34 38 38
rect 17 30 21 34
rect 17 26 28 30
rect 2 18 14 22
rect 18 18 19 22
rect 2 17 19 18
rect 24 21 28 26
rect 34 25 38 34
rect 42 33 46 38
rect 43 23 47 24
rect 24 19 43 21
rect 24 17 47 19
rect -2 8 3 12
rect 7 8 25 12
rect 29 8 58 12
rect -2 2 58 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
<< ntransistor >>
rect 10 16 12 30
rect 20 16 22 30
rect 32 18 34 30
rect 39 18 41 30
<< ptransistor >>
rect 9 42 11 70
rect 19 42 21 70
rect 29 46 31 61
rect 39 46 41 61
<< polycontact >>
rect 17 34 21 38
rect 29 34 33 38
rect 42 38 46 42
<< ndcontact >>
rect 14 18 18 22
rect 43 19 47 23
rect 3 8 7 12
rect 25 8 29 12
<< pdcontact >>
rect 3 65 7 69
rect 3 58 7 62
rect 13 58 17 62
rect 13 51 17 55
rect 23 56 27 60
rect 33 56 37 60
rect 33 49 37 53
rect 43 56 47 60
rect 43 49 47 53
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
<< psubstratepdiff >>
rect 0 2 56 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 56 2
rect 0 -3 56 -2
<< nsubstratendiff >>
rect 0 82 56 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 56 82
rect 0 77 56 78
<< labels >>
rlabel polysilicon 15 36 15 36 6 zn
rlabel metal1 4 32 4 32 6 z
rlabel metal1 12 20 12 20 6 z
rlabel polycontact 19 36 19 36 6 zn
rlabel metal1 12 52 12 52 6 z
rlabel metal1 28 6 28 6 6 vss
rlabel metal1 28 36 28 36 6 a
rlabel metal1 36 28 36 28 6 a
rlabel metal1 36 44 36 44 6 b
rlabel metal1 30 51 30 51 6 zn
rlabel metal1 35 54 35 54 6 zn
rlabel metal1 28 74 28 74 6 vdd
rlabel metal1 35 19 35 19 6 zn
rlabel metal1 44 36 44 36 6 b
<< end >>
