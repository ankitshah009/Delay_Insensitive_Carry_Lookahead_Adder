magic
tech scmos
timestamp 1179386269
<< checkpaint >>
rect -22 -25 118 105
<< ab >>
rect 0 0 96 80
<< pwell >>
rect -4 -7 100 36
<< nwell >>
rect -4 36 100 87
<< polysilicon >>
rect 9 66 11 71
rect 19 66 21 71
rect 29 66 31 71
rect 39 66 41 71
rect 49 66 51 71
rect 59 66 61 71
rect 69 66 71 71
rect 79 58 81 63
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 39 39 41 42
rect 49 39 51 42
rect 59 39 61 42
rect 69 39 71 42
rect 79 39 81 42
rect 9 38 15 39
rect 9 34 10 38
rect 14 34 15 38
rect 9 33 15 34
rect 19 38 33 39
rect 19 34 27 38
rect 31 34 33 38
rect 19 33 33 34
rect 12 30 14 33
rect 19 30 21 33
rect 31 30 33 33
rect 38 38 51 39
rect 38 34 39 38
rect 43 34 46 38
rect 50 34 51 38
rect 38 33 51 34
rect 55 38 62 39
rect 55 34 57 38
rect 61 34 62 38
rect 55 33 62 34
rect 66 38 81 39
rect 66 34 76 38
rect 80 34 81 38
rect 66 33 81 34
rect 38 30 40 33
rect 48 30 50 33
rect 55 30 57 33
rect 66 30 68 33
rect 12 6 14 10
rect 19 6 21 10
rect 31 6 33 10
rect 38 6 40 10
rect 48 6 50 10
rect 55 6 57 10
rect 66 6 68 10
<< ndiffusion >>
rect 5 29 12 30
rect 5 25 6 29
rect 10 25 12 29
rect 5 22 12 25
rect 5 18 6 22
rect 10 18 12 22
rect 5 17 12 18
rect 7 10 12 17
rect 14 10 19 30
rect 21 15 31 30
rect 21 11 24 15
rect 28 11 31 15
rect 21 10 31 11
rect 33 10 38 30
rect 40 29 48 30
rect 40 25 42 29
rect 46 25 48 29
rect 40 22 48 25
rect 40 18 42 22
rect 46 18 48 22
rect 40 10 48 18
rect 50 10 55 30
rect 57 22 66 30
rect 57 18 60 22
rect 64 18 66 22
rect 57 15 66 18
rect 57 11 60 15
rect 64 11 66 15
rect 57 10 66 11
rect 68 29 75 30
rect 68 25 70 29
rect 74 25 75 29
rect 68 22 75 25
rect 68 18 70 22
rect 74 18 75 22
rect 68 17 75 18
rect 68 10 73 17
<< pdiffusion >>
rect 2 65 9 66
rect 2 61 3 65
rect 7 61 9 65
rect 2 42 9 61
rect 11 62 19 66
rect 11 58 13 62
rect 17 58 19 62
rect 11 54 19 58
rect 11 50 13 54
rect 17 50 19 54
rect 11 42 19 50
rect 21 65 29 66
rect 21 61 23 65
rect 27 61 29 65
rect 21 42 29 61
rect 31 62 39 66
rect 31 58 33 62
rect 37 58 39 62
rect 31 54 39 58
rect 31 50 33 54
rect 37 50 39 54
rect 31 42 39 50
rect 41 65 49 66
rect 41 61 43 65
rect 47 61 49 65
rect 41 42 49 61
rect 51 62 59 66
rect 51 58 53 62
rect 57 58 59 62
rect 51 55 59 58
rect 51 51 53 55
rect 57 51 59 55
rect 51 42 59 51
rect 61 65 69 66
rect 61 61 63 65
rect 67 61 69 65
rect 61 57 69 61
rect 61 53 63 57
rect 67 53 69 57
rect 61 42 69 53
rect 71 58 76 66
rect 71 54 79 58
rect 71 50 73 54
rect 77 50 79 54
rect 71 47 79 50
rect 71 43 73 47
rect 77 43 79 47
rect 71 42 79 43
rect 81 57 89 58
rect 81 53 83 57
rect 87 53 89 57
rect 81 49 89 53
rect 81 45 83 49
rect 87 45 89 49
rect 81 42 89 45
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect -2 68 98 78
rect 3 65 7 68
rect 23 65 27 68
rect 3 60 7 61
rect 13 62 17 63
rect 43 65 47 68
rect 23 60 27 61
rect 33 62 38 63
rect 13 55 17 58
rect 2 54 17 55
rect 37 58 38 62
rect 63 65 67 68
rect 43 60 47 61
rect 53 62 57 63
rect 33 54 38 58
rect 53 55 57 58
rect 2 50 13 54
rect 17 50 33 54
rect 37 51 53 54
rect 63 57 67 61
rect 83 57 87 68
rect 63 52 67 53
rect 73 54 77 55
rect 37 50 57 51
rect 2 25 6 50
rect 73 47 77 50
rect 17 39 23 46
rect 10 38 23 39
rect 14 34 23 38
rect 10 33 23 34
rect 27 43 73 46
rect 83 49 87 53
rect 83 44 87 45
rect 27 42 77 43
rect 27 38 31 42
rect 57 38 61 42
rect 27 33 31 34
rect 17 30 23 33
rect 35 30 39 38
rect 43 34 46 38
rect 50 34 51 38
rect 57 30 61 34
rect 74 38 86 39
rect 74 34 76 38
rect 80 34 86 38
rect 74 33 86 34
rect 10 25 11 29
rect 17 26 39 30
rect 42 29 47 30
rect 5 22 11 25
rect 46 25 47 29
rect 57 29 74 30
rect 57 26 70 29
rect 42 22 47 25
rect 70 22 74 25
rect 5 18 6 22
rect 10 18 42 22
rect 46 18 47 22
rect 59 18 60 22
rect 64 18 65 22
rect 59 15 65 18
rect 70 17 74 18
rect 82 17 86 33
rect 23 12 24 15
rect -2 11 24 12
rect 28 12 29 15
rect 59 12 60 15
rect 28 11 60 12
rect 64 12 65 15
rect 64 11 98 12
rect -2 2 98 11
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
<< ntransistor >>
rect 12 10 14 30
rect 19 10 21 30
rect 31 10 33 30
rect 38 10 40 30
rect 48 10 50 30
rect 55 10 57 30
rect 66 10 68 30
<< ptransistor >>
rect 9 42 11 66
rect 19 42 21 66
rect 29 42 31 66
rect 39 42 41 66
rect 49 42 51 66
rect 59 42 61 66
rect 69 42 71 66
rect 79 42 81 58
<< polycontact >>
rect 10 34 14 38
rect 27 34 31 38
rect 39 34 43 38
rect 46 34 50 38
rect 57 34 61 38
rect 76 34 80 38
<< ndcontact >>
rect 6 25 10 29
rect 6 18 10 22
rect 24 11 28 15
rect 42 25 46 29
rect 42 18 46 22
rect 60 18 64 22
rect 60 11 64 15
rect 70 25 74 29
rect 70 18 74 22
<< pdcontact >>
rect 3 61 7 65
rect 13 58 17 62
rect 13 50 17 54
rect 23 61 27 65
rect 33 58 37 62
rect 33 50 37 54
rect 43 61 47 65
rect 53 58 57 62
rect 53 51 57 55
rect 63 61 67 65
rect 63 53 67 57
rect 73 50 77 54
rect 73 43 77 47
rect 83 53 87 57
rect 83 45 87 49
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
rect 90 -2 94 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
rect 90 78 94 82
<< psubstratepdiff >>
rect 0 2 96 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 96 2
rect 0 -3 96 -2
<< nsubstratendiff >>
rect 0 82 96 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 96 82
rect 0 77 96 78
<< labels >>
rlabel polycontact 58 36 58 36 6 an
rlabel metal1 12 20 12 20 6 z
rlabel metal1 4 40 4 40 6 z
rlabel polycontact 12 36 12 36 6 b
rlabel metal1 12 52 12 52 6 z
rlabel metal1 20 20 20 20 6 z
rlabel metal1 28 20 28 20 6 z
rlabel metal1 28 28 28 28 6 b
rlabel metal1 29 39 29 39 6 an
rlabel metal1 20 36 20 36 6 b
rlabel metal1 28 52 28 52 6 z
rlabel metal1 20 52 20 52 6 z
rlabel metal1 48 6 48 6 6 vss
rlabel metal1 36 20 36 20 6 z
rlabel metal1 36 28 36 28 6 b
rlabel ndcontact 44 20 44 20 6 z
rlabel metal1 44 36 44 36 6 b
rlabel metal1 44 52 44 52 6 z
rlabel metal1 52 52 52 52 6 z
rlabel metal1 36 56 36 56 6 z
rlabel metal1 48 74 48 74 6 vdd
rlabel metal1 72 23 72 23 6 an
rlabel polycontact 59 36 59 36 6 an
rlabel metal1 76 36 76 36 6 a
rlabel metal1 75 48 75 48 6 an
rlabel metal1 84 28 84 28 6 a
<< end >>
