magic
tech scmos
timestamp 1179386692
<< checkpaint >>
rect -22 -25 94 105
<< ab >>
rect 0 0 72 80
<< pwell >>
rect -4 -7 76 36
<< nwell >>
rect -4 36 76 87
<< polysilicon >>
rect 9 70 11 74
rect 16 70 18 74
rect 27 70 29 74
rect 34 70 36 74
rect 44 70 46 74
rect 51 70 53 74
rect 61 70 63 74
rect 9 39 11 45
rect 2 38 12 39
rect 2 34 3 38
rect 7 34 12 38
rect 2 33 12 34
rect 16 35 18 45
rect 27 35 29 45
rect 34 42 36 45
rect 44 42 46 45
rect 34 40 46 42
rect 40 39 46 40
rect 40 35 41 39
rect 45 35 46 39
rect 16 33 36 35
rect 40 34 46 35
rect 10 30 12 33
rect 20 30 22 33
rect 34 30 36 33
rect 51 30 53 45
rect 61 39 63 42
rect 57 38 63 39
rect 57 34 58 38
rect 62 34 63 38
rect 57 33 63 34
rect 61 30 63 33
rect 34 29 53 30
rect 34 28 45 29
rect 44 25 45 28
rect 49 28 53 29
rect 49 25 50 28
rect 44 24 50 25
rect 10 6 12 10
rect 20 6 22 10
rect 61 11 63 16
<< ndiffusion >>
rect 2 12 10 30
rect 2 8 3 12
rect 7 10 10 12
rect 12 29 20 30
rect 12 25 14 29
rect 18 25 20 29
rect 12 10 20 25
rect 22 12 31 30
rect 56 26 61 30
rect 53 21 61 26
rect 53 17 55 21
rect 59 17 61 21
rect 53 16 61 17
rect 63 29 70 30
rect 63 25 65 29
rect 69 25 70 29
rect 63 22 70 25
rect 63 18 65 22
rect 69 18 70 22
rect 63 16 70 18
rect 22 10 25 12
rect 7 8 8 10
rect 2 7 8 8
rect 24 8 25 10
rect 29 8 31 12
rect 24 7 31 8
<< pdiffusion >>
rect 4 62 9 70
rect 2 61 9 62
rect 2 57 3 61
rect 7 57 9 61
rect 2 54 9 57
rect 2 50 3 54
rect 7 50 9 54
rect 2 49 9 50
rect 4 45 9 49
rect 11 45 16 70
rect 18 69 27 70
rect 18 65 21 69
rect 25 65 27 69
rect 18 62 27 65
rect 18 58 21 62
rect 25 58 27 62
rect 18 45 27 58
rect 29 45 34 70
rect 36 62 44 70
rect 36 58 38 62
rect 42 58 44 62
rect 36 55 44 58
rect 36 51 38 55
rect 42 51 44 55
rect 36 45 44 51
rect 46 45 51 70
rect 53 69 61 70
rect 53 65 55 69
rect 59 65 61 69
rect 53 62 61 65
rect 53 58 55 62
rect 59 58 61 62
rect 53 45 61 58
rect 56 42 61 45
rect 63 55 68 70
rect 63 54 70 55
rect 63 50 65 54
rect 69 50 70 54
rect 63 47 70 50
rect 63 43 65 47
rect 69 43 70 47
rect 63 42 70 43
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect -2 69 74 78
rect -2 68 21 69
rect 20 65 21 68
rect 25 68 55 69
rect 25 65 26 68
rect 2 61 7 63
rect 2 57 3 61
rect 20 62 26 65
rect 54 65 55 68
rect 59 68 74 69
rect 59 65 60 68
rect 20 58 21 62
rect 25 58 26 62
rect 38 62 46 63
rect 42 58 46 62
rect 54 62 60 65
rect 54 58 55 62
rect 59 58 60 62
rect 2 54 7 57
rect 38 57 46 58
rect 38 55 42 57
rect 2 50 3 54
rect 7 51 38 54
rect 7 50 42 51
rect 65 54 69 55
rect 2 38 7 39
rect 2 34 3 38
rect 2 21 7 34
rect 13 25 14 29
rect 18 25 22 50
rect 65 47 69 50
rect 50 39 54 47
rect 26 35 41 39
rect 45 35 46 39
rect 26 33 46 35
rect 50 38 62 39
rect 50 34 58 38
rect 50 33 62 34
rect 26 21 30 33
rect 65 29 69 43
rect 44 25 45 29
rect 49 25 65 29
rect 65 22 69 25
rect 2 17 30 21
rect 54 17 55 21
rect 59 17 60 21
rect 65 17 69 18
rect 54 12 60 17
rect -2 8 3 12
rect 7 8 25 12
rect 29 8 74 12
rect -2 2 74 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
<< ntransistor >>
rect 10 10 12 30
rect 20 10 22 30
rect 61 16 63 30
<< ptransistor >>
rect 9 45 11 70
rect 16 45 18 70
rect 27 45 29 70
rect 34 45 36 70
rect 44 45 46 70
rect 51 45 53 70
rect 61 42 63 70
<< polycontact >>
rect 3 34 7 38
rect 41 35 45 39
rect 58 34 62 38
rect 45 25 49 29
<< ndcontact >>
rect 3 8 7 12
rect 14 25 18 29
rect 55 17 59 21
rect 65 25 69 29
rect 65 18 69 22
rect 25 8 29 12
<< pdcontact >>
rect 3 57 7 61
rect 3 50 7 54
rect 21 65 25 69
rect 21 58 25 62
rect 38 58 42 62
rect 38 51 42 55
rect 55 65 59 69
rect 55 58 59 62
rect 65 50 69 54
rect 65 43 69 47
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
<< psubstratepdiff >>
rect 0 2 72 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 72 2
rect 0 -3 72 -2
<< nsubstratendiff >>
rect 0 82 72 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 72 82
rect 0 77 72 78
<< labels >>
rlabel polycontact 47 27 47 27 6 an
rlabel metal1 4 28 4 28 6 b
rlabel pdcontact 4 60 4 60 6 z
rlabel metal1 20 40 20 40 6 z
rlabel metal1 20 52 20 52 6 z
rlabel metal1 12 52 12 52 6 z
rlabel metal1 36 6 36 6 6 vss
rlabel metal1 28 28 28 28 6 b
rlabel metal1 36 36 36 36 6 b
rlabel metal1 36 52 36 52 6 z
rlabel metal1 28 52 28 52 6 z
rlabel metal1 36 74 36 74 6 vdd
rlabel polycontact 44 36 44 36 6 b
rlabel metal1 52 40 52 40 6 a
rlabel metal1 44 60 44 60 6 z
rlabel metal1 56 27 56 27 6 an
rlabel polycontact 60 36 60 36 6 a
rlabel metal1 67 36 67 36 6 an
<< end >>
