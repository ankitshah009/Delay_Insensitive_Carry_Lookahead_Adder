magic
tech scmos
timestamp 1185038928
<< checkpaint >>
rect -22 -24 102 124
<< ab >>
rect 0 0 80 100
<< pwell >>
rect -2 -4 82 49
<< nwell >>
rect -2 49 82 104
<< polysilicon >>
rect 55 95 57 98
rect 67 95 69 98
rect 11 85 13 88
rect 31 85 33 88
rect 43 85 45 88
rect 11 63 13 65
rect 11 62 23 63
rect 11 61 18 62
rect 17 58 18 61
rect 22 58 23 62
rect 17 57 23 58
rect 3 52 9 53
rect 3 48 4 52
rect 8 51 9 52
rect 31 51 33 65
rect 8 49 33 51
rect 8 48 9 49
rect 3 47 9 48
rect 31 29 33 49
rect 43 53 45 65
rect 43 52 51 53
rect 43 48 46 52
rect 50 48 51 52
rect 43 47 51 48
rect 37 42 43 43
rect 37 38 38 42
rect 42 41 43 42
rect 55 41 57 55
rect 67 41 69 55
rect 42 39 69 41
rect 42 38 43 39
rect 37 37 43 38
rect 43 32 51 33
rect 31 27 37 29
rect 17 26 23 27
rect 17 23 18 26
rect 11 22 18 23
rect 22 22 23 26
rect 35 25 37 27
rect 43 28 46 32
rect 50 28 51 32
rect 43 27 51 28
rect 43 25 45 27
rect 55 25 57 39
rect 67 25 69 39
rect 11 21 23 22
rect 11 19 13 21
rect 11 6 13 9
rect 35 2 37 5
rect 43 2 45 5
rect 55 2 57 5
rect 67 2 69 5
<< ndiffusion >>
rect 3 22 9 23
rect 3 18 4 22
rect 8 19 9 22
rect 27 22 35 25
rect 8 18 11 19
rect 3 9 11 18
rect 13 12 21 19
rect 13 9 16 12
rect 15 8 16 9
rect 20 8 21 12
rect 15 7 21 8
rect 27 18 28 22
rect 32 18 35 22
rect 27 5 35 18
rect 37 5 43 25
rect 45 12 55 25
rect 45 8 48 12
rect 52 8 55 12
rect 45 5 55 8
rect 57 22 67 25
rect 57 18 60 22
rect 64 18 67 22
rect 57 5 67 18
rect 69 22 77 25
rect 69 18 72 22
rect 76 18 77 22
rect 69 12 77 18
rect 69 8 72 12
rect 76 8 77 12
rect 69 5 77 8
<< pdiffusion >>
rect 15 92 29 93
rect 15 88 16 92
rect 20 88 24 92
rect 28 88 29 92
rect 47 92 55 95
rect 47 88 48 92
rect 52 88 55 92
rect 15 85 29 88
rect 47 85 55 88
rect 3 82 11 85
rect 3 78 4 82
rect 8 78 11 82
rect 3 72 11 78
rect 3 68 4 72
rect 8 68 11 72
rect 3 65 11 68
rect 13 65 31 85
rect 33 82 43 85
rect 33 78 36 82
rect 40 78 43 82
rect 33 72 43 78
rect 33 68 36 72
rect 40 68 43 72
rect 33 65 43 68
rect 45 65 55 85
rect 47 55 55 65
rect 57 82 67 95
rect 57 78 60 82
rect 64 78 67 82
rect 57 72 67 78
rect 57 68 60 72
rect 64 68 67 72
rect 57 62 67 68
rect 57 58 60 62
rect 64 58 67 62
rect 57 55 67 58
rect 69 92 77 95
rect 69 88 72 92
rect 76 88 77 92
rect 69 82 77 88
rect 69 78 72 82
rect 76 78 77 82
rect 69 72 77 78
rect 69 68 72 72
rect 76 68 77 72
rect 69 62 77 68
rect 69 58 72 62
rect 76 58 77 62
rect 69 55 77 58
<< metal1 >>
rect -2 92 82 101
rect -2 88 16 92
rect 20 88 24 92
rect 28 88 48 92
rect 52 88 72 92
rect 76 88 82 92
rect -2 87 82 88
rect 3 82 9 83
rect 35 82 41 83
rect 59 82 65 83
rect 3 78 4 82
rect 8 78 9 82
rect 3 77 9 78
rect 4 73 8 77
rect 3 72 9 73
rect 3 68 4 72
rect 8 68 9 72
rect 3 67 9 68
rect 4 53 8 67
rect 17 62 23 82
rect 35 78 36 82
rect 40 78 41 82
rect 35 77 41 78
rect 37 73 41 77
rect 35 72 41 73
rect 35 68 36 72
rect 40 68 41 72
rect 35 67 41 68
rect 17 58 18 62
rect 22 58 23 62
rect 3 52 9 53
rect 3 48 4 52
rect 8 48 9 52
rect 3 47 9 48
rect 4 23 8 47
rect 17 26 23 58
rect 3 22 9 23
rect 3 18 4 22
rect 8 18 9 22
rect 17 22 18 26
rect 22 22 23 26
rect 37 43 41 67
rect 47 53 53 82
rect 45 52 53 53
rect 45 48 46 52
rect 50 48 53 52
rect 45 47 53 48
rect 37 42 43 43
rect 37 38 38 42
rect 42 38 43 42
rect 37 37 43 38
rect 17 18 23 22
rect 27 22 33 23
rect 37 22 41 37
rect 47 33 53 47
rect 45 32 53 33
rect 45 28 46 32
rect 50 28 53 32
rect 45 27 53 28
rect 27 18 28 22
rect 32 18 41 22
rect 47 18 53 27
rect 57 78 60 82
rect 64 78 65 82
rect 57 77 65 78
rect 71 82 77 87
rect 71 78 72 82
rect 76 78 77 82
rect 57 73 63 77
rect 57 72 65 73
rect 57 68 60 72
rect 64 68 65 72
rect 57 67 65 68
rect 71 72 77 78
rect 71 68 72 72
rect 76 68 77 72
rect 57 63 63 67
rect 57 62 65 63
rect 57 58 60 62
rect 64 58 65 62
rect 57 57 65 58
rect 71 62 77 68
rect 71 58 72 62
rect 76 58 77 62
rect 71 57 77 58
rect 57 23 63 57
rect 57 22 65 23
rect 57 18 60 22
rect 64 18 65 22
rect 3 17 9 18
rect 27 17 33 18
rect 59 17 65 18
rect 71 22 77 23
rect 71 18 72 22
rect 76 18 77 22
rect 71 13 77 18
rect -2 12 82 13
rect -2 8 16 12
rect 20 8 48 12
rect 52 8 72 12
rect 76 8 82 12
rect -2 -1 82 8
<< ntransistor >>
rect 11 9 13 19
rect 35 5 37 25
rect 43 5 45 25
rect 55 5 57 25
rect 67 5 69 25
<< ptransistor >>
rect 11 65 13 85
rect 31 65 33 85
rect 43 65 45 85
rect 55 55 57 95
rect 67 55 69 95
<< polycontact >>
rect 18 58 22 62
rect 4 48 8 52
rect 46 48 50 52
rect 38 38 42 42
rect 18 22 22 26
rect 46 28 50 32
<< ndcontact >>
rect 4 18 8 22
rect 16 8 20 12
rect 28 18 32 22
rect 48 8 52 12
rect 60 18 64 22
rect 72 18 76 22
rect 72 8 76 12
<< pdcontact >>
rect 16 88 20 92
rect 24 88 28 92
rect 48 88 52 92
rect 4 78 8 82
rect 4 68 8 72
rect 36 78 40 82
rect 36 68 40 72
rect 60 78 64 82
rect 60 68 64 72
rect 60 58 64 62
rect 72 88 76 92
rect 72 78 76 82
rect 72 68 76 72
rect 72 58 76 62
<< labels >>
rlabel metal1 20 50 20 50 6 i0
rlabel metal1 20 50 20 50 6 i0
rlabel metal1 40 6 40 6 6 vss
rlabel metal1 40 6 40 6 6 vss
rlabel metal1 50 50 50 50 6 i1
rlabel metal1 60 50 60 50 6 q
rlabel metal1 50 50 50 50 6 i1
rlabel metal1 60 50 60 50 6 q
rlabel metal1 40 94 40 94 6 vdd
rlabel metal1 40 94 40 94 6 vdd
<< end >>
