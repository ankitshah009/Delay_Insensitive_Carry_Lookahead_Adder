magic
tech scmos
timestamp 1179385194
<< checkpaint >>
rect -22 -25 110 105
<< ab >>
rect 0 0 88 80
<< pwell >>
rect -4 -7 92 36
<< nwell >>
rect -4 36 92 87
<< polysilicon >>
rect 9 70 11 74
rect 16 70 18 74
rect 26 70 28 74
rect 33 70 35 74
rect 43 70 45 74
rect 53 70 55 74
rect 63 70 65 74
rect 73 70 75 74
rect 9 33 11 42
rect 16 39 18 42
rect 26 39 28 42
rect 16 38 28 39
rect 16 37 23 38
rect 20 34 23 37
rect 27 34 28 38
rect 20 33 28 34
rect 9 32 15 33
rect 9 28 10 32
rect 14 28 15 32
rect 9 27 15 28
rect 10 24 12 27
rect 20 24 22 33
rect 33 31 35 42
rect 43 39 45 42
rect 53 39 55 42
rect 63 39 65 42
rect 43 38 49 39
rect 43 34 44 38
rect 48 34 49 38
rect 43 33 49 34
rect 53 38 65 39
rect 53 34 54 38
rect 58 37 65 38
rect 73 39 75 42
rect 73 38 79 39
rect 58 34 59 37
rect 53 33 59 34
rect 73 34 74 38
rect 78 34 79 38
rect 73 33 79 34
rect 33 30 39 31
rect 47 30 49 33
rect 54 30 56 33
rect 33 26 34 30
rect 38 26 39 30
rect 33 25 39 26
rect 10 9 12 14
rect 20 9 22 14
rect 47 8 49 13
rect 54 8 56 13
<< ndiffusion >>
rect 2 14 10 24
rect 12 22 20 24
rect 12 18 14 22
rect 18 18 20 22
rect 12 14 20 18
rect 22 14 31 24
rect 42 23 47 30
rect 40 22 47 23
rect 40 18 41 22
rect 45 18 47 22
rect 40 17 47 18
rect 2 12 8 14
rect 2 8 3 12
rect 7 8 8 12
rect 24 12 31 14
rect 42 13 47 17
rect 49 13 54 30
rect 56 25 63 30
rect 56 21 58 25
rect 62 21 63 25
rect 56 18 63 21
rect 56 14 58 18
rect 62 14 63 18
rect 56 13 63 14
rect 2 7 8 8
rect 24 8 25 12
rect 29 8 31 12
rect 24 7 31 8
<< pdiffusion >>
rect 4 64 9 70
rect 2 63 9 64
rect 2 59 3 63
rect 7 59 9 63
rect 2 58 9 59
rect 4 42 9 58
rect 11 42 16 70
rect 18 55 26 70
rect 18 51 20 55
rect 24 51 26 55
rect 18 48 26 51
rect 18 44 20 48
rect 24 44 26 48
rect 18 42 26 44
rect 28 42 33 70
rect 35 62 43 70
rect 35 58 37 62
rect 41 58 43 62
rect 35 55 43 58
rect 35 51 37 55
rect 41 51 43 55
rect 35 42 43 51
rect 45 69 53 70
rect 45 65 47 69
rect 51 65 53 69
rect 45 62 53 65
rect 45 58 47 62
rect 51 58 53 62
rect 45 42 53 58
rect 55 61 63 70
rect 55 57 57 61
rect 61 57 63 61
rect 55 54 63 57
rect 55 50 57 54
rect 61 50 63 54
rect 55 42 63 50
rect 65 69 73 70
rect 65 65 67 69
rect 71 65 73 69
rect 65 62 73 65
rect 65 58 67 62
rect 71 58 73 62
rect 65 42 73 58
rect 75 63 80 70
rect 75 62 82 63
rect 75 58 77 62
rect 81 58 82 62
rect 75 55 82 58
rect 75 51 77 55
rect 81 51 82 55
rect 75 50 82 51
rect 75 42 80 50
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect -2 69 90 78
rect -2 68 47 69
rect 46 65 47 68
rect 51 68 67 69
rect 51 65 52 68
rect 2 59 3 63
rect 7 62 41 63
rect 7 59 37 62
rect 46 62 52 65
rect 66 65 67 68
rect 71 68 90 69
rect 71 65 72 68
rect 66 62 72 65
rect 46 58 47 62
rect 51 58 52 62
rect 57 61 61 62
rect 37 55 41 58
rect 2 51 20 55
rect 24 51 25 55
rect 2 50 25 51
rect 66 58 67 62
rect 71 58 72 62
rect 77 62 81 63
rect 57 54 61 57
rect 77 55 81 58
rect 41 51 57 54
rect 37 50 57 51
rect 61 51 77 54
rect 61 50 81 51
rect 2 22 6 50
rect 19 48 25 50
rect 10 32 14 47
rect 19 44 20 48
rect 24 44 25 48
rect 33 38 39 46
rect 22 34 23 38
rect 27 34 39 38
rect 43 42 78 46
rect 43 38 49 42
rect 74 38 78 42
rect 43 34 44 38
rect 48 34 49 38
rect 53 34 54 38
rect 58 34 70 38
rect 14 28 34 30
rect 10 26 34 28
rect 38 26 39 30
rect 58 25 62 26
rect 2 18 14 22
rect 18 18 41 22
rect 45 18 47 22
rect 58 18 62 21
rect 66 17 70 34
rect 74 25 78 34
rect 58 12 62 14
rect -2 8 3 12
rect 7 8 25 12
rect 29 8 90 12
rect -2 2 90 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
<< ntransistor >>
rect 10 14 12 24
rect 20 14 22 24
rect 47 13 49 30
rect 54 13 56 30
<< ptransistor >>
rect 9 42 11 70
rect 16 42 18 70
rect 26 42 28 70
rect 33 42 35 70
rect 43 42 45 70
rect 53 42 55 70
rect 63 42 65 70
rect 73 42 75 70
<< polycontact >>
rect 23 34 27 38
rect 10 28 14 32
rect 44 34 48 38
rect 54 34 58 38
rect 74 34 78 38
rect 34 26 38 30
<< ndcontact >>
rect 14 18 18 22
rect 41 18 45 22
rect 3 8 7 12
rect 58 21 62 25
rect 58 14 62 18
rect 25 8 29 12
<< pdcontact >>
rect 3 59 7 63
rect 20 51 24 55
rect 20 44 24 48
rect 37 58 41 62
rect 37 51 41 55
rect 47 65 51 69
rect 47 58 51 62
rect 57 57 61 61
rect 57 50 61 54
rect 67 65 71 69
rect 67 58 71 62
rect 77 58 81 62
rect 77 51 81 55
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
<< psubstratepdiff >>
rect 0 2 88 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 88 2
rect 0 -3 88 -2
<< nsubstratendiff >>
rect 0 82 88 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 88 82
rect 0 77 88 78
<< labels >>
rlabel metal1 12 20 12 20 6 z
rlabel metal1 4 40 4 40 6 z
rlabel metal1 12 40 12 40 6 b
rlabel metal1 20 20 20 20 6 z
rlabel metal1 20 28 20 28 6 b
rlabel metal1 28 20 28 20 6 z
rlabel metal1 28 28 28 28 6 b
rlabel metal1 28 36 28 36 6 c
rlabel metal1 20 52 20 52 6 z
rlabel metal1 44 6 44 6 6 vss
rlabel metal1 36 20 36 20 6 z
rlabel polycontact 36 28 36 28 6 b
rlabel ndcontact 44 20 44 20 6 z
rlabel metal1 36 40 36 40 6 c
rlabel metal1 39 56 39 56 6 n1
rlabel metal1 21 61 21 61 6 n1
rlabel metal1 44 74 44 74 6 vdd
rlabel metal1 68 24 68 24 6 a1
rlabel metal1 52 44 52 44 6 a2
rlabel metal1 60 36 60 36 6 a1
rlabel metal1 60 44 60 44 6 a2
rlabel metal1 68 44 68 44 6 a2
rlabel metal1 59 56 59 56 6 n1
rlabel metal1 76 32 76 32 6 a2
rlabel metal1 79 56 79 56 6 n1
rlabel pdcontact 59 52 59 52 6 n1
<< end >>
