.subckt nd2v3x05 a b vdd vss z
*   SPICE3 file   created from nd2v3x05.ext -      technology: scmos
m00 z      b      vdd    vdd p w=10u  l=2.3636u ad=40p      pd=18u      as=146p     ps=58u
m01 vdd    a      z      vdd p w=10u  l=2.3636u ad=146p     pd=58u      as=40p      ps=18u
m02 w1     b      z      vss n w=17u  l=2.3636u ad=42.5p    pd=22u      as=111p     ps=48u
m03 vss    a      w1     vss n w=17u  l=2.3636u ad=136p     pd=50u      as=42.5p    ps=22u
C0  z      a      0.052f
C1  vss    vdd    0.005f
C2  a      b      0.079f
C3  z      vdd    0.037f
C4  b      vdd    0.138f
C5  vss    z      0.048f
C6  vss    b      0.010f
C7  z      b      0.071f
C8  a      vdd    0.018f
C9  vss    a      0.058f
C11 z      vss    0.006f
C12 a      vss    0.021f
C13 b      vss    0.023f
.ends
