magic
tech scmos
timestamp 1179387159
<< checkpaint >>
rect -22 -25 62 105
<< ab >>
rect 0 0 40 80
<< pwell >>
rect -4 -7 44 36
<< nwell >>
rect -4 36 44 87
<< polysilicon >>
rect 22 70 24 74
rect 29 70 31 74
rect 9 60 11 65
rect 9 39 11 42
rect 22 39 24 49
rect 29 46 31 49
rect 29 45 35 46
rect 29 41 30 45
rect 34 41 35 45
rect 29 40 35 41
rect 9 38 15 39
rect 9 34 10 38
rect 14 34 15 38
rect 9 33 15 34
rect 19 38 25 39
rect 19 34 20 38
rect 24 34 25 38
rect 19 33 25 34
rect 9 30 11 33
rect 19 30 21 33
rect 29 30 31 40
rect 9 16 11 21
rect 19 19 21 24
rect 29 19 31 24
<< ndiffusion >>
rect 2 29 9 30
rect 2 25 3 29
rect 7 25 9 29
rect 2 24 9 25
rect 4 21 9 24
rect 11 24 19 30
rect 21 29 29 30
rect 21 25 23 29
rect 27 25 29 29
rect 21 24 29 25
rect 31 24 38 30
rect 11 21 17 24
rect 13 17 17 21
rect 33 17 38 24
rect 13 16 19 17
rect 13 12 14 16
rect 18 12 19 16
rect 13 11 19 12
rect 32 16 38 17
rect 32 12 33 16
rect 37 12 38 16
rect 32 11 38 12
<< pdiffusion >>
rect 13 69 22 70
rect 13 65 14 69
rect 18 65 22 69
rect 13 60 22 65
rect 2 59 9 60
rect 2 55 3 59
rect 7 55 9 59
rect 2 52 9 55
rect 2 48 3 52
rect 7 48 9 52
rect 2 47 9 48
rect 4 42 9 47
rect 11 49 22 60
rect 24 49 29 70
rect 31 63 36 70
rect 31 62 38 63
rect 31 58 33 62
rect 37 58 38 62
rect 31 57 38 58
rect 31 49 36 57
rect 11 42 19 49
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect -2 69 42 78
rect -2 68 14 69
rect 13 65 14 68
rect 18 68 42 69
rect 18 65 19 68
rect 2 62 6 63
rect 2 59 15 62
rect 2 55 3 59
rect 7 58 15 59
rect 21 58 33 62
rect 37 58 38 62
rect 2 52 7 55
rect 21 54 25 58
rect 2 48 3 52
rect 2 47 7 48
rect 10 50 25 54
rect 2 30 6 47
rect 10 38 14 50
rect 34 46 38 55
rect 17 45 38 46
rect 17 42 30 45
rect 29 41 30 42
rect 34 42 38 45
rect 34 41 35 42
rect 17 34 20 38
rect 24 34 38 38
rect 2 29 7 30
rect 2 25 3 29
rect 10 29 14 34
rect 10 25 23 29
rect 27 25 28 29
rect 34 25 38 34
rect 2 24 7 25
rect 13 12 14 16
rect 18 12 19 16
rect 32 12 33 16
rect 37 12 38 16
rect -2 2 42 12
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
<< ntransistor >>
rect 9 21 11 30
rect 19 24 21 30
rect 29 24 31 30
<< ptransistor >>
rect 9 42 11 60
rect 22 49 24 70
rect 29 49 31 70
<< polycontact >>
rect 30 41 34 45
rect 10 34 14 38
rect 20 34 24 38
<< ndcontact >>
rect 3 25 7 29
rect 23 25 27 29
rect 14 12 18 16
rect 33 12 37 16
<< pdcontact >>
rect 14 65 18 69
rect 3 55 7 59
rect 3 48 7 52
rect 33 58 37 62
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
<< psubstratepdiff >>
rect 0 2 40 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 40 2
rect 0 -3 40 -2
<< nsubstratendiff >>
rect 0 82 40 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 40 82
rect 0 77 40 78
<< labels >>
rlabel polycontact 12 36 12 36 6 zn
rlabel metal1 4 44 4 44 6 z
rlabel metal1 12 39 12 39 6 zn
rlabel metal1 12 60 12 60 6 z
rlabel metal1 20 6 20 6 6 vss
rlabel metal1 20 36 20 36 6 a
rlabel metal1 19 27 19 27 6 zn
rlabel metal1 28 36 28 36 6 a
rlabel metal1 28 44 28 44 6 b
rlabel metal1 20 44 20 44 6 b
rlabel metal1 20 74 20 74 6 vdd
rlabel metal1 36 28 36 28 6 a
rlabel metal1 36 52 36 52 6 b
rlabel metal1 29 60 29 60 6 zn
<< end >>
