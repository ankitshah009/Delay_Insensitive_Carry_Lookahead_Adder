magic
tech scmos
timestamp 1179385279
<< checkpaint >>
rect -22 -25 94 105
<< ab >>
rect 0 0 72 80
<< pwell >>
rect -4 -7 76 36
<< nwell >>
rect -4 36 76 87
<< polysilicon >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 39 70 41 74
rect 51 70 53 74
rect 61 70 63 74
rect 9 40 11 43
rect 9 39 15 40
rect 9 35 10 39
rect 14 35 15 39
rect 9 34 15 35
rect 19 39 21 43
rect 29 39 31 43
rect 19 38 31 39
rect 39 40 41 43
rect 51 40 53 43
rect 61 40 63 43
rect 39 38 54 40
rect 19 34 26 38
rect 30 34 31 38
rect 41 34 42 38
rect 46 34 54 38
rect 58 39 64 40
rect 58 35 59 39
rect 63 35 64 39
rect 58 34 64 35
rect 19 33 31 34
rect 20 29 22 33
rect 35 29 37 34
rect 41 33 54 34
rect 42 29 44 33
rect 52 29 54 33
rect 59 29 61 34
rect 20 9 22 14
rect 35 8 37 16
rect 42 12 44 16
rect 52 12 54 16
rect 59 8 61 16
rect 35 6 61 8
<< ndiffusion >>
rect 15 23 20 29
rect 13 22 20 23
rect 13 18 14 22
rect 18 18 20 22
rect 13 17 20 18
rect 15 14 20 17
rect 22 16 35 29
rect 37 16 42 29
rect 44 22 52 29
rect 44 18 46 22
rect 50 18 52 22
rect 44 16 52 18
rect 54 16 59 29
rect 61 16 69 29
rect 22 15 33 16
rect 22 14 26 15
rect 24 11 26 14
rect 30 11 33 15
rect 24 10 33 11
rect 63 12 69 16
rect 63 8 64 12
rect 68 8 69 12
rect 63 7 69 8
<< pdiffusion >>
rect 43 72 49 73
rect 43 70 44 72
rect 2 69 9 70
rect 2 65 3 69
rect 7 65 9 69
rect 2 62 9 65
rect 2 58 3 62
rect 7 58 9 62
rect 2 43 9 58
rect 11 63 19 70
rect 11 59 13 63
rect 17 59 19 63
rect 11 43 19 59
rect 21 54 29 70
rect 21 50 23 54
rect 27 50 29 54
rect 21 43 29 50
rect 31 62 39 70
rect 31 58 33 62
rect 37 58 39 62
rect 31 55 39 58
rect 31 51 33 55
rect 37 51 39 55
rect 31 43 39 51
rect 41 68 44 70
rect 48 70 49 72
rect 48 68 51 70
rect 41 43 51 68
rect 53 62 61 70
rect 53 58 55 62
rect 59 58 61 62
rect 53 55 61 58
rect 53 51 55 55
rect 59 51 61 55
rect 53 43 61 51
rect 63 69 70 70
rect 63 65 65 69
rect 69 65 70 69
rect 63 61 70 65
rect 63 57 65 61
rect 69 57 70 61
rect 63 43 70 57
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect -2 72 74 78
rect -2 69 44 72
rect -2 68 3 69
rect 2 65 3 68
rect 7 68 44 69
rect 48 69 74 72
rect 48 68 65 69
rect 7 65 8 68
rect 2 62 8 65
rect 69 68 74 69
rect 2 58 3 62
rect 7 58 8 62
rect 12 59 13 63
rect 17 62 59 63
rect 17 59 33 62
rect 37 59 55 62
rect 33 55 37 58
rect 55 55 59 58
rect 65 61 69 65
rect 65 56 69 57
rect 2 54 28 55
rect 2 50 23 54
rect 27 50 28 54
rect 33 50 37 51
rect 2 22 6 50
rect 42 46 46 55
rect 55 50 59 51
rect 10 42 63 46
rect 10 39 14 42
rect 57 39 63 42
rect 10 34 14 35
rect 25 34 26 38
rect 30 34 31 38
rect 25 30 31 34
rect 17 26 31 30
rect 41 34 42 38
rect 46 34 47 38
rect 57 35 59 39
rect 57 34 63 35
rect 41 30 47 34
rect 41 26 55 30
rect 2 18 14 22
rect 18 18 46 22
rect 50 18 55 22
rect 25 12 26 15
rect -2 11 26 12
rect 30 12 31 15
rect 30 11 64 12
rect -2 8 64 11
rect 68 8 74 12
rect -2 2 74 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
<< ntransistor >>
rect 20 14 22 29
rect 35 16 37 29
rect 42 16 44 29
rect 52 16 54 29
rect 59 16 61 29
<< ptransistor >>
rect 9 43 11 70
rect 19 43 21 70
rect 29 43 31 70
rect 39 43 41 70
rect 51 43 53 70
rect 61 43 63 70
<< polycontact >>
rect 10 35 14 39
rect 26 34 30 38
rect 42 34 46 38
rect 59 35 63 39
<< ndcontact >>
rect 14 18 18 22
rect 46 18 50 22
rect 26 11 30 15
rect 64 8 68 12
<< pdcontact >>
rect 3 65 7 69
rect 3 58 7 62
rect 13 59 17 63
rect 23 50 27 54
rect 33 58 37 62
rect 33 51 37 55
rect 44 68 48 72
rect 55 58 59 62
rect 55 51 59 55
rect 65 65 69 69
rect 65 57 69 61
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
<< psubstratepdiff >>
rect 0 2 72 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 72 2
rect 0 -3 72 -2
<< nsubstratendiff >>
rect 0 82 72 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 72 82
rect 0 77 72 78
<< labels >>
rlabel metal1 4 40 4 40 6 z
rlabel metal1 12 20 12 20 6 z
rlabel metal1 20 20 20 20 6 z
rlabel metal1 20 28 20 28 6 b
rlabel metal1 20 44 20 44 6 a1
rlabel metal1 20 52 20 52 6 z
rlabel metal1 12 52 12 52 6 z
rlabel metal1 36 6 36 6 6 vss
rlabel metal1 28 20 28 20 6 z
rlabel metal1 36 20 36 20 6 z
rlabel metal1 28 32 28 32 6 b
rlabel metal1 28 44 28 44 6 a1
rlabel metal1 36 44 36 44 6 a1
rlabel metal1 35 56 35 56 6 n1
rlabel metal1 36 74 36 74 6 vdd
rlabel metal1 44 20 44 20 6 z
rlabel metal1 52 20 52 20 6 z
rlabel metal1 52 28 52 28 6 a2
rlabel metal1 44 32 44 32 6 a2
rlabel metal1 52 44 52 44 6 a1
rlabel metal1 44 48 44 48 6 a1
rlabel metal1 60 40 60 40 6 a1
rlabel metal1 57 56 57 56 6 n1
rlabel pdcontact 35 61 35 61 6 n1
<< end >>
