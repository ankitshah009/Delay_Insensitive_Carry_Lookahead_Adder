.subckt nr2v1x3 a b vdd vss z
*   SPICE3 file   created from nr2v1x3.ext -      technology: scmos
m00 w1     b      z      vdd p w=28u  l=2.3636u ad=70p      pd=33u      as=130p     ps=47.3333u
m01 vdd    a      w1     vdd p w=28u  l=2.3636u ad=140p     pd=47.3333u as=70p      ps=33u
m02 w2     a      vdd    vdd p w=28u  l=2.3636u ad=70p      pd=33u      as=140p     ps=47.3333u
m03 z      b      w2     vdd p w=28u  l=2.3636u ad=130p     pd=47.3333u as=70p      ps=33u
m04 w3     b      z      vdd p w=28u  l=2.3636u ad=70p      pd=33u      as=130p     ps=47.3333u
m05 vdd    a      w3     vdd p w=28u  l=2.3636u ad=140p     pd=47.3333u as=70p      ps=33u
m06 z      b      vss    vss n w=20u  l=2.3636u ad=80p      pd=28u      as=165p     ps=46.5u
m07 vss    a      z      vss n w=20u  l=2.3636u ad=165p     pd=46.5u    as=80p      ps=28u
m08 z      b      vss    vss n w=20u  l=2.3636u ad=80p      pd=28u      as=165p     ps=46.5u
m09 vss    a      z      vss n w=20u  l=2.3636u ad=165p     pd=46.5u    as=80p      ps=28u
C0  w3     vdd    0.005f
C1  z      b      0.425f
C2  w1     vdd    0.005f
C3  a      vdd    0.082f
C4  vss    a      0.051f
C5  vss    vdd    0.003f
C6  w1     z      0.010f
C7  w2     a      0.007f
C8  z      a      0.305f
C9  w2     vdd    0.005f
C10 a      b      0.426f
C11 z      vdd    0.214f
C12 b      vdd    0.042f
C13 vss    z      0.437f
C14 w2     z      0.010f
C15 w3     a      0.007f
C16 vss    b      0.098f
C18 z      vss    0.012f
C19 a      vss    0.038f
C20 b      vss    0.041f
.ends
