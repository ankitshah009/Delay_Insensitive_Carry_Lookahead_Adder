.subckt nr2v0x1 a b vdd vss z
*   SPICE3 file   created from nr2v0x1.ext -      technology: scmos
m00 w1     a      vdd    vdd p w=26u  l=2.3636u ad=130p     pd=36u      as=182p     ps=66u
m01 z      b      w1     vdd p w=26u  l=2.3636u ad=182p     pd=66u      as=130p     ps=36u
m02 z      a      vss    vss n w=18u  l=2.3636u ad=90p      pd=28u      as=126p     ps=50u
m03 vss    b      z      vss n w=18u  l=2.3636u ad=126p     pd=50u      as=90p      ps=28u
C0  z      b      0.224f
C1  vss    a      0.041f
C2  z      vdd    0.010f
C3  b      vdd    0.006f
C4  vss    z      0.073f
C5  z      w1     0.021f
C6  vss    b      0.024f
C7  z      a      0.214f
C8  b      a      0.176f
C9  a      vdd    0.017f
C11 z      vss    0.006f
C12 b      vss    0.062f
C13 a      vss    0.061f
.ends
