.subckt nd3_x05 a b c vdd vss z
*   SPICE3 file   created from nd3_x05.ext -      technology: scmos
m00 vdd    c      z      vdd p w=12u  l=2.3636u ad=92p      pd=34.6667u as=66p      ps=28u
m01 z      b      vdd    vdd p w=12u  l=2.3636u ad=66p      pd=28u      as=92p      ps=34.6667u
m02 vdd    a      z      vdd p w=12u  l=2.3636u ad=92p      pd=34.6667u as=66p      ps=28u
m03 w1     c      z      vss n w=12u  l=2.3636u ad=36p      pd=18u      as=78p      ps=40u
m04 w2     b      w1     vss n w=12u  l=2.3636u ad=36p      pd=18u      as=36p      ps=18u
m05 vss    a      w2     vss n w=12u  l=2.3636u ad=96p      pd=40u      as=36p      ps=18u
C0  z      c      0.217f
C1  a      b      0.201f
C2  b      c      0.155f
C3  a      vdd    0.006f
C4  c      vdd    0.021f
C5  vss    a      0.042f
C6  w1     a      0.009f
C7  vss    c      0.015f
C8  z      b      0.133f
C9  a      c      0.138f
C10 z      vdd    0.092f
C11 b      vdd    0.065f
C12 vss    z      0.045f
C13 w2     a      0.013f
C14 w1     z      0.003f
C15 z      a      0.070f
C17 z      vss    0.029f
C18 a      vss    0.029f
C19 b      vss    0.033f
C20 c      vss    0.037f
.ends
