.subckt inv_x4 i nq vdd vss
*   SPICE3 file   created from inv_x4.ext -      technology: scmos
m00 nq     i      vdd    vdd p w=40u  l=2.3636u ad=221.176p pd=58.8235u as=320p     ps=98.8235u
m01 vdd    i      nq     vdd p w=28u  l=2.3636u ad=224p     pd=69.1765u as=154.824p ps=41.1765u
m02 nq     i      vss    vss n w=20u  l=2.3636u ad=100p     pd=30u      as=160p     ps=56u
m03 vss    i      nq     vss n w=20u  l=2.3636u ad=160p     pd=56u      as=100p     ps=30u
C0  nq     i      0.504f
C1  vss    nq     0.099f
C2  vss    i      0.072f
C3  nq     vdd    0.150f
C4  vdd    i      0.129f
C6  nq     vss    0.018f
C8  i      vss    0.073f
.ends
