magic
tech scmos
timestamp 1179385917
<< checkpaint >>
rect -22 -25 54 105
<< ab >>
rect 0 0 32 80
<< pwell >>
rect -4 -7 36 36
<< nwell >>
rect -4 36 36 87
<< polysilicon >>
rect 9 63 11 67
rect 19 61 21 65
rect 9 39 11 42
rect 19 39 21 42
rect 9 38 21 39
rect 9 34 15 38
rect 19 34 21 38
rect 9 33 21 34
rect 9 30 11 33
rect 19 30 21 33
rect 9 6 11 10
rect 19 6 21 10
<< ndiffusion >>
rect 2 22 9 30
rect 2 18 3 22
rect 7 18 9 22
rect 2 15 9 18
rect 2 11 3 15
rect 7 11 9 15
rect 2 10 9 11
rect 11 28 19 30
rect 11 24 13 28
rect 17 24 19 28
rect 11 21 19 24
rect 11 17 13 21
rect 17 17 19 21
rect 11 10 19 17
rect 21 22 28 30
rect 21 18 23 22
rect 27 18 28 22
rect 21 15 28 18
rect 21 11 23 15
rect 27 11 28 15
rect 21 10 28 11
<< pdiffusion >>
rect 2 62 9 63
rect 2 58 3 62
rect 7 58 9 62
rect 2 42 9 58
rect 11 61 16 63
rect 11 60 19 61
rect 11 56 13 60
rect 17 56 19 60
rect 11 53 19 56
rect 11 49 13 53
rect 17 49 19 53
rect 11 42 19 49
rect 21 60 28 61
rect 21 56 23 60
rect 27 56 28 60
rect 21 53 28 56
rect 21 49 23 53
rect 27 49 28 53
rect 21 42 28 49
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect -2 68 34 78
rect 2 62 8 68
rect 2 58 3 62
rect 7 58 8 62
rect 22 60 28 68
rect 12 56 13 60
rect 17 56 18 60
rect 12 55 18 56
rect 2 53 18 55
rect 2 49 13 53
rect 17 49 18 53
rect 22 56 23 60
rect 27 56 28 60
rect 22 53 28 56
rect 22 49 23 53
rect 27 49 28 53
rect 2 29 6 49
rect 17 39 23 46
rect 10 38 23 39
rect 10 34 15 38
rect 19 34 23 38
rect 10 33 23 34
rect 2 28 17 29
rect 2 25 13 28
rect 2 18 3 22
rect 7 18 8 22
rect 2 15 8 18
rect 13 21 17 24
rect 13 16 17 17
rect 22 18 23 22
rect 27 18 28 22
rect 2 12 3 15
rect -2 11 3 12
rect 7 12 8 15
rect 22 15 28 18
rect 22 12 23 15
rect 7 11 23 12
rect 27 12 28 15
rect 27 11 34 12
rect -2 2 34 11
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
<< ntransistor >>
rect 9 10 11 30
rect 19 10 21 30
<< ptransistor >>
rect 9 42 11 63
rect 19 42 21 61
<< polycontact >>
rect 15 34 19 38
<< ndcontact >>
rect 3 18 7 22
rect 3 11 7 15
rect 13 24 17 28
rect 13 17 17 21
rect 23 18 27 22
rect 23 11 27 15
<< pdcontact >>
rect 3 58 7 62
rect 13 56 17 60
rect 13 49 17 53
rect 23 56 27 60
rect 23 49 27 53
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
<< psubstratepdiff >>
rect 0 2 32 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 32 2
rect 0 -3 32 -2
<< nsubstratendiff >>
rect 0 82 32 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 32 82
rect 0 77 32 78
<< labels >>
rlabel metal1 4 40 4 40 6 z
rlabel metal1 12 36 12 36 6 a
rlabel metal1 12 52 12 52 6 z
rlabel metal1 16 6 16 6 6 vss
rlabel metal1 20 40 20 40 6 a
rlabel metal1 16 74 16 74 6 vdd
<< end >>
