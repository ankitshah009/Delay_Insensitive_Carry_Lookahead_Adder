magic
tech scmos
timestamp 1179385568
<< checkpaint >>
rect -22 -22 54 94
<< ab >>
rect 0 0 32 72
<< pwell >>
rect -4 -4 36 32
<< nwell >>
rect -4 32 36 76
<< polysilicon >>
rect 9 50 11 55
rect 21 58 27 59
rect 21 54 22 58
rect 26 54 27 58
rect 21 53 27 54
rect 21 50 23 53
rect 9 35 11 38
rect 9 34 15 35
rect 9 30 10 34
rect 14 30 15 34
rect 9 29 15 30
rect 9 26 11 29
rect 21 26 23 38
rect 9 15 11 20
rect 21 15 23 20
<< ndiffusion >>
rect 2 25 9 26
rect 2 21 3 25
rect 7 21 9 25
rect 2 20 9 21
rect 11 25 21 26
rect 11 21 14 25
rect 18 21 21 25
rect 11 20 21 21
rect 23 25 30 26
rect 23 21 25 25
rect 29 21 30 25
rect 23 20 30 21
<< pdiffusion >>
rect 13 68 19 69
rect 13 64 14 68
rect 18 64 19 68
rect 13 50 19 64
rect 4 44 9 50
rect 2 43 9 44
rect 2 39 3 43
rect 7 39 9 43
rect 2 38 9 39
rect 11 38 21 50
rect 23 44 28 50
rect 23 43 30 44
rect 23 39 25 43
rect 29 39 30 43
rect 23 38 30 39
<< metal1 >>
rect -2 68 34 72
rect -2 64 4 68
rect 8 64 14 68
rect 18 64 24 68
rect 28 64 34 68
rect 18 58 30 59
rect 18 54 22 58
rect 26 54 30 58
rect 18 53 30 54
rect 2 45 14 51
rect 18 45 22 53
rect 2 43 7 45
rect 2 39 3 43
rect 2 38 7 39
rect 25 43 29 44
rect 2 25 6 38
rect 25 34 29 39
rect 9 30 10 34
rect 14 30 29 34
rect 14 25 18 26
rect 2 21 3 25
rect 7 21 8 25
rect 14 8 18 21
rect 25 25 29 30
rect 25 20 29 21
rect -2 4 4 8
rect 8 4 24 8
rect 28 4 34 8
rect -2 0 34 4
<< ntransistor >>
rect 9 20 11 26
rect 21 20 23 26
<< ptransistor >>
rect 9 38 11 50
rect 21 38 23 50
<< polycontact >>
rect 22 54 26 58
rect 10 30 14 34
<< ndcontact >>
rect 3 21 7 25
rect 14 21 18 25
rect 25 21 29 25
<< pdcontact >>
rect 14 64 18 68
rect 3 39 7 43
rect 25 39 29 43
<< psubstratepcontact >>
rect 4 4 8 8
rect 24 4 28 8
<< nsubstratencontact >>
rect 4 64 8 68
rect 24 64 28 68
<< psubstratepdiff >>
rect 3 8 29 9
rect 3 4 4 8
rect 8 4 24 8
rect 28 4 29 8
rect 3 3 29 4
<< nsubstratendiff >>
rect 3 68 9 69
rect 3 64 4 68
rect 8 64 9 68
rect 3 57 9 64
rect 23 68 29 69
rect 23 64 24 68
rect 28 64 29 68
rect 23 63 29 64
<< labels >>
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 48 12 48 6 z
rlabel metal1 16 4 16 4 6 vss
rlabel metal1 20 52 20 52 6 a
rlabel metal1 16 68 16 68 6 vdd
rlabel metal1 19 32 19 32 6 an
rlabel metal1 28 56 28 56 6 a
<< end >>
