magic
tech scmos
timestamp 1179386278
<< checkpaint >>
rect -22 -25 134 105
<< ab >>
rect 0 0 112 80
<< pwell >>
rect -4 -7 116 36
<< nwell >>
rect -4 36 116 87
<< polysilicon >>
rect 9 68 11 73
rect 19 68 21 73
rect 29 68 31 73
rect 39 68 41 73
rect 49 68 51 73
rect 59 68 61 73
rect 69 60 71 65
rect 79 60 81 65
rect 91 64 93 69
rect 101 64 103 69
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 39 39 41 42
rect 9 38 15 39
rect 9 34 10 38
rect 14 34 15 38
rect 9 33 15 34
rect 19 38 31 39
rect 19 34 26 38
rect 30 34 31 38
rect 19 33 31 34
rect 35 38 41 39
rect 35 34 36 38
rect 40 35 41 38
rect 49 35 51 42
rect 59 39 61 42
rect 69 39 71 42
rect 59 38 71 39
rect 40 34 54 35
rect 35 33 54 34
rect 12 30 14 33
rect 19 30 21 33
rect 29 30 31 33
rect 36 30 38 33
rect 52 30 54 33
rect 59 34 60 38
rect 64 34 71 38
rect 79 39 81 42
rect 91 39 93 42
rect 101 39 103 42
rect 79 38 87 39
rect 79 35 82 38
rect 59 33 71 34
rect 59 30 61 33
rect 69 30 71 33
rect 76 34 82 35
rect 86 34 87 38
rect 76 33 87 34
rect 91 38 103 39
rect 91 34 98 38
rect 102 34 103 38
rect 91 33 103 34
rect 76 30 78 33
rect 91 30 93 33
rect 101 30 103 33
rect 91 14 93 19
rect 101 15 103 19
rect 12 6 14 10
rect 19 6 21 10
rect 29 6 31 10
rect 36 6 38 10
rect 52 6 54 10
rect 59 6 61 10
rect 69 6 71 10
rect 76 6 78 10
<< ndiffusion >>
rect 4 15 12 30
rect 4 11 6 15
rect 10 11 12 15
rect 4 10 12 11
rect 14 10 19 30
rect 21 22 29 30
rect 21 18 23 22
rect 27 18 29 22
rect 21 10 29 18
rect 31 10 36 30
rect 38 15 52 30
rect 38 11 43 15
rect 47 11 52 15
rect 38 10 52 11
rect 54 10 59 30
rect 61 22 69 30
rect 61 18 63 22
rect 67 18 69 22
rect 61 10 69 18
rect 71 10 76 30
rect 78 22 91 30
rect 78 18 82 22
rect 86 19 91 22
rect 93 29 101 30
rect 93 25 95 29
rect 99 25 101 29
rect 93 19 101 25
rect 103 24 110 30
rect 103 20 105 24
rect 109 20 110 24
rect 103 19 110 20
rect 86 18 89 19
rect 78 15 89 18
rect 78 11 82 15
rect 86 11 89 15
rect 78 10 89 11
<< pdiffusion >>
rect 2 67 9 68
rect 2 63 3 67
rect 7 63 9 67
rect 2 42 9 63
rect 11 61 19 68
rect 11 57 13 61
rect 17 57 19 61
rect 11 54 19 57
rect 11 50 13 54
rect 17 50 19 54
rect 11 42 19 50
rect 21 67 29 68
rect 21 63 23 67
rect 27 63 29 67
rect 21 42 29 63
rect 31 62 39 68
rect 31 58 33 62
rect 37 58 39 62
rect 31 54 39 58
rect 31 50 33 54
rect 37 50 39 54
rect 31 42 39 50
rect 41 67 49 68
rect 41 63 43 67
rect 47 63 49 67
rect 41 42 49 63
rect 51 54 59 68
rect 51 50 53 54
rect 57 50 59 54
rect 51 47 59 50
rect 51 43 53 47
rect 57 43 59 47
rect 51 42 59 43
rect 61 60 67 68
rect 83 60 91 64
rect 61 59 69 60
rect 61 55 63 59
rect 67 55 69 59
rect 61 42 69 55
rect 71 54 79 60
rect 71 50 73 54
rect 77 50 79 54
rect 71 47 79 50
rect 71 43 73 47
rect 77 43 79 47
rect 71 42 79 43
rect 81 59 91 60
rect 81 55 83 59
rect 87 55 91 59
rect 81 42 91 55
rect 93 54 101 64
rect 93 50 95 54
rect 99 50 101 54
rect 93 47 101 50
rect 93 43 95 47
rect 99 43 101 47
rect 93 42 101 43
rect 103 63 110 64
rect 103 59 105 63
rect 109 59 110 63
rect 103 42 110 59
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect -2 68 114 78
rect 3 67 7 68
rect 3 62 7 63
rect 23 67 27 68
rect 43 67 47 68
rect 23 62 27 63
rect 33 62 38 63
rect 43 62 47 63
rect 13 61 17 62
rect 13 55 17 57
rect 2 54 17 55
rect 37 58 38 62
rect 33 54 38 58
rect 63 59 67 68
rect 83 59 87 68
rect 104 63 110 68
rect 104 59 105 63
rect 109 59 110 63
rect 63 54 67 55
rect 73 54 78 55
rect 83 54 87 55
rect 95 54 99 55
rect 2 50 13 54
rect 17 50 33 54
rect 37 50 53 54
rect 57 50 58 54
rect 2 22 6 50
rect 53 47 58 50
rect 25 42 49 46
rect 57 46 58 47
rect 77 50 78 54
rect 73 47 78 50
rect 57 43 73 46
rect 77 43 78 47
rect 95 47 99 50
rect 53 42 78 43
rect 82 43 95 46
rect 82 42 99 43
rect 10 38 14 39
rect 25 38 31 42
rect 45 38 49 42
rect 82 38 86 42
rect 106 38 110 55
rect 25 34 26 38
rect 30 34 31 38
rect 35 34 36 38
rect 40 34 41 38
rect 45 34 60 38
rect 64 34 71 38
rect 97 34 98 38
rect 102 34 110 38
rect 10 30 14 34
rect 35 30 41 34
rect 82 30 86 34
rect 10 29 100 30
rect 10 26 95 29
rect 94 25 95 26
rect 99 25 100 29
rect 105 24 109 25
rect 2 18 23 22
rect 27 18 63 22
rect 67 18 71 22
rect 81 18 82 22
rect 86 18 87 22
rect 81 15 87 18
rect 5 12 6 15
rect -2 11 6 12
rect 10 12 11 15
rect 42 12 43 15
rect 10 11 43 12
rect 47 12 48 15
rect 81 12 82 15
rect 47 11 82 12
rect 86 12 87 15
rect 105 12 109 20
rect 86 11 114 12
rect -2 2 114 11
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
<< ntransistor >>
rect 12 10 14 30
rect 19 10 21 30
rect 29 10 31 30
rect 36 10 38 30
rect 52 10 54 30
rect 59 10 61 30
rect 69 10 71 30
rect 76 10 78 30
rect 91 19 93 30
rect 101 19 103 30
<< ptransistor >>
rect 9 42 11 68
rect 19 42 21 68
rect 29 42 31 68
rect 39 42 41 68
rect 49 42 51 68
rect 59 42 61 68
rect 69 42 71 60
rect 79 42 81 60
rect 91 42 93 64
rect 101 42 103 64
<< polycontact >>
rect 10 34 14 38
rect 26 34 30 38
rect 36 34 40 38
rect 60 34 64 38
rect 82 34 86 38
rect 98 34 102 38
<< ndcontact >>
rect 6 11 10 15
rect 23 18 27 22
rect 43 11 47 15
rect 63 18 67 22
rect 82 18 86 22
rect 95 25 99 29
rect 105 20 109 24
rect 82 11 86 15
<< pdcontact >>
rect 3 63 7 67
rect 13 57 17 61
rect 13 50 17 54
rect 23 63 27 67
rect 33 58 37 62
rect 33 50 37 54
rect 43 63 47 67
rect 53 50 57 54
rect 53 43 57 47
rect 63 55 67 59
rect 73 50 77 54
rect 73 43 77 47
rect 83 55 87 59
rect 95 50 99 54
rect 95 43 99 47
rect 105 59 109 63
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
rect 90 -2 94 2
rect 98 -2 102 2
rect 106 -2 110 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
rect 90 78 94 82
rect 98 78 102 82
rect 106 78 110 82
<< psubstratepdiff >>
rect 0 2 112 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 112 2
rect 0 -3 112 -2
<< nsubstratendiff >>
rect 0 82 112 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 112 82
rect 0 77 112 78
<< labels >>
rlabel ntransistor 13 22 13 22 6 an
rlabel ntransistor 37 22 37 22 6 an
rlabel polycontact 83 36 83 36 6 an
rlabel metal1 12 20 12 20 6 z
rlabel metal1 12 32 12 32 6 an
rlabel metal1 4 40 4 40 6 z
rlabel metal1 12 52 12 52 6 z
rlabel metal1 20 20 20 20 6 z
rlabel metal1 28 20 28 20 6 z
rlabel metal1 36 20 36 20 6 z
rlabel metal1 38 32 38 32 6 an
rlabel metal1 28 40 28 40 6 b
rlabel metal1 36 44 36 44 6 b
rlabel metal1 28 52 28 52 6 z
rlabel metal1 20 52 20 52 6 z
rlabel metal1 36 56 36 56 6 z
rlabel metal1 56 6 56 6 6 vss
rlabel metal1 44 20 44 20 6 z
rlabel metal1 52 20 52 20 6 z
rlabel metal1 60 20 60 20 6 z
rlabel metal1 44 44 44 44 6 b
rlabel metal1 52 36 52 36 6 b
rlabel metal1 60 36 60 36 6 b
rlabel metal1 60 44 60 44 6 z
rlabel metal1 52 52 52 52 6 z
rlabel metal1 44 52 44 52 6 z
rlabel metal1 56 74 56 74 6 vdd
rlabel metal1 68 20 68 20 6 z
rlabel polycontact 84 36 84 36 6 an
rlabel metal1 68 36 68 36 6 b
rlabel metal1 68 44 68 44 6 z
rlabel pdcontact 76 52 76 52 6 z
rlabel ndcontact 97 27 97 27 6 an
rlabel polycontact 100 36 100 36 6 a
rlabel metal1 108 48 108 48 6 a
rlabel metal1 97 48 97 48 6 an
<< end >>
