magic
tech scmos
timestamp 1179387705
<< checkpaint >>
rect -22 -25 94 105
<< ab >>
rect 0 0 72 80
<< pwell >>
rect -4 -7 76 36
<< nwell >>
rect -4 36 76 87
<< polysilicon >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 40 70 42 74
rect 50 70 52 74
rect 40 53 42 56
rect 50 53 52 56
rect 40 52 63 53
rect 40 51 42 52
rect 41 48 42 51
rect 46 51 63 52
rect 46 48 47 51
rect 41 47 47 48
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 9 38 15 39
rect 9 34 10 38
rect 14 34 15 38
rect 9 33 15 34
rect 19 38 25 39
rect 19 34 20 38
rect 24 34 25 38
rect 29 36 33 39
rect 19 33 25 34
rect 12 30 14 33
rect 19 30 21 33
rect 31 30 33 36
rect 41 30 43 47
rect 51 38 57 39
rect 51 34 52 38
rect 56 34 57 38
rect 51 33 57 34
rect 51 30 53 33
rect 61 30 63 51
rect 12 6 14 11
rect 19 6 21 11
rect 31 8 33 23
rect 61 18 63 23
rect 41 12 43 16
rect 51 8 53 16
rect 31 6 53 8
<< ndiffusion >>
rect 7 23 12 30
rect 5 22 12 23
rect 5 18 6 22
rect 10 18 12 22
rect 5 17 12 18
rect 7 11 12 17
rect 14 11 19 30
rect 21 23 31 30
rect 33 29 41 30
rect 33 25 35 29
rect 39 25 41 29
rect 33 23 41 25
rect 21 12 29 23
rect 21 11 24 12
rect 23 8 24 11
rect 28 8 29 12
rect 23 7 29 8
rect 36 16 41 23
rect 43 22 51 30
rect 43 18 45 22
rect 49 18 51 22
rect 43 16 51 18
rect 53 29 61 30
rect 53 25 55 29
rect 59 25 61 29
rect 53 23 61 25
rect 63 28 70 30
rect 63 24 65 28
rect 69 24 70 28
rect 63 23 70 24
rect 53 16 58 23
<< pdiffusion >>
rect 4 63 9 70
rect 2 62 9 63
rect 2 58 3 62
rect 7 58 9 62
rect 2 57 9 58
rect 4 42 9 57
rect 11 54 19 70
rect 11 50 13 54
rect 17 50 19 54
rect 11 42 19 50
rect 21 54 29 70
rect 21 50 23 54
rect 27 50 29 54
rect 21 47 29 50
rect 21 43 23 47
rect 27 43 29 47
rect 21 42 29 43
rect 31 69 40 70
rect 31 65 34 69
rect 38 65 40 69
rect 31 56 40 65
rect 42 62 50 70
rect 42 58 44 62
rect 48 58 50 62
rect 42 56 50 58
rect 52 69 59 70
rect 52 65 54 69
rect 58 65 59 69
rect 52 62 59 65
rect 52 58 54 62
rect 58 58 59 62
rect 52 56 59 58
rect 31 42 38 56
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect -2 69 74 78
rect -2 68 34 69
rect 33 65 34 68
rect 38 68 54 69
rect 38 65 39 68
rect 53 65 54 68
rect 58 68 74 69
rect 58 65 59 68
rect 53 62 59 65
rect 2 58 3 62
rect 7 58 44 62
rect 48 58 49 62
rect 53 58 54 62
rect 58 58 59 62
rect 23 54 27 55
rect 2 50 13 54
rect 17 50 18 54
rect 2 18 6 50
rect 23 47 27 50
rect 10 43 23 46
rect 10 42 27 43
rect 10 38 14 42
rect 31 38 35 58
rect 41 52 55 54
rect 41 48 42 52
rect 46 48 55 52
rect 49 42 55 48
rect 66 38 70 47
rect 19 34 20 38
rect 24 34 48 38
rect 10 30 14 34
rect 10 29 40 30
rect 10 26 35 29
rect 34 25 35 26
rect 39 25 40 29
rect 44 29 48 34
rect 51 34 52 38
rect 56 34 70 38
rect 51 33 70 34
rect 44 25 55 29
rect 59 25 60 29
rect 65 28 69 29
rect 10 18 45 22
rect 49 18 50 22
rect 65 12 69 24
rect -2 8 24 12
rect 28 8 74 12
rect -2 2 74 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
<< ntransistor >>
rect 12 11 14 30
rect 19 11 21 30
rect 31 23 33 30
rect 41 16 43 30
rect 51 16 53 30
rect 61 23 63 30
<< ptransistor >>
rect 9 42 11 70
rect 19 42 21 70
rect 29 42 31 70
rect 40 56 42 70
rect 50 56 52 70
<< polycontact >>
rect 42 48 46 52
rect 10 34 14 38
rect 20 34 24 38
rect 52 34 56 38
<< ndcontact >>
rect 6 18 10 22
rect 35 25 39 29
rect 24 8 28 12
rect 45 18 49 22
rect 55 25 59 29
rect 65 24 69 28
<< pdcontact >>
rect 3 58 7 62
rect 13 50 17 54
rect 23 50 27 54
rect 23 43 27 47
rect 34 65 38 69
rect 44 58 48 62
rect 54 65 58 69
rect 54 58 58 62
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
<< psubstratepdiff >>
rect 0 2 72 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 72 2
rect 0 -3 72 -2
<< nsubstratendiff >>
rect 0 82 72 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 72 82
rect 0 77 72 78
<< labels >>
rlabel polycontact 12 36 12 36 6 bn
rlabel polycontact 22 36 22 36 6 an
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 20 12 20 6 z
rlabel metal1 20 20 20 20 6 z
rlabel polycontact 12 36 12 36 6 bn
rlabel metal1 25 48 25 48 6 bn
rlabel metal1 12 52 12 52 6 z
rlabel metal1 36 6 36 6 6 vss
rlabel metal1 28 20 28 20 6 z
rlabel metal1 25 28 25 28 6 bn
rlabel metal1 36 20 36 20 6 z
rlabel metal1 36 74 36 74 6 vdd
rlabel metal1 44 20 44 20 6 z
rlabel metal1 33 36 33 36 6 an
rlabel metal1 52 48 52 48 6 a
rlabel metal1 44 52 44 52 6 a
rlabel metal1 25 60 25 60 6 an
rlabel metal1 52 27 52 27 6 an
rlabel metal1 60 36 60 36 6 b
rlabel metal1 68 40 68 40 6 b
<< end >>
