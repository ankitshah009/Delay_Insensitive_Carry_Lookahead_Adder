.subckt buf_x2 i q vdd vss
*   SPICE3 file   created from buf_x2.ext -      technology: scmos
m00 vdd    i      w1     vdd p w=12u  l=2.3636u ad=79.3846p pd=23.0769u as=96p      ps=40u
m01 q      w1     vdd    vdd p w=40u  l=2.3636u ad=320p     pd=96u      as=264.615p ps=76.9231u
m02 vss    i      w1     vss n w=6u   l=2.3636u ad=39.6923p pd=13.8462u as=48p      ps=28u
m03 q      w1     vss    vss n w=20u  l=2.3636u ad=160p     pd=56u      as=132.308p ps=46.1538u
C0  vss    q      0.064f
C1  vss    w1     0.038f
C2  q      i      0.485f
C3  q      vdd    0.068f
C4  i      w1     0.377f
C5  w1     vdd    0.021f
C6  vss    i      0.065f
C7  q      w1     0.072f
C8  i      vdd    0.098f
C10 q      vss    0.022f
C11 i      vss    0.040f
C12 w1     vss    0.046f
.ends
