magic
tech scmos
timestamp 1179385492
<< checkpaint >>
rect -22 -22 86 94
<< ab >>
rect 0 0 64 72
<< pwell >>
rect -4 -4 68 32
<< nwell >>
rect -4 32 68 76
<< polysilicon >>
rect 9 65 11 70
rect 19 65 21 70
rect 29 65 31 70
rect 39 56 41 61
rect 49 56 51 61
rect 9 35 11 38
rect 19 35 21 38
rect 29 35 31 38
rect 39 35 41 38
rect 49 35 51 38
rect 9 34 31 35
rect 9 33 26 34
rect 14 30 26 33
rect 30 30 31 34
rect 14 29 31 30
rect 37 34 51 35
rect 37 30 42 34
rect 46 33 51 34
rect 46 30 47 33
rect 37 29 47 30
rect 14 26 16 29
rect 24 26 26 29
rect 37 26 39 29
rect 14 2 16 6
rect 24 2 26 6
rect 37 2 39 7
<< ndiffusion >>
rect 6 18 14 26
rect 6 14 8 18
rect 12 14 14 18
rect 6 11 14 14
rect 6 7 8 11
rect 12 7 14 11
rect 6 6 14 7
rect 16 25 24 26
rect 16 21 18 25
rect 22 21 24 25
rect 16 18 24 21
rect 16 14 18 18
rect 22 14 24 18
rect 16 6 24 14
rect 26 18 37 26
rect 26 14 30 18
rect 34 14 37 18
rect 26 11 37 14
rect 26 7 30 11
rect 34 7 37 11
rect 39 25 46 26
rect 39 21 41 25
rect 45 21 46 25
rect 39 18 46 21
rect 39 14 41 18
rect 45 14 46 18
rect 39 13 46 14
rect 39 7 44 13
rect 26 6 35 7
<< pdiffusion >>
rect 4 51 9 65
rect 2 50 9 51
rect 2 46 3 50
rect 7 46 9 50
rect 2 43 9 46
rect 2 39 3 43
rect 7 39 9 43
rect 2 38 9 39
rect 11 63 19 65
rect 11 59 13 63
rect 17 59 19 63
rect 11 55 19 59
rect 11 51 13 55
rect 17 51 19 55
rect 11 38 19 51
rect 21 50 29 65
rect 21 46 23 50
rect 27 46 29 50
rect 21 43 29 46
rect 21 39 23 43
rect 27 39 29 43
rect 21 38 29 39
rect 31 56 37 65
rect 31 55 39 56
rect 31 51 33 55
rect 37 51 39 55
rect 31 38 39 51
rect 41 50 49 56
rect 41 46 43 50
rect 47 46 49 50
rect 41 43 49 46
rect 41 39 43 43
rect 47 39 49 43
rect 41 38 49 39
rect 51 55 58 56
rect 51 51 53 55
rect 57 51 58 55
rect 51 47 58 51
rect 51 43 53 47
rect 57 43 58 47
rect 51 38 58 43
<< metal1 >>
rect -2 68 66 72
rect -2 64 44 68
rect 48 64 52 68
rect 56 64 66 68
rect 13 63 17 64
rect 13 55 17 59
rect 33 55 37 64
rect 53 55 57 64
rect 2 50 7 51
rect 13 50 17 51
rect 23 50 27 51
rect 33 50 37 51
rect 43 50 47 51
rect 2 46 3 50
rect 2 43 7 46
rect 2 39 3 43
rect 23 43 27 46
rect 7 39 23 42
rect 43 43 47 46
rect 2 38 27 39
rect 33 39 43 42
rect 53 47 57 51
rect 53 42 57 43
rect 33 38 47 39
rect 2 37 14 38
rect 9 26 14 37
rect 33 34 37 38
rect 25 30 26 34
rect 30 30 37 34
rect 41 30 42 34
rect 46 30 55 34
rect 33 26 37 30
rect 9 25 23 26
rect 9 22 18 25
rect 22 21 23 25
rect 33 25 45 26
rect 33 22 41 25
rect 18 18 23 21
rect 49 22 55 30
rect 41 18 45 21
rect 7 14 8 18
rect 12 14 13 18
rect 7 11 13 14
rect 22 14 23 18
rect 18 13 23 14
rect 29 14 30 18
rect 34 14 35 18
rect 7 8 8 11
rect -2 7 8 8
rect 12 8 13 11
rect 29 11 35 14
rect 41 13 45 14
rect 29 8 30 11
rect 12 7 30 8
rect 34 8 35 11
rect 34 7 52 8
rect -2 4 52 7
rect 56 4 66 8
rect -2 0 66 4
<< ntransistor >>
rect 14 6 16 26
rect 24 6 26 26
rect 37 7 39 26
<< ptransistor >>
rect 9 38 11 65
rect 19 38 21 65
rect 29 38 31 65
rect 39 38 41 56
rect 49 38 51 56
<< polycontact >>
rect 26 30 30 34
rect 42 30 46 34
<< ndcontact >>
rect 8 14 12 18
rect 8 7 12 11
rect 18 21 22 25
rect 18 14 22 18
rect 30 14 34 18
rect 30 7 34 11
rect 41 21 45 25
rect 41 14 45 18
<< pdcontact >>
rect 3 46 7 50
rect 3 39 7 43
rect 13 59 17 63
rect 13 51 17 55
rect 23 46 27 50
rect 23 39 27 43
rect 33 51 37 55
rect 43 46 47 50
rect 43 39 47 43
rect 53 51 57 55
rect 53 43 57 47
<< psubstratepcontact >>
rect 52 4 56 8
<< nsubstratencontact >>
rect 44 64 48 68
rect 52 64 56 68
<< psubstratepdiff >>
rect 51 8 57 24
rect 51 4 52 8
rect 56 4 57 8
rect 51 3 57 4
<< nsubstratendiff >>
rect 43 68 57 69
rect 43 64 44 68
rect 48 64 52 68
rect 56 64 57 68
rect 43 63 57 64
<< labels >>
rlabel polysilicon 22 32 22 32 6 an
rlabel metal1 12 32 12 32 6 z
rlabel metal1 4 44 4 44 6 z
rlabel metal1 20 20 20 20 6 z
rlabel metal1 20 40 20 40 6 z
rlabel metal1 32 4 32 4 6 vss
rlabel metal1 43 19 43 19 6 an
rlabel metal1 31 32 31 32 6 an
rlabel polycontact 44 32 44 32 6 a
rlabel metal1 45 44 45 44 6 an
rlabel metal1 32 68 32 68 6 vdd
rlabel metal1 52 28 52 28 6 a
<< end >>
