magic
tech scmos
timestamp 1179387737
<< checkpaint >>
rect -22 -25 94 105
<< ab >>
rect 0 0 72 80
<< pwell >>
rect -4 -7 76 36
<< nwell >>
rect -4 36 76 87
<< polysilicon >>
rect 18 70 20 74
rect 25 70 27 74
rect 36 70 38 74
rect 43 70 45 74
rect 2 62 8 63
rect 2 58 3 62
rect 7 59 8 62
rect 7 58 11 59
rect 2 57 11 58
rect 9 54 11 57
rect 54 61 56 66
rect 54 46 56 50
rect 54 45 64 46
rect 9 30 11 43
rect 18 40 20 43
rect 15 39 21 40
rect 15 35 16 39
rect 20 35 21 39
rect 15 34 21 35
rect 25 30 27 43
rect 36 39 38 43
rect 43 40 45 43
rect 54 41 59 45
rect 63 41 64 45
rect 54 40 64 41
rect 9 28 27 30
rect 31 38 38 39
rect 31 34 32 38
rect 36 34 38 38
rect 31 33 38 34
rect 42 38 64 40
rect 9 25 11 28
rect 21 25 23 28
rect 31 25 33 33
rect 42 30 44 38
rect 51 33 57 34
rect 9 15 11 19
rect 51 29 52 33
rect 56 29 57 33
rect 51 28 57 29
rect 52 24 54 28
rect 61 26 63 38
rect 21 8 23 13
rect 31 9 33 14
rect 42 13 44 18
rect 61 16 63 20
rect 52 6 54 10
<< ndiffusion >>
rect 35 29 42 30
rect 35 25 36 29
rect 40 25 42 29
rect 2 24 9 25
rect 2 20 3 24
rect 7 20 9 24
rect 2 19 9 20
rect 11 19 21 25
rect 13 18 21 19
rect 13 14 14 18
rect 18 14 21 18
rect 13 13 21 14
rect 23 22 31 25
rect 23 18 25 22
rect 29 18 31 22
rect 23 14 31 18
rect 33 18 42 25
rect 44 24 49 30
rect 56 24 61 26
rect 44 23 52 24
rect 44 19 46 23
rect 50 19 52 23
rect 44 18 52 19
rect 33 14 38 18
rect 23 13 28 14
rect 47 10 52 18
rect 54 20 61 24
rect 63 25 70 26
rect 63 21 65 25
rect 69 21 70 25
rect 63 20 70 21
rect 54 14 59 20
rect 54 13 62 14
rect 54 10 57 13
rect 56 9 57 10
rect 61 9 62 13
rect 56 8 62 9
<< pdiffusion >>
rect 11 66 18 70
rect 11 62 12 66
rect 16 62 18 66
rect 11 61 18 62
rect 13 54 18 61
rect 4 49 9 54
rect 2 48 9 49
rect 2 44 3 48
rect 7 44 9 48
rect 2 43 9 44
rect 11 43 18 54
rect 20 43 25 70
rect 27 48 36 70
rect 27 44 30 48
rect 34 44 36 48
rect 27 43 36 44
rect 38 43 43 70
rect 45 64 52 70
rect 45 60 47 64
rect 51 61 52 64
rect 51 60 54 61
rect 45 50 54 60
rect 56 56 61 61
rect 56 55 63 56
rect 56 51 58 55
rect 62 51 63 55
rect 56 50 63 51
rect 45 43 52 50
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect -2 68 74 78
rect 11 66 17 68
rect 2 62 7 63
rect 11 62 12 66
rect 16 62 17 66
rect 47 64 51 68
rect 2 58 3 62
rect 47 59 51 60
rect 2 54 14 58
rect 10 49 14 54
rect 18 51 58 55
rect 62 51 63 55
rect 3 48 7 49
rect 3 30 7 44
rect 18 39 22 51
rect 29 44 30 48
rect 34 47 35 48
rect 34 44 46 47
rect 29 42 46 44
rect 15 35 16 39
rect 20 35 22 39
rect 27 34 32 38
rect 36 34 37 38
rect 27 30 31 34
rect 42 30 46 42
rect 3 26 31 30
rect 35 29 46 30
rect 50 33 54 51
rect 66 47 70 55
rect 58 45 70 47
rect 58 41 59 45
rect 63 41 70 45
rect 50 29 52 33
rect 56 29 69 33
rect 3 24 7 26
rect 35 25 36 29
rect 40 26 46 29
rect 40 25 41 26
rect 65 25 69 29
rect 45 22 46 23
rect 3 19 7 20
rect 14 18 18 19
rect 24 18 25 22
rect 29 19 46 22
rect 50 19 51 23
rect 65 20 69 21
rect 29 18 51 19
rect 14 12 18 14
rect 56 12 57 13
rect -2 9 57 12
rect 61 12 62 13
rect 61 9 74 12
rect -2 2 74 9
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
<< ntransistor >>
rect 9 19 11 25
rect 21 13 23 25
rect 31 14 33 25
rect 42 18 44 30
rect 52 10 54 24
rect 61 20 63 26
<< ptransistor >>
rect 9 43 11 54
rect 18 43 20 70
rect 25 43 27 70
rect 36 43 38 70
rect 43 43 45 70
rect 54 50 56 61
<< polycontact >>
rect 3 58 7 62
rect 16 35 20 39
rect 59 41 63 45
rect 32 34 36 38
rect 52 29 56 33
<< ndcontact >>
rect 36 25 40 29
rect 3 20 7 24
rect 14 14 18 18
rect 25 18 29 22
rect 46 19 50 23
rect 65 21 69 25
rect 57 9 61 13
<< pdcontact >>
rect 12 62 16 66
rect 3 44 7 48
rect 30 44 34 48
rect 47 60 51 64
rect 58 51 62 55
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
<< psubstratepdiff >>
rect 0 2 72 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 72 2
rect 0 -3 72 -2
<< nsubstratendiff >>
rect 0 82 72 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 72 82
rect 0 77 72 78
<< labels >>
rlabel ptransistor 19 54 19 54 6 an
rlabel polycontact 34 36 34 36 6 bn
rlabel polycontact 54 31 54 31 6 an
rlabel metal1 5 34 5 34 6 bn
rlabel polycontact 4 60 4 60 6 b
rlabel metal1 20 45 20 45 6 an
rlabel metal1 12 52 12 52 6 b
rlabel metal1 36 6 36 6 6 vss
rlabel metal1 32 36 32 36 6 bn
rlabel metal1 36 44 36 44 6 z
rlabel metal1 36 74 36 74 6 vdd
rlabel metal1 37 20 37 20 6 n3
rlabel metal1 44 40 44 40 6 z
rlabel metal1 67 26 67 26 6 an
rlabel metal1 59 31 59 31 6 an
rlabel polycontact 60 44 60 44 6 a
rlabel metal1 68 48 68 48 6 a
rlabel metal1 40 53 40 53 6 an
<< end >>
