.subckt iv1_x1 a vdd vss z
*   SPICE3 file   created from iv1_x1.ext -      technology: scmos
m00 vdd    a      z      vdd p w=20u  l=2.3636u ad=180p     pd=58u      as=142p     ps=56u
m01 vss    a      z      vss n w=10u  l=2.3636u ad=132p     pd=50u      as=68p      ps=36u
C0  z      a      0.161f
C1  a      vdd    0.037f
C2  vss    a      0.009f
C3  z      vdd    0.036f
C4  vss    z      0.068f
C6  z      vss    0.012f
C7  a      vss    0.027f
.ends
