.subckt o4_x4 i0 i1 i2 i3 q vdd vss
*   SPICE3 file   created from o4_x4.ext -      technology: scmos
m00 w1     i1     w2     vdd p w=40u  l=2.3636u ad=120p     pd=46u      as=440p     ps=104u
m01 w3     i0     w1     vdd p w=40u  l=2.3636u ad=120p     pd=46u      as=120p     ps=46u
m02 w4     i2     w3     vdd p w=40u  l=2.3636u ad=120p     pd=46u      as=120p     ps=46u
m03 vdd    i3     w4     vdd p w=40u  l=2.3636u ad=240p     pd=65.3333u as=120p     ps=46u
m04 q      w2     vdd    vdd p w=40u  l=2.3636u ad=200p     pd=50u      as=240p     ps=65.3333u
m05 vdd    w2     q      vdd p w=40u  l=2.3636u ad=240p     pd=65.3333u as=200p     ps=50u
m06 w2     i1     vss    vss n w=10u  l=2.3636u ad=50p      pd=20u      as=73.5p    ps=29.5u
m07 vss    i0     w2     vss n w=10u  l=2.3636u ad=73.5p    pd=29.5u    as=50p      ps=20u
m08 w2     i2     vss    vss n w=10u  l=2.3636u ad=50p      pd=20u      as=73.5p    ps=29.5u
m09 vss    i3     w2     vss n w=10u  l=2.3636u ad=73.5p    pd=29.5u    as=50p      ps=20u
m10 q      w2     vss    vss n w=20u  l=2.3636u ad=100p     pd=30u      as=147p     ps=59u
m11 vss    w2     q      vss n w=20u  l=2.3636u ad=147p     pd=59u      as=100p     ps=30u
C0  vdd    w4     0.014f
C1  i3     i0     0.132f
C2  w2     i1     0.482f
C3  vss    i3     0.010f
C4  vdd    w1     0.014f
C5  q      w2     0.330f
C6  i2     i1     0.149f
C7  vss    i0     0.015f
C8  vdd    i3     0.135f
C9  q      i2     0.091f
C10 q      i1     0.022f
C11 vdd    i0     0.053f
C12 w4     i2     0.040f
C13 w2     i3     0.237f
C14 w3     i0     0.041f
C15 w2     i0     0.195f
C16 i3     i2     0.468f
C17 w1     i1     0.027f
C18 vdd    w3     0.014f
C19 vss    w2     0.388f
C20 i3     i1     0.077f
C21 i2     i0     0.497f
C22 vss    i2     0.015f
C23 vdd    w2     0.087f
C24 q      i3     0.230f
C25 i0     i1     0.498f
C26 vdd    i2     0.058f
C27 vss    i1     0.015f
C28 q      i0     0.057f
C29 vss    q      0.141f
C30 vdd    i1     0.041f
C31 q      vdd    0.200f
C32 w2     i2     0.197f
C33 w1     i0     0.014f
C35 q      vss    0.020f
C37 w2     vss    0.054f
C38 i3     vss    0.029f
C39 i2     vss    0.033f
C40 i0     vss    0.034f
C41 i1     vss    0.038f
.ends
