magic
tech scmos
timestamp 1179386216
<< checkpaint >>
rect -22 -25 118 105
<< ab >>
rect 0 0 96 80
<< pwell >>
rect -4 -7 100 36
<< nwell >>
rect -4 36 100 87
<< polysilicon >>
rect 29 70 31 74
rect 39 70 41 74
rect 9 65 11 70
rect 19 65 21 70
rect 9 47 11 50
rect 19 47 21 50
rect 9 46 21 47
rect 9 42 10 46
rect 14 45 21 46
rect 14 42 15 45
rect 51 70 53 74
rect 61 70 63 74
rect 71 70 73 74
rect 81 60 83 65
rect 71 47 73 50
rect 81 47 83 50
rect 71 46 83 47
rect 71 42 74 46
rect 78 42 83 46
rect 9 41 15 42
rect 9 28 11 41
rect 29 37 31 42
rect 15 36 31 37
rect 15 32 16 36
rect 20 35 31 36
rect 39 39 41 42
rect 51 39 53 42
rect 61 39 63 42
rect 71 41 83 42
rect 39 38 53 39
rect 39 35 44 38
rect 20 32 21 35
rect 15 31 21 32
rect 29 28 31 35
rect 36 34 44 35
rect 48 37 53 38
rect 57 38 63 39
rect 48 34 49 37
rect 36 33 49 34
rect 57 34 58 38
rect 62 34 63 38
rect 57 33 63 34
rect 71 36 77 37
rect 36 28 38 33
rect 47 28 49 33
rect 54 31 66 33
rect 54 28 56 31
rect 64 28 66 31
rect 71 32 72 36
rect 76 32 77 36
rect 71 31 77 32
rect 71 28 73 31
rect 81 28 83 41
rect 9 8 11 13
rect 29 6 31 10
rect 36 6 38 10
rect 47 8 49 13
rect 54 8 56 13
rect 64 8 66 13
rect 71 8 73 13
rect 81 8 83 13
<< ndiffusion >>
rect 2 27 9 28
rect 2 23 3 27
rect 7 23 9 27
rect 2 22 9 23
rect 4 13 9 22
rect 11 26 18 28
rect 11 22 13 26
rect 17 22 18 26
rect 22 27 29 28
rect 22 23 23 27
rect 27 23 29 27
rect 22 22 29 23
rect 11 18 18 22
rect 11 14 13 18
rect 17 14 18 18
rect 11 13 18 14
rect 24 10 29 22
rect 31 10 36 28
rect 38 15 47 28
rect 38 11 40 15
rect 44 13 47 15
rect 49 13 54 28
rect 56 22 64 28
rect 56 18 58 22
rect 62 18 64 22
rect 56 13 64 18
rect 66 13 71 28
rect 73 18 81 28
rect 73 14 75 18
rect 79 14 81 18
rect 73 13 81 14
rect 83 27 90 28
rect 83 23 85 27
rect 89 23 90 27
rect 83 22 90 23
rect 83 13 88 22
rect 44 11 45 13
rect 38 10 45 11
<< pdiffusion >>
rect 43 72 49 73
rect 43 70 44 72
rect 23 65 29 70
rect 2 64 9 65
rect 2 60 3 64
rect 7 60 9 64
rect 2 50 9 60
rect 11 63 19 65
rect 11 59 13 63
rect 17 59 19 63
rect 11 56 19 59
rect 11 52 13 56
rect 17 52 19 56
rect 11 50 19 52
rect 21 64 29 65
rect 21 60 23 64
rect 27 60 29 64
rect 21 50 29 60
rect 23 42 29 50
rect 31 63 39 70
rect 31 59 33 63
rect 37 59 39 63
rect 31 47 39 59
rect 31 43 33 47
rect 37 43 39 47
rect 31 42 39 43
rect 41 68 44 70
rect 48 70 49 72
rect 48 68 51 70
rect 41 42 51 68
rect 53 63 61 70
rect 53 59 55 63
rect 59 59 61 63
rect 53 56 61 59
rect 53 52 55 56
rect 59 52 61 56
rect 53 42 61 52
rect 63 69 71 70
rect 63 65 65 69
rect 69 65 71 69
rect 63 62 71 65
rect 63 58 65 62
rect 69 58 71 62
rect 63 50 71 58
rect 73 60 78 70
rect 73 55 81 60
rect 73 51 75 55
rect 79 51 81 55
rect 73 50 81 51
rect 83 59 90 60
rect 83 55 85 59
rect 89 55 90 59
rect 83 50 90 55
rect 63 42 69 50
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect -2 72 98 78
rect -2 68 44 72
rect 48 69 98 72
rect 48 68 65 69
rect 3 64 7 68
rect 23 64 27 68
rect 3 59 7 60
rect 13 63 17 64
rect 64 65 65 68
rect 69 68 98 69
rect 69 65 70 68
rect 23 59 27 60
rect 32 59 33 63
rect 37 59 55 63
rect 59 59 60 63
rect 13 56 17 59
rect 2 47 6 55
rect 55 56 60 59
rect 64 62 70 65
rect 64 58 65 62
rect 69 58 70 62
rect 85 59 89 68
rect 17 52 49 55
rect 13 51 49 52
rect 59 52 60 56
rect 55 51 60 52
rect 67 51 75 55
rect 79 51 80 55
rect 85 54 89 55
rect 2 46 14 47
rect 2 42 10 46
rect 2 41 14 42
rect 18 36 22 51
rect 45 47 49 51
rect 3 32 16 36
rect 20 32 22 36
rect 26 43 33 47
rect 37 43 39 47
rect 45 43 62 47
rect 26 42 39 43
rect 3 27 7 32
rect 26 27 30 42
rect 58 38 62 43
rect 43 34 44 38
rect 3 22 7 23
rect 13 26 17 27
rect 22 23 23 27
rect 27 23 30 27
rect 48 29 52 38
rect 58 33 62 34
rect 67 36 71 51
rect 74 46 86 47
rect 78 42 86 46
rect 74 41 86 42
rect 67 32 72 36
rect 76 32 77 36
rect 82 33 86 41
rect 67 29 71 32
rect 48 27 71 29
rect 48 25 85 27
rect 67 23 85 25
rect 89 23 90 27
rect 13 18 17 22
rect 26 22 30 23
rect 26 18 58 22
rect 62 18 63 22
rect 75 18 79 19
rect 13 12 17 14
rect 39 12 40 15
rect -2 11 40 12
rect 44 12 45 15
rect 75 12 79 14
rect 44 11 98 12
rect -2 2 98 11
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
<< ntransistor >>
rect 9 13 11 28
rect 29 10 31 28
rect 36 10 38 28
rect 47 13 49 28
rect 54 13 56 28
rect 64 13 66 28
rect 71 13 73 28
rect 81 13 83 28
<< ptransistor >>
rect 9 50 11 65
rect 19 50 21 65
rect 29 42 31 70
rect 39 42 41 70
rect 51 42 53 70
rect 61 42 63 70
rect 71 50 73 70
rect 81 50 83 60
<< polycontact >>
rect 10 42 14 46
rect 74 42 78 46
rect 16 32 20 36
rect 44 34 48 38
rect 58 34 62 38
rect 72 32 76 36
<< ndcontact >>
rect 3 23 7 27
rect 13 22 17 26
rect 23 23 27 27
rect 13 14 17 18
rect 40 11 44 15
rect 58 18 62 22
rect 75 14 79 18
rect 85 23 89 27
<< pdcontact >>
rect 3 60 7 64
rect 13 59 17 63
rect 13 52 17 56
rect 23 60 27 64
rect 33 59 37 63
rect 33 43 37 47
rect 44 68 48 72
rect 55 59 59 63
rect 55 52 59 56
rect 65 65 69 69
rect 65 58 69 62
rect 75 51 79 55
rect 85 55 89 59
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
rect 90 -2 94 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
rect 90 78 94 82
<< psubstratepdiff >>
rect 0 2 96 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 96 2
rect 0 -3 96 -2
<< nsubstratendiff >>
rect 0 82 96 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 96 82
rect 0 77 96 78
<< labels >>
rlabel polycontact 18 34 18 34 6 bn
rlabel polycontact 60 35 60 35 6 bn
rlabel polycontact 74 34 74 34 6 an
rlabel metal1 5 29 5 29 6 bn
rlabel polycontact 12 44 12 44 6 b
rlabel metal1 4 48 4 48 6 b
rlabel metal1 15 57 15 57 6 bn
rlabel metal1 12 34 12 34 6 bn
rlabel metal1 28 36 28 36 6 z
rlabel metal1 48 6 48 6 6 vss
rlabel metal1 36 20 36 20 6 z
rlabel metal1 52 20 52 20 6 z
rlabel metal1 44 20 44 20 6 z
rlabel pdcontact 36 44 36 44 6 z
rlabel polycontact 47 36 47 36 6 an
rlabel metal1 48 74 48 74 6 vdd
rlabel ndcontact 60 20 60 20 6 z
rlabel metal1 72 34 72 34 6 an
rlabel metal1 60 40 60 40 6 bn
rlabel polycontact 76 44 76 44 6 a
rlabel metal1 78 25 78 25 6 an
rlabel metal1 84 40 84 40 6 a
rlabel metal1 73 53 73 53 6 an
<< end >>
