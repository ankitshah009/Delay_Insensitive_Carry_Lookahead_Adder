magic
tech scmos
timestamp 1180600768
<< checkpaint >>
rect -22 -22 72 122
<< ab >>
rect 0 0 50 100
<< pwell >>
rect -4 -4 54 48
<< nwell >>
rect -4 48 54 104
<< polysilicon >>
rect 35 94 37 98
rect 15 85 17 89
rect 23 85 25 89
rect 15 53 17 56
rect 11 51 17 53
rect 23 53 25 56
rect 23 52 31 53
rect 11 43 13 51
rect 23 48 26 52
rect 30 48 31 52
rect 23 47 31 48
rect 7 42 13 43
rect 7 38 8 42
rect 12 38 13 42
rect 7 37 13 38
rect 17 42 23 43
rect 17 38 18 42
rect 22 41 23 42
rect 35 41 37 55
rect 22 39 37 41
rect 22 38 23 39
rect 17 37 23 38
rect 11 25 13 37
rect 23 32 31 33
rect 23 28 26 32
rect 30 28 31 32
rect 23 27 31 28
rect 23 24 25 27
rect 35 25 37 39
rect 11 11 13 15
rect 23 10 25 14
rect 35 2 37 6
<< ndiffusion >>
rect 3 15 11 25
rect 13 24 18 25
rect 30 24 35 25
rect 13 22 23 24
rect 13 18 16 22
rect 20 18 23 22
rect 13 15 23 18
rect 3 12 9 15
rect 3 8 4 12
rect 8 8 9 12
rect 15 14 23 15
rect 25 14 35 24
rect 27 12 35 14
rect 3 7 9 8
rect 27 8 28 12
rect 32 8 35 12
rect 27 6 35 8
rect 37 22 45 25
rect 37 18 40 22
rect 44 18 45 22
rect 37 6 45 18
<< pdiffusion >>
rect 27 92 35 94
rect 27 88 28 92
rect 32 88 35 92
rect 27 85 35 88
rect 3 82 15 85
rect 3 78 4 82
rect 8 78 15 82
rect 3 56 15 78
rect 17 56 23 85
rect 25 56 35 85
rect 3 55 9 56
rect 30 55 35 56
rect 37 82 45 94
rect 37 78 40 82
rect 44 78 45 82
rect 37 72 45 78
rect 37 68 40 72
rect 44 68 45 72
rect 37 62 45 68
rect 37 58 40 62
rect 44 58 45 62
rect 37 55 45 58
<< metal1 >>
rect -2 96 52 100
rect -2 92 4 96
rect 8 92 16 96
rect 20 92 52 96
rect -2 88 28 92
rect 32 88 52 92
rect 3 78 4 82
rect 8 78 21 82
rect 8 42 12 73
rect 8 27 12 38
rect 17 42 21 78
rect 28 52 32 83
rect 25 48 26 52
rect 30 48 32 52
rect 17 38 18 42
rect 22 38 23 42
rect 17 22 21 38
rect 28 32 32 48
rect 25 28 26 32
rect 30 28 32 32
rect 15 18 16 22
rect 20 18 21 22
rect 28 17 32 28
rect 38 82 42 83
rect 38 78 40 82
rect 44 78 45 82
rect 38 72 42 78
rect 38 68 40 72
rect 44 68 45 72
rect 38 62 42 68
rect 38 58 40 62
rect 44 58 45 62
rect 38 22 42 58
rect 38 18 40 22
rect 44 18 45 22
rect 38 17 42 18
rect -2 8 4 12
rect 8 8 28 12
rect 32 8 52 12
rect -2 0 52 8
<< ntransistor >>
rect 11 15 13 25
rect 23 14 25 24
rect 35 6 37 25
<< ptransistor >>
rect 15 56 17 85
rect 23 56 25 85
rect 35 55 37 94
<< polycontact >>
rect 26 48 30 52
rect 8 38 12 42
rect 18 38 22 42
rect 26 28 30 32
<< ndcontact >>
rect 16 18 20 22
rect 4 8 8 12
rect 28 8 32 12
rect 40 18 44 22
<< pdcontact >>
rect 28 88 32 92
rect 4 78 8 82
rect 40 78 44 82
rect 40 68 44 72
rect 40 58 44 62
<< nsubstratencontact >>
rect 4 92 8 96
rect 16 92 20 96
<< nsubstratendiff >>
rect 3 96 21 97
rect 3 92 4 96
rect 8 92 16 96
rect 20 92 21 96
rect 3 91 21 92
<< labels >>
rlabel metal1 10 50 10 50 6 i1
rlabel metal1 25 6 25 6 6 vss
rlabel metal1 30 50 30 50 6 i0
rlabel metal1 25 94 25 94 6 vdd
rlabel metal1 40 50 40 50 6 q
<< end >>
