magic
tech scmos
timestamp 1179386914
<< checkpaint >>
rect -22 -25 158 105
<< ab >>
rect 0 0 136 80
<< pwell >>
rect -4 -7 140 36
<< nwell >>
rect -4 36 140 87
<< polysilicon >>
rect 39 70 41 74
rect 46 70 48 74
rect 53 70 55 74
rect 63 70 65 74
rect 70 70 72 74
rect 77 70 79 74
rect 87 70 89 74
rect 94 70 96 74
rect 101 70 103 74
rect 111 70 113 74
rect 118 70 120 74
rect 125 70 127 74
rect 15 62 17 67
rect 22 62 24 67
rect 29 62 31 67
rect 15 39 17 42
rect 9 38 17 39
rect 9 34 10 38
rect 14 34 17 38
rect 9 33 17 34
rect 9 22 11 33
rect 22 31 24 42
rect 29 39 31 42
rect 39 39 41 42
rect 29 38 41 39
rect 29 37 36 38
rect 35 34 36 37
rect 40 34 41 38
rect 46 39 48 42
rect 53 39 55 42
rect 63 39 65 42
rect 46 36 49 39
rect 53 37 65 39
rect 35 33 41 34
rect 21 30 27 31
rect 21 28 22 30
rect 19 26 22 28
rect 26 26 27 30
rect 39 27 41 33
rect 47 31 49 36
rect 47 30 55 31
rect 19 25 27 26
rect 31 25 43 27
rect 47 26 49 30
rect 53 26 55 30
rect 47 25 55 26
rect 19 22 21 25
rect 31 22 33 25
rect 41 22 43 25
rect 53 22 55 25
rect 63 24 65 37
rect 70 31 72 42
rect 77 39 79 42
rect 87 39 89 42
rect 77 38 90 39
rect 77 37 85 38
rect 84 34 85 37
rect 89 34 90 38
rect 84 33 90 34
rect 70 30 80 31
rect 70 29 75 30
rect 74 26 75 29
rect 79 26 80 30
rect 74 25 80 26
rect 9 6 11 10
rect 19 6 21 10
rect 31 6 33 10
rect 41 6 43 10
rect 94 23 96 42
rect 90 22 96 23
rect 90 18 91 22
rect 95 18 96 22
rect 90 17 96 18
rect 101 39 103 42
rect 111 39 113 42
rect 101 38 113 39
rect 101 34 106 38
rect 110 34 113 38
rect 101 33 113 34
rect 53 6 55 10
rect 63 9 65 12
rect 101 9 103 33
rect 118 23 120 42
rect 125 31 127 42
rect 125 30 131 31
rect 125 26 126 30
rect 130 26 131 30
rect 125 25 131 26
rect 113 22 120 23
rect 113 18 114 22
rect 118 18 120 22
rect 113 17 120 18
rect 63 7 103 9
<< ndiffusion >>
rect 58 22 63 24
rect 2 15 9 22
rect 2 11 3 15
rect 7 11 9 15
rect 2 10 9 11
rect 11 21 19 22
rect 11 17 13 21
rect 17 17 19 21
rect 11 10 19 17
rect 21 12 31 22
rect 21 10 24 12
rect 23 8 24 10
rect 28 10 31 12
rect 33 21 41 22
rect 33 17 35 21
rect 39 17 41 21
rect 33 10 41 17
rect 43 12 53 22
rect 43 10 46 12
rect 28 8 29 10
rect 23 7 29 8
rect 45 8 46 10
rect 50 10 53 12
rect 55 21 63 22
rect 55 17 57 21
rect 61 17 63 21
rect 55 12 63 17
rect 65 17 72 24
rect 65 13 67 17
rect 71 13 72 17
rect 65 12 72 13
rect 55 10 60 12
rect 50 8 51 10
rect 45 7 51 8
<< pdiffusion >>
rect 33 62 39 70
rect 8 61 15 62
rect 8 57 9 61
rect 13 57 15 61
rect 8 54 15 57
rect 8 50 9 54
rect 13 50 15 54
rect 8 49 15 50
rect 10 42 15 49
rect 17 42 22 62
rect 24 42 29 62
rect 31 61 39 62
rect 31 57 33 61
rect 37 57 39 61
rect 31 42 39 57
rect 41 42 46 70
rect 48 42 53 70
rect 55 62 63 70
rect 55 58 57 62
rect 61 58 63 62
rect 55 54 63 58
rect 55 50 57 54
rect 61 50 63 54
rect 55 42 63 50
rect 65 42 70 70
rect 72 42 77 70
rect 79 69 87 70
rect 79 65 81 69
rect 85 65 87 69
rect 79 62 87 65
rect 79 58 81 62
rect 85 58 87 62
rect 79 42 87 58
rect 89 42 94 70
rect 96 42 101 70
rect 103 62 111 70
rect 103 58 105 62
rect 109 58 111 62
rect 103 54 111 58
rect 103 50 105 54
rect 109 50 111 54
rect 103 42 111 50
rect 113 42 118 70
rect 120 42 125 70
rect 127 69 134 70
rect 127 65 129 69
rect 133 65 134 69
rect 127 62 134 65
rect 127 58 129 62
rect 133 58 134 62
rect 127 42 134 58
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect 118 78 122 82
rect 126 78 130 82
rect 134 78 138 82
rect -2 69 138 78
rect -2 68 81 69
rect 9 61 14 63
rect 13 57 14 61
rect 32 61 38 68
rect 80 65 81 68
rect 85 68 129 69
rect 85 65 86 68
rect 32 57 33 61
rect 37 57 38 61
rect 57 62 62 63
rect 61 58 62 62
rect 80 62 86 65
rect 128 65 129 68
rect 133 68 138 69
rect 133 65 134 68
rect 80 58 81 62
rect 85 58 86 62
rect 105 62 111 63
rect 109 58 111 62
rect 128 62 134 65
rect 128 58 129 62
rect 133 58 134 62
rect 9 55 14 57
rect 2 54 14 55
rect 57 54 62 58
rect 105 54 111 58
rect 2 50 9 54
rect 13 50 57 54
rect 61 50 105 54
rect 109 50 111 54
rect 2 29 6 50
rect 10 42 111 46
rect 10 38 14 42
rect 105 38 111 42
rect 10 33 14 34
rect 25 30 31 38
rect 35 34 36 38
rect 40 34 85 38
rect 89 34 98 38
rect 105 34 106 38
rect 110 34 111 38
rect 94 30 98 34
rect 2 25 14 29
rect 21 26 22 30
rect 26 26 49 30
rect 53 26 75 30
rect 79 26 87 30
rect 94 26 126 30
rect 130 26 131 30
rect 10 22 14 25
rect 81 22 87 26
rect 10 21 63 22
rect 10 17 13 21
rect 17 17 35 21
rect 39 17 57 21
rect 61 17 63 21
rect 81 18 91 22
rect 95 18 114 22
rect 118 18 119 22
rect 67 17 71 18
rect 3 15 7 16
rect -2 11 3 12
rect 67 12 71 13
rect 7 11 24 12
rect -2 8 24 11
rect 28 8 46 12
rect 50 8 138 12
rect -2 2 138 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 122 2
rect 126 -2 130 2
rect 134 -2 138 2
<< ntransistor >>
rect 9 10 11 22
rect 19 10 21 22
rect 31 10 33 22
rect 41 10 43 22
rect 53 10 55 22
rect 63 12 65 24
<< ptransistor >>
rect 15 42 17 62
rect 22 42 24 62
rect 29 42 31 62
rect 39 42 41 70
rect 46 42 48 70
rect 53 42 55 70
rect 63 42 65 70
rect 70 42 72 70
rect 77 42 79 70
rect 87 42 89 70
rect 94 42 96 70
rect 101 42 103 70
rect 111 42 113 70
rect 118 42 120 70
rect 125 42 127 70
<< polycontact >>
rect 10 34 14 38
rect 36 34 40 38
rect 22 26 26 30
rect 49 26 53 30
rect 85 34 89 38
rect 75 26 79 30
rect 91 18 95 22
rect 106 34 110 38
rect 126 26 130 30
rect 114 18 118 22
<< ndcontact >>
rect 3 11 7 15
rect 13 17 17 21
rect 24 8 28 12
rect 35 17 39 21
rect 46 8 50 12
rect 57 17 61 21
rect 67 13 71 17
<< pdcontact >>
rect 9 57 13 61
rect 9 50 13 54
rect 33 57 37 61
rect 57 58 61 62
rect 57 50 61 54
rect 81 65 85 69
rect 81 58 85 62
rect 105 58 109 62
rect 105 50 109 54
rect 129 65 133 69
rect 129 58 133 62
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
rect 90 -2 94 2
rect 98 -2 102 2
rect 106 -2 110 2
rect 114 -2 118 2
rect 122 -2 126 2
rect 130 -2 134 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
rect 90 78 94 82
rect 98 78 102 82
rect 106 78 110 82
rect 114 78 118 82
rect 122 78 126 82
rect 130 78 134 82
<< psubstratepdiff >>
rect 0 2 136 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 122 2
rect 126 -2 130 2
rect 134 -2 136 2
rect 0 -3 136 -2
<< nsubstratendiff >>
rect 0 82 136 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect 118 78 122 82
rect 126 78 130 82
rect 134 78 136 82
rect 0 77 136 78
<< labels >>
rlabel metal1 12 20 12 20 6 z
rlabel polycontact 12 36 12 36 6 c
rlabel metal1 4 40 4 40 6 z
rlabel metal1 12 56 12 56 6 z
rlabel metal1 20 20 20 20 6 z
rlabel metal1 28 20 28 20 6 z
rlabel ndcontact 36 20 36 20 6 z
rlabel metal1 36 28 36 28 6 b
rlabel metal1 28 32 28 32 6 b
rlabel metal1 28 44 28 44 6 c
rlabel metal1 36 44 36 44 6 c
rlabel metal1 20 44 20 44 6 c
rlabel metal1 20 52 20 52 6 z
rlabel metal1 28 52 28 52 6 z
rlabel metal1 36 52 36 52 6 z
rlabel metal1 44 20 44 20 6 z
rlabel metal1 52 20 52 20 6 z
rlabel ndcontact 60 20 60 20 6 z
rlabel polycontact 52 28 52 28 6 b
rlabel metal1 60 28 60 28 6 b
rlabel metal1 44 28 44 28 6 b
rlabel metal1 44 36 44 36 6 a
rlabel metal1 52 36 52 36 6 a
rlabel metal1 60 36 60 36 6 a
rlabel metal1 52 44 52 44 6 c
rlabel metal1 60 44 60 44 6 c
rlabel metal1 44 44 44 44 6 c
rlabel metal1 44 52 44 52 6 z
rlabel metal1 52 52 52 52 6 z
rlabel metal1 60 56 60 56 6 z
rlabel metal1 68 6 68 6 6 vss
rlabel metal1 84 20 84 20 6 b
rlabel polycontact 76 28 76 28 6 b
rlabel metal1 84 28 84 28 6 b
rlabel metal1 68 28 68 28 6 b
rlabel metal1 68 36 68 36 6 a
rlabel metal1 76 36 76 36 6 a
rlabel metal1 84 36 84 36 6 a
rlabel metal1 76 44 76 44 6 c
rlabel metal1 84 44 84 44 6 c
rlabel metal1 68 44 68 44 6 c
rlabel metal1 68 52 68 52 6 z
rlabel metal1 76 52 76 52 6 z
rlabel metal1 84 52 84 52 6 z
rlabel metal1 68 74 68 74 6 vdd
rlabel polycontact 92 20 92 20 6 b
rlabel metal1 100 20 100 20 6 b
rlabel metal1 108 20 108 20 6 b
rlabel metal1 100 28 100 28 6 a
rlabel metal1 108 28 108 28 6 a
rlabel metal1 92 36 92 36 6 a
rlabel metal1 100 44 100 44 6 c
rlabel metal1 108 40 108 40 6 c
rlabel metal1 92 44 92 44 6 c
rlabel metal1 92 52 92 52 6 z
rlabel metal1 100 52 100 52 6 z
rlabel metal1 108 56 108 56 6 z
rlabel polycontact 116 20 116 20 6 b
rlabel metal1 124 28 124 28 6 a
rlabel metal1 116 28 116 28 6 a
<< end >>
