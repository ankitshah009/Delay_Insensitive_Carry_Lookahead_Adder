.subckt a2_x4 i0 i1 q vdd vss
*   SPICE3 file   created from a2_x4.ext -      technology: scmos
m00 w1     i0     vdd    vdd p w=20u  l=2.3636u ad=100p     pd=30u      as=148p     ps=44.6667u
m01 vdd    i1     w1     vdd p w=20u  l=2.3636u ad=148p     pd=44.6667u as=100p     ps=30u
m02 q      w1     vdd    vdd p w=40u  l=2.3636u ad=200p     pd=50u      as=296p     ps=89.3333u
m03 vdd    w1     q      vdd p w=40u  l=2.3636u ad=296p     pd=89.3333u as=200p     ps=50u
m04 w2     i0     w1     vss n w=20u  l=2.3636u ad=100p     pd=30u      as=160p     ps=56u
m05 vss    i1     w2     vss n w=20u  l=2.3636u ad=120p     pd=38.6667u as=100p     ps=30u
m06 q      w1     vss    vss n w=20u  l=2.3636u ad=100p     pd=30u      as=120p     ps=38.6667u
m07 vss    w1     q      vss n w=20u  l=2.3636u ad=120p     pd=38.6667u as=100p     ps=30u
C0  vss    i0     0.018f
C1  vss    w1     0.156f
C2  q      i0     0.057f
C3  i1     vdd    0.154f
C4  q      w1     0.199f
C5  i0     w1     0.403f
C6  vss    w2     0.023f
C7  vss    i1     0.076f
C8  q      i1     0.485f
C9  vss    vdd    0.005f
C10 q      vdd    0.216f
C11 i1     i0     0.138f
C12 w2     w1     0.021f
C13 i1     w1     0.501f
C14 i0     vdd    0.047f
C15 vdd    w1     0.112f
C16 vss    q      0.111f
C18 q      vss    0.020f
C19 i1     vss    0.043f
C20 i0     vss    0.038f
C22 w1     vss    0.064f
.ends
