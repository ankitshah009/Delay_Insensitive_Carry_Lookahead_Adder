.subckt noa2a2a23_x4 i0 i1 i2 i3 i4 i5 nq vdd vss
*   SPICE3 file   created from noa2a2a23_x4.ext -      technology: scmos
m00 w1     i5     w2     vdd p w=40u  l=2.3636u ad=200p     pd=50u      as=248p     ps=73u
m01 w2     i4     w1     vdd p w=40u  l=2.3636u ad=248p     pd=73u      as=200p     ps=50u
m02 w3     i3     w2     vdd p w=40u  l=2.3636u ad=200p     pd=50u      as=248p     ps=73u
m03 w2     i2     w3     vdd p w=40u  l=2.3636u ad=248p     pd=73u      as=200p     ps=50u
m04 w3     i1     vdd    vdd p w=40u  l=2.3636u ad=200p     pd=50u      as=224.889p ps=65.7778u
m05 vdd    i0     w3     vdd p w=40u  l=2.3636u ad=224.889p pd=65.7778u as=200p     ps=50u
m06 nq     w4     vdd    vdd p w=40u  l=2.3636u ad=200p     pd=50u      as=224.889p ps=65.7778u
m07 vdd    w4     nq     vdd p w=40u  l=2.3636u ad=224.889p pd=65.7778u as=200p     ps=50u
m08 w4     w1     vdd    vdd p w=20u  l=2.3636u ad=160p     pd=56u      as=112.444p ps=32.8889u
m09 w5     i5     vss    vss n w=20u  l=2.3636u ad=60p      pd=26u      as=127.273p ps=42.1818u
m10 w1     i4     w5     vss n w=20u  l=2.3636u ad=120p     pd=38.6667u as=60p      ps=26u
m11 w6     i3     w1     vss n w=20u  l=2.3636u ad=60p      pd=26u      as=120p     ps=38.6667u
m12 vss    i2     w6     vss n w=20u  l=2.3636u ad=127.273p pd=42.1818u as=60p      ps=26u
m13 w7     i1     w1     vss n w=20u  l=2.3636u ad=60p      pd=26u      as=120p     ps=38.6667u
m14 vss    i0     w7     vss n w=20u  l=2.3636u ad=127.273p pd=42.1818u as=60p      ps=26u
m15 nq     w4     vss    vss n w=20u  l=2.3636u ad=124p     pd=38u      as=127.273p ps=42.1818u
m16 vss    w4     nq     vss n w=20u  l=2.3636u ad=127.273p pd=42.1818u as=124p     ps=38u
m17 w4     w1     vss    vss n w=10u  l=2.3636u ad=80p      pd=36u      as=63.6364p ps=21.0909u
C0  i3     i5     0.108f
C1  w6     w1     0.012f
C2  w3     i3     0.041f
C3  w4     i0     0.116f
C4  vdd    i4     0.017f
C5  w1     i2     0.065f
C6  nq     w3     0.024f
C7  vss    w1     0.800f
C8  w4     i2     0.002f
C9  i0     i1     0.340f
C10 w2     i3     0.017f
C11 w1     i4     0.146f
C12 vdd    w1     0.053f
C13 nq     w2     0.005f
C14 vss    w4     0.074f
C15 w2     i5     0.017f
C16 i0     i3     0.041f
C17 i1     i2     0.104f
C18 w7     vss    0.014f
C19 w3     w2     0.151f
C20 vss    i1     0.017f
C21 vdd    w4     0.072f
C22 nq     i0     0.074f
C23 i1     i4     0.042f
C24 i2     i3     0.351f
C25 w5     vss    0.014f
C26 w3     i0     0.019f
C27 vdd    i1     0.020f
C28 vss    i3     0.017f
C29 w1     w4     0.263f
C30 i3     i4     0.343f
C31 i2     i5     0.065f
C32 w7     w1     0.012f
C33 vss    nq     0.036f
C34 vss    i5     0.017f
C35 vdd    i3     0.012f
C36 w1     i1     0.047f
C37 w3     i2     0.039f
C38 i4     i5     0.367f
C39 nq     vdd    0.231f
C40 w5     w1     0.012f
C41 w1     i3     0.077f
C42 w4     i1     0.051f
C43 vdd    i5     0.012f
C44 w2     i2     0.029f
C45 w3     i4     0.025f
C46 vdd    w3     0.262f
C47 nq     w1     0.079f
C48 i0     i2     0.062f
C49 w2     i4     0.086f
C50 w1     i5     0.306f
C51 vss    i0     0.017f
C52 w3     w1     0.010f
C53 vdd    w2     0.413f
C54 nq     w4     0.120f
C55 i1     i3     0.063f
C56 w6     vss    0.014f
C57 w1     w2     0.108f
C58 vss    i2     0.017f
C59 vdd    i0     0.016f
C60 nq     i1     0.043f
C61 w3     w4     0.004f
C62 i2     i4     0.108f
C63 vdd    i2     0.012f
C64 vss    i4     0.017f
C65 w3     i1     0.043f
C66 w1     i0     0.056f
C68 nq     vss    0.015f
C70 w3     vss    0.003f
C71 w1     vss    0.044f
C72 w4     vss    0.060f
C73 i0     vss    0.030f
C74 i1     vss    0.032f
C75 i2     vss    0.032f
C76 i3     vss    0.033f
C77 i4     vss    0.034f
C78 i5     vss    0.034f
.ends
