magic
tech scmos
timestamp 1179387419
<< checkpaint >>
rect -22 -22 174 94
<< ab >>
rect 0 0 152 72
<< pwell >>
rect -4 -4 156 32
<< nwell >>
rect -4 32 156 76
<< polysilicon >>
rect 9 66 11 70
rect 19 66 21 70
rect 51 66 53 70
rect 58 66 60 70
rect 68 66 70 70
rect 78 66 80 70
rect 88 66 90 70
rect 95 66 97 70
rect 111 66 113 70
rect 121 66 123 70
rect 131 66 133 70
rect 141 66 143 70
rect 35 42 41 43
rect 35 38 36 42
rect 40 38 41 42
rect 9 35 11 38
rect 19 35 21 38
rect 9 34 21 35
rect 9 30 16 34
rect 20 30 21 34
rect 35 35 41 38
rect 51 35 53 38
rect 35 33 53 35
rect 35 31 41 33
rect 9 29 21 30
rect 9 26 11 29
rect 19 26 21 29
rect 29 29 41 31
rect 29 26 31 29
rect 39 26 41 29
rect 58 26 60 38
rect 68 35 70 38
rect 78 35 80 38
rect 64 34 80 35
rect 64 30 65 34
rect 69 33 80 34
rect 88 35 90 38
rect 95 35 97 38
rect 111 35 113 38
rect 121 35 123 38
rect 131 35 133 38
rect 69 30 70 33
rect 88 32 91 35
rect 95 34 107 35
rect 95 33 102 34
rect 64 29 70 30
rect 54 25 60 26
rect 54 21 55 25
rect 59 22 60 25
rect 79 24 81 29
rect 89 26 91 32
rect 101 30 102 33
rect 106 30 107 34
rect 101 29 107 30
rect 111 34 117 35
rect 111 30 112 34
rect 116 30 117 34
rect 111 29 117 30
rect 121 34 133 35
rect 121 30 122 34
rect 126 30 133 34
rect 141 35 143 38
rect 141 34 150 35
rect 141 31 145 34
rect 121 29 133 30
rect 114 26 116 29
rect 121 26 123 29
rect 131 26 133 29
rect 138 30 145 31
rect 149 30 150 34
rect 138 29 150 30
rect 138 26 140 29
rect 59 21 70 22
rect 54 20 70 21
rect 9 7 11 12
rect 19 7 21 12
rect 29 7 31 12
rect 39 7 41 12
rect 68 4 70 20
rect 79 4 81 7
rect 89 4 91 7
rect 68 2 91 4
rect 114 3 116 8
rect 121 3 123 8
rect 131 3 133 8
rect 138 3 140 8
<< ndiffusion >>
rect 2 25 9 26
rect 2 21 3 25
rect 7 21 9 25
rect 2 18 9 21
rect 2 14 3 18
rect 7 14 9 18
rect 2 12 9 14
rect 11 17 19 26
rect 11 13 13 17
rect 17 13 19 17
rect 11 12 19 13
rect 21 25 29 26
rect 21 21 23 25
rect 27 21 29 25
rect 21 18 29 21
rect 21 14 23 18
rect 27 14 29 18
rect 21 12 29 14
rect 31 18 39 26
rect 31 14 33 18
rect 37 14 39 18
rect 31 12 39 14
rect 41 25 48 26
rect 41 21 43 25
rect 47 21 48 25
rect 41 20 48 21
rect 84 24 89 26
rect 41 12 46 20
rect 74 19 79 24
rect 72 18 79 19
rect 72 14 73 18
rect 77 14 79 18
rect 72 13 79 14
rect 74 7 79 13
rect 81 17 89 24
rect 81 13 83 17
rect 87 13 89 17
rect 81 7 89 13
rect 91 25 98 26
rect 91 21 93 25
rect 97 21 98 25
rect 91 20 98 21
rect 91 7 96 20
rect 105 8 114 26
rect 116 8 121 26
rect 123 17 131 26
rect 123 13 125 17
rect 129 13 131 17
rect 123 8 131 13
rect 133 8 138 26
rect 140 22 148 26
rect 140 18 142 22
rect 146 18 148 22
rect 140 14 148 18
rect 140 10 142 14
rect 146 10 148 14
rect 140 8 148 10
rect 105 4 107 8
rect 111 4 112 8
rect 105 3 112 4
<< pdiffusion >>
rect 2 65 9 66
rect 2 61 3 65
rect 7 61 9 65
rect 2 57 9 61
rect 2 53 3 57
rect 7 53 9 57
rect 2 38 9 53
rect 11 51 19 66
rect 11 47 13 51
rect 17 47 19 51
rect 11 44 19 47
rect 11 40 13 44
rect 17 40 19 44
rect 11 38 19 40
rect 21 65 29 66
rect 21 61 23 65
rect 27 61 29 65
rect 21 58 29 61
rect 21 54 23 58
rect 27 54 29 58
rect 21 38 29 54
rect 99 66 109 68
rect 43 65 51 66
rect 43 61 45 65
rect 49 61 51 65
rect 43 58 51 61
rect 43 54 45 58
rect 49 54 51 58
rect 43 38 51 54
rect 53 38 58 66
rect 60 43 68 66
rect 60 39 62 43
rect 66 39 68 43
rect 60 38 68 39
rect 70 58 78 66
rect 70 54 72 58
rect 76 54 78 58
rect 70 51 78 54
rect 70 47 72 51
rect 76 47 78 51
rect 70 38 78 47
rect 80 43 88 66
rect 80 39 82 43
rect 86 39 88 43
rect 80 38 88 39
rect 90 38 95 66
rect 97 62 102 66
rect 106 62 111 66
rect 97 59 111 62
rect 97 55 102 59
rect 106 55 111 59
rect 97 38 111 55
rect 113 58 121 66
rect 113 54 115 58
rect 119 54 121 58
rect 113 51 121 54
rect 113 47 115 51
rect 119 47 121 51
rect 113 38 121 47
rect 123 65 131 66
rect 123 61 125 65
rect 129 61 131 65
rect 123 58 131 61
rect 123 54 125 58
rect 129 54 131 58
rect 123 38 131 54
rect 133 58 141 66
rect 133 54 135 58
rect 139 54 141 58
rect 133 51 141 54
rect 133 47 135 51
rect 139 47 141 51
rect 133 38 141 47
rect 143 65 150 66
rect 143 61 145 65
rect 149 61 150 65
rect 143 58 150 61
rect 143 54 145 58
rect 149 54 150 58
rect 143 38 150 54
<< metal1 >>
rect -2 68 154 72
rect -2 65 34 68
rect -2 64 3 65
rect 7 64 23 65
rect 3 57 7 61
rect 22 61 23 64
rect 27 64 34 65
rect 38 66 154 68
rect 38 65 102 66
rect 38 64 45 65
rect 27 61 28 64
rect 22 58 28 61
rect 22 54 23 58
rect 27 54 28 58
rect 44 61 45 64
rect 49 64 102 65
rect 49 61 50 64
rect 44 58 50 61
rect 101 62 102 64
rect 106 65 154 66
rect 106 64 125 65
rect 106 62 107 64
rect 101 59 107 62
rect 124 61 125 64
rect 129 64 145 65
rect 129 61 130 64
rect 44 54 45 58
rect 49 54 50 58
rect 72 58 76 59
rect 101 55 102 59
rect 106 55 107 59
rect 115 58 119 59
rect 3 52 7 53
rect 13 51 17 52
rect 72 51 76 54
rect 124 58 130 61
rect 144 61 145 64
rect 149 64 154 65
rect 149 61 150 64
rect 124 54 125 58
rect 129 54 130 58
rect 135 58 140 59
rect 139 54 140 58
rect 144 58 150 61
rect 144 54 145 58
rect 149 54 150 58
rect 115 51 119 54
rect 135 51 140 54
rect 13 44 17 47
rect 2 40 13 43
rect 2 39 17 40
rect 2 25 6 39
rect 26 34 30 51
rect 46 47 72 51
rect 76 47 115 51
rect 119 47 135 51
rect 139 47 140 51
rect 46 42 50 47
rect 35 38 36 42
rect 40 38 50 42
rect 57 39 62 43
rect 66 39 82 43
rect 86 39 87 43
rect 57 38 87 39
rect 15 30 16 34
rect 20 30 65 34
rect 69 30 71 34
rect 82 26 87 38
rect 102 34 106 47
rect 146 42 150 51
rect 111 38 150 42
rect 111 34 117 38
rect 145 34 150 38
rect 111 30 112 34
rect 116 30 117 34
rect 121 30 122 34
rect 126 30 127 34
rect 73 25 98 26
rect 2 21 3 25
rect 7 21 23 25
rect 27 21 43 25
rect 47 21 55 25
rect 59 21 60 25
rect 73 21 93 25
rect 97 21 98 25
rect 3 18 7 21
rect 23 18 27 21
rect 73 18 78 21
rect 3 13 7 14
rect 12 13 13 17
rect 17 13 18 17
rect 32 14 33 18
rect 37 14 73 18
rect 77 14 78 18
rect 102 17 106 30
rect 121 26 127 30
rect 149 30 150 34
rect 145 29 150 30
rect 121 22 135 26
rect 142 22 146 23
rect 23 13 27 14
rect 82 13 83 17
rect 87 13 125 17
rect 129 13 130 17
rect 142 14 146 18
rect 12 8 18 13
rect 142 8 146 10
rect -2 4 52 8
rect 56 4 60 8
rect 64 4 107 8
rect 111 4 154 8
rect -2 0 154 4
<< ntransistor >>
rect 9 12 11 26
rect 19 12 21 26
rect 29 12 31 26
rect 39 12 41 26
rect 79 7 81 24
rect 89 7 91 26
rect 114 8 116 26
rect 121 8 123 26
rect 131 8 133 26
rect 138 8 140 26
<< ptransistor >>
rect 9 38 11 66
rect 19 38 21 66
rect 51 38 53 66
rect 58 38 60 66
rect 68 38 70 66
rect 78 38 80 66
rect 88 38 90 66
rect 95 38 97 66
rect 111 38 113 66
rect 121 38 123 66
rect 131 38 133 66
rect 141 38 143 66
<< polycontact >>
rect 36 38 40 42
rect 16 30 20 34
rect 65 30 69 34
rect 55 21 59 25
rect 102 30 106 34
rect 112 30 116 34
rect 122 30 126 34
rect 145 30 149 34
<< ndcontact >>
rect 3 21 7 25
rect 3 14 7 18
rect 13 13 17 17
rect 23 21 27 25
rect 23 14 27 18
rect 33 14 37 18
rect 43 21 47 25
rect 73 14 77 18
rect 83 13 87 17
rect 93 21 97 25
rect 125 13 129 17
rect 142 18 146 22
rect 142 10 146 14
rect 107 4 111 8
<< pdcontact >>
rect 3 61 7 65
rect 3 53 7 57
rect 13 47 17 51
rect 13 40 17 44
rect 23 61 27 65
rect 23 54 27 58
rect 45 61 49 65
rect 45 54 49 58
rect 62 39 66 43
rect 72 54 76 58
rect 72 47 76 51
rect 82 39 86 43
rect 102 62 106 66
rect 102 55 106 59
rect 115 54 119 58
rect 115 47 119 51
rect 125 61 129 65
rect 125 54 129 58
rect 135 54 139 58
rect 135 47 139 51
rect 145 61 149 65
rect 145 54 149 58
<< psubstratepcontact >>
rect 52 4 56 8
rect 60 4 64 8
<< nsubstratencontact >>
rect 34 64 38 68
<< psubstratepdiff >>
rect 51 8 65 9
rect 51 4 52 8
rect 56 4 60 8
rect 64 4 65 8
rect 51 3 65 4
<< nsubstratendiff >>
rect 33 68 39 69
rect 33 64 34 68
rect 38 64 39 68
rect 33 47 39 64
<< labels >>
rlabel polysilicon 38 36 38 36 6 an
rlabel polycontact 57 23 57 23 6 bn
rlabel polycontact 104 32 104 32 6 an
rlabel metal1 25 19 25 19 6 bn
rlabel metal1 5 19 5 19 6 bn
rlabel metal1 20 32 20 32 6 b
rlabel metal1 15 45 15 45 6 bn
rlabel ndcontact 36 16 36 16 6 z
rlabel metal1 44 16 44 16 6 z
rlabel metal1 52 16 52 16 6 z
rlabel metal1 36 32 36 32 6 b
rlabel metal1 44 32 44 32 6 b
rlabel metal1 52 32 52 32 6 b
rlabel metal1 28 40 28 40 6 b
rlabel metal1 42 40 42 40 6 an
rlabel metal1 76 4 76 4 6 vss
rlabel metal1 68 16 68 16 6 z
rlabel metal1 60 16 60 16 6 z
rlabel metal1 31 23 31 23 6 bn
rlabel metal1 76 24 76 24 6 z
rlabel polycontact 68 32 68 32 6 b
rlabel metal1 84 32 84 32 6 z
rlabel metal1 60 32 60 32 6 b
rlabel metal1 60 40 60 40 6 z
rlabel metal1 68 40 68 40 6 z
rlabel metal1 76 40 76 40 6 z
rlabel metal1 74 53 74 53 6 an
rlabel metal1 76 68 76 68 6 vdd
rlabel metal1 92 24 92 24 6 z
rlabel metal1 116 40 116 40 6 a1
rlabel polycontact 104 32 104 32 6 an
rlabel metal1 117 53 117 53 6 an
rlabel metal1 106 15 106 15 6 an
rlabel metal1 132 24 132 24 6 a2
rlabel metal1 124 28 124 28 6 a2
rlabel metal1 124 40 124 40 6 a1
rlabel metal1 148 40 148 40 6 a1
rlabel metal1 132 40 132 40 6 a1
rlabel metal1 140 40 140 40 6 a1
rlabel metal1 93 49 93 49 6 an
rlabel metal1 137 53 137 53 6 an
<< end >>
