magic
tech scmos
timestamp 1179386304
<< checkpaint >>
rect -22 -25 54 105
<< ab >>
rect 0 0 32 80
<< pwell >>
rect -4 -7 36 36
<< nwell >>
rect -4 36 36 87
<< polysilicon >>
rect 9 70 11 74
rect 19 70 21 74
rect 9 39 11 46
rect 19 43 21 46
rect 19 42 30 43
rect 9 38 15 39
rect 9 34 10 38
rect 14 34 15 38
rect 9 33 15 34
rect 19 38 25 42
rect 29 38 30 42
rect 19 37 30 38
rect 12 30 14 33
rect 19 30 21 37
rect 12 6 14 10
rect 19 6 21 10
<< ndiffusion >>
rect 7 22 12 30
rect 5 21 12 22
rect 5 17 6 21
rect 10 17 12 21
rect 5 16 12 17
rect 7 10 12 16
rect 14 10 19 30
rect 21 22 30 30
rect 21 18 25 22
rect 29 18 30 22
rect 21 15 30 18
rect 21 11 25 15
rect 29 11 30 15
rect 21 10 30 11
<< pdiffusion >>
rect 2 69 9 70
rect 2 65 3 69
rect 7 65 9 69
rect 2 62 9 65
rect 2 58 3 62
rect 7 58 9 62
rect 2 46 9 58
rect 11 62 19 70
rect 11 58 13 62
rect 17 58 19 62
rect 11 55 19 58
rect 11 51 13 55
rect 17 51 19 55
rect 11 46 19 51
rect 21 69 29 70
rect 21 65 23 69
rect 27 65 29 69
rect 21 62 29 65
rect 21 58 23 62
rect 27 58 29 62
rect 21 46 29 58
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect -2 69 34 78
rect -2 68 3 69
rect 2 65 3 68
rect 7 68 23 69
rect 7 65 8 68
rect 2 62 8 65
rect 22 65 23 68
rect 27 68 34 69
rect 27 65 28 68
rect 2 58 3 62
rect 7 58 8 62
rect 13 62 17 63
rect 22 62 28 65
rect 22 58 23 62
rect 27 58 28 62
rect 13 55 17 58
rect 2 51 13 55
rect 2 50 17 51
rect 2 49 14 50
rect 2 17 6 49
rect 18 42 30 47
rect 18 41 25 42
rect 10 38 14 39
rect 29 38 30 42
rect 25 37 30 38
rect 10 31 14 34
rect 26 33 30 37
rect 10 25 22 31
rect 25 22 29 23
rect 10 17 11 21
rect 25 15 29 18
rect -2 11 25 12
rect 29 11 34 12
rect -2 2 34 11
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
<< ntransistor >>
rect 12 10 14 30
rect 19 10 21 30
<< ptransistor >>
rect 9 46 11 70
rect 19 46 21 70
<< polycontact >>
rect 10 34 14 38
rect 25 38 29 42
<< ndcontact >>
rect 6 17 10 21
rect 25 18 29 22
rect 25 11 29 15
<< pdcontact >>
rect 3 65 7 69
rect 3 58 7 62
rect 13 58 17 62
rect 13 51 17 55
rect 23 65 27 69
rect 23 58 27 62
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
<< psubstratepdiff >>
rect 0 2 32 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 32 2
rect 0 -3 32 -2
<< nsubstratendiff >>
rect 0 82 32 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 32 82
rect 0 77 32 78
<< labels >>
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 32 12 32 6 b
rlabel metal1 12 52 12 52 6 z
rlabel metal1 16 6 16 6 6 vss
rlabel metal1 20 28 20 28 6 b
rlabel metal1 20 44 20 44 6 a
rlabel metal1 16 74 16 74 6 vdd
rlabel polycontact 28 40 28 40 6 a
<< end >>
