magic
tech scmos
timestamp 1179387299
<< checkpaint >>
rect -22 -25 118 105
<< ab >>
rect 0 0 96 80
<< pwell >>
rect -4 -7 100 36
<< nwell >>
rect -4 36 100 87
<< polysilicon >>
rect 33 70 35 74
rect 40 70 42 74
rect 47 70 49 74
rect 54 70 56 74
rect 64 70 66 74
rect 71 70 73 74
rect 78 70 80 74
rect 85 70 87 74
rect 9 61 11 65
rect 19 63 21 68
rect 9 39 11 42
rect 19 39 21 42
rect 33 39 35 42
rect 9 38 21 39
rect 9 34 16 38
rect 20 34 21 38
rect 9 33 21 34
rect 28 38 35 39
rect 28 34 29 38
rect 33 36 35 38
rect 33 34 34 36
rect 28 33 34 34
rect 9 30 11 33
rect 28 22 30 33
rect 40 32 42 42
rect 47 39 49 42
rect 54 39 56 42
rect 64 39 66 42
rect 47 36 50 39
rect 54 38 66 39
rect 54 37 59 38
rect 38 31 44 32
rect 38 27 39 31
rect 43 27 44 31
rect 38 26 44 27
rect 48 31 50 36
rect 58 34 59 37
rect 63 37 66 38
rect 63 34 64 37
rect 58 33 64 34
rect 48 30 54 31
rect 48 26 49 30
rect 53 26 54 30
rect 38 22 40 26
rect 48 25 54 26
rect 50 22 52 25
rect 60 22 62 33
rect 71 31 73 42
rect 78 33 80 42
rect 85 39 87 42
rect 85 38 94 39
rect 85 37 89 38
rect 88 34 89 37
rect 93 34 94 38
rect 88 33 94 34
rect 78 32 84 33
rect 68 30 74 31
rect 68 26 69 30
rect 73 26 74 30
rect 78 28 79 32
rect 83 28 84 32
rect 78 27 84 28
rect 68 25 74 26
rect 9 6 11 10
rect 28 9 30 14
rect 38 9 40 14
rect 50 9 52 14
rect 60 9 62 14
<< ndiffusion >>
rect 2 29 9 30
rect 2 25 3 29
rect 7 25 9 29
rect 2 22 9 25
rect 2 18 3 22
rect 7 18 9 22
rect 2 17 9 18
rect 4 10 9 17
rect 11 22 26 30
rect 11 21 28 22
rect 11 17 13 21
rect 17 17 28 21
rect 11 14 28 17
rect 30 21 38 22
rect 30 17 32 21
rect 36 17 38 21
rect 30 14 38 17
rect 40 14 50 22
rect 52 21 60 22
rect 52 17 54 21
rect 58 17 60 21
rect 52 14 60 17
rect 62 14 71 22
rect 11 12 26 14
rect 11 10 14 12
rect 13 8 14 10
rect 18 8 21 12
rect 25 8 26 12
rect 42 12 48 14
rect 13 7 26 8
rect 42 8 43 12
rect 47 8 48 12
rect 64 12 71 14
rect 42 7 48 8
rect 64 8 65 12
rect 69 8 71 12
rect 64 7 71 8
<< pdiffusion >>
rect 23 69 33 70
rect 23 65 25 69
rect 29 65 33 69
rect 23 63 33 65
rect 14 61 19 63
rect 2 60 9 61
rect 2 56 3 60
rect 7 56 9 60
rect 2 53 9 56
rect 2 49 3 53
rect 7 49 9 53
rect 2 42 9 49
rect 11 54 19 61
rect 11 50 13 54
rect 17 50 19 54
rect 11 47 19 50
rect 11 43 13 47
rect 17 43 19 47
rect 11 42 19 43
rect 21 42 33 63
rect 35 42 40 70
rect 42 42 47 70
rect 49 42 54 70
rect 56 62 64 70
rect 56 58 58 62
rect 62 58 64 62
rect 56 42 64 58
rect 66 42 71 70
rect 73 42 78 70
rect 80 42 85 70
rect 87 69 94 70
rect 87 65 89 69
rect 93 65 94 69
rect 87 62 94 65
rect 87 58 89 62
rect 93 58 94 62
rect 87 42 94 58
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect -2 69 98 78
rect -2 68 25 69
rect 2 60 8 68
rect 24 65 25 68
rect 29 68 89 69
rect 29 65 30 68
rect 88 65 89 68
rect 93 68 98 69
rect 93 65 94 68
rect 2 56 3 60
rect 7 56 8 60
rect 2 53 8 56
rect 21 58 58 62
rect 62 58 63 62
rect 2 49 3 53
rect 7 49 8 53
rect 13 54 17 55
rect 13 47 17 50
rect 2 43 13 46
rect 2 42 17 43
rect 2 30 6 42
rect 21 38 25 58
rect 74 54 78 63
rect 88 62 94 65
rect 88 58 89 62
rect 93 58 94 62
rect 15 34 16 38
rect 20 34 25 38
rect 2 29 15 30
rect 2 25 3 29
rect 7 26 15 29
rect 2 22 7 25
rect 2 18 3 22
rect 2 17 7 18
rect 13 21 17 22
rect 21 21 25 34
rect 29 50 94 54
rect 29 38 33 50
rect 29 33 33 34
rect 39 42 79 46
rect 39 31 43 42
rect 73 38 79 42
rect 89 38 94 50
rect 49 34 59 38
rect 63 34 64 38
rect 73 34 83 38
rect 79 32 83 34
rect 93 34 94 38
rect 89 33 94 34
rect 39 26 43 27
rect 48 26 49 30
rect 53 26 69 30
rect 73 26 74 30
rect 79 27 83 28
rect 21 17 32 21
rect 36 17 54 21
rect 58 17 59 21
rect 66 17 70 26
rect 13 12 17 17
rect -2 8 14 12
rect 18 8 21 12
rect 25 8 43 12
rect 47 8 65 12
rect 69 8 98 12
rect -2 2 98 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
<< ntransistor >>
rect 9 10 11 30
rect 28 14 30 22
rect 38 14 40 22
rect 50 14 52 22
rect 60 14 62 22
<< ptransistor >>
rect 9 42 11 61
rect 19 42 21 63
rect 33 42 35 70
rect 40 42 42 70
rect 47 42 49 70
rect 54 42 56 70
rect 64 42 66 70
rect 71 42 73 70
rect 78 42 80 70
rect 85 42 87 70
<< polycontact >>
rect 16 34 20 38
rect 29 34 33 38
rect 39 27 43 31
rect 59 34 63 38
rect 49 26 53 30
rect 89 34 93 38
rect 69 26 73 30
rect 79 28 83 32
<< ndcontact >>
rect 3 25 7 29
rect 3 18 7 22
rect 13 17 17 21
rect 32 17 36 21
rect 54 17 58 21
rect 14 8 18 12
rect 21 8 25 12
rect 43 8 47 12
rect 65 8 69 12
<< pdcontact >>
rect 25 65 29 69
rect 3 56 7 60
rect 3 49 7 53
rect 13 50 17 54
rect 13 43 17 47
rect 58 58 62 62
rect 89 65 93 69
rect 89 58 93 62
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
rect 90 -2 94 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
rect 90 78 94 82
<< psubstratepdiff >>
rect 0 2 96 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 96 2
rect 0 -3 96 -2
<< nsubstratendiff >>
rect 0 82 96 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 96 82
rect 0 77 96 78
<< labels >>
rlabel polysilicon 15 36 15 36 6 zn
rlabel ndcontact 4 28 4 28 6 z
rlabel metal1 12 28 12 28 6 z
rlabel metal1 12 44 12 44 6 z
rlabel metal1 20 36 20 36 6 zn
rlabel metal1 48 6 48 6 6 vss
rlabel polycontact 52 28 52 28 6 c
rlabel metal1 44 44 44 44 6 b
rlabel metal1 52 36 52 36 6 d
rlabel metal1 52 44 52 44 6 b
rlabel metal1 44 52 44 52 6 a
rlabel metal1 52 52 52 52 6 a
rlabel metal1 36 52 36 52 6 a
rlabel metal1 48 74 48 74 6 vdd
rlabel metal1 60 28 60 28 6 c
rlabel metal1 40 19 40 19 6 zn
rlabel metal1 68 20 68 20 6 c
rlabel metal1 68 24 68 24 6 c
rlabel polycontact 60 36 60 36 6 d
rlabel metal1 60 44 60 44 6 b
rlabel metal1 68 44 68 44 6 b
rlabel metal1 76 40 76 40 6 b
rlabel metal1 68 52 68 52 6 a
rlabel metal1 60 52 60 52 6 a
rlabel metal1 42 60 42 60 6 zn
rlabel metal1 76 56 76 56 6 a
rlabel metal1 92 40 92 40 6 a
rlabel metal1 84 52 84 52 6 a
<< end >>
