magic
tech scmos
timestamp 1179386961
<< checkpaint >>
rect -22 -25 70 105
<< ab >>
rect 0 0 48 80
<< pwell >>
rect -4 -7 52 36
<< nwell >>
rect -4 36 52 87
<< polysilicon >>
rect 30 68 32 73
rect 37 68 39 73
rect 10 61 12 65
rect 20 61 22 65
rect 10 47 12 52
rect 9 46 15 47
rect 9 42 10 46
rect 14 42 15 46
rect 9 41 15 42
rect 9 23 11 41
rect 20 32 22 52
rect 30 38 32 52
rect 37 49 39 52
rect 37 48 46 49
rect 37 44 41 48
rect 45 44 46 48
rect 37 43 46 44
rect 16 31 22 32
rect 16 27 17 31
rect 21 27 22 31
rect 16 26 22 27
rect 26 37 33 38
rect 26 33 28 37
rect 32 33 33 37
rect 26 32 33 33
rect 16 23 18 26
rect 26 23 28 32
rect 37 29 39 43
rect 37 15 39 19
rect 9 8 11 13
rect 16 8 18 13
rect 26 8 28 13
<< ndiffusion >>
rect 30 23 37 29
rect 2 22 9 23
rect 2 18 3 22
rect 7 18 9 22
rect 2 17 9 18
rect 4 13 9 17
rect 11 13 16 23
rect 18 21 26 23
rect 18 17 20 21
rect 24 17 26 21
rect 18 13 26 17
rect 28 19 37 23
rect 39 25 44 29
rect 39 24 46 25
rect 39 20 41 24
rect 45 20 46 24
rect 39 19 46 20
rect 28 13 35 19
rect 30 12 36 13
rect 30 8 31 12
rect 35 8 36 12
rect 30 7 36 8
<< pdiffusion >>
rect 2 72 8 73
rect 2 68 3 72
rect 7 68 8 72
rect 2 61 8 68
rect 22 72 28 73
rect 22 68 23 72
rect 27 68 28 72
rect 22 67 30 68
rect 24 61 30 67
rect 2 52 10 61
rect 12 60 20 61
rect 12 56 14 60
rect 18 56 20 60
rect 12 52 20 56
rect 22 52 30 61
rect 32 52 37 68
rect 39 64 44 68
rect 39 63 46 64
rect 39 59 41 63
rect 45 59 46 63
rect 39 58 46 59
rect 39 52 44 58
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect -2 72 50 78
rect -2 68 3 72
rect 7 68 23 72
rect 27 68 50 72
rect 2 60 41 63
rect 2 57 14 60
rect 2 23 6 57
rect 13 56 14 57
rect 18 59 41 60
rect 45 59 46 63
rect 18 57 22 59
rect 18 56 19 57
rect 26 47 30 55
rect 34 49 46 55
rect 10 46 30 47
rect 14 43 30 46
rect 41 48 46 49
rect 45 44 46 48
rect 41 43 46 44
rect 14 42 22 43
rect 10 41 22 42
rect 42 41 46 43
rect 26 37 38 39
rect 26 33 28 37
rect 32 33 38 37
rect 10 27 17 31
rect 21 27 22 31
rect 10 25 22 27
rect 34 25 38 33
rect 2 22 7 23
rect 2 18 3 22
rect 2 17 7 18
rect 10 17 14 25
rect 41 24 45 25
rect 19 17 20 21
rect 24 20 41 21
rect 24 17 45 20
rect -2 8 31 12
rect 35 8 50 12
rect -2 2 50 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
<< ntransistor >>
rect 9 13 11 23
rect 16 13 18 23
rect 26 13 28 23
rect 37 19 39 29
<< ptransistor >>
rect 10 52 12 61
rect 20 52 22 61
rect 30 52 32 68
rect 37 52 39 68
<< polycontact >>
rect 10 42 14 46
rect 41 44 45 48
rect 17 27 21 31
rect 28 33 32 37
<< ndcontact >>
rect 3 18 7 22
rect 20 17 24 21
rect 41 20 45 24
rect 31 8 35 12
<< pdcontact >>
rect 3 68 7 72
rect 23 68 27 72
rect 14 56 18 60
rect 41 59 45 63
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
<< psubstratepdiff >>
rect 0 2 48 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 48 2
rect 0 -3 48 -2
<< nsubstratendiff >>
rect 0 82 48 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 48 82
rect 0 77 48 78
<< labels >>
rlabel metal1 4 40 4 40 6 z
rlabel metal1 12 24 12 24 6 b
rlabel polycontact 12 44 12 44 6 c
rlabel metal1 12 60 12 60 6 z
rlabel metal1 24 6 24 6 6 vss
rlabel polycontact 20 28 20 28 6 b
rlabel metal1 20 44 20 44 6 c
rlabel metal1 20 60 20 60 6 z
rlabel metal1 24 74 24 74 6 vdd
rlabel metal1 36 32 36 32 6 a1
rlabel metal1 28 36 28 36 6 a1
rlabel metal1 36 52 36 52 6 a2
rlabel metal1 28 52 28 52 6 c
rlabel metal1 32 19 32 19 6 n1
rlabel metal1 44 48 44 48 6 a2
<< end >>
