magic
tech scmos
timestamp 1179387502
<< checkpaint >>
rect -22 -25 126 105
<< ab >>
rect 0 0 104 80
<< pwell >>
rect -4 -7 108 36
<< nwell >>
rect -4 36 108 87
<< polysilicon >>
rect 9 70 11 74
rect 16 70 18 74
rect 26 70 28 74
rect 33 70 35 74
rect 43 70 45 74
rect 53 70 55 74
rect 63 68 65 73
rect 73 68 75 73
rect 83 61 85 66
rect 93 61 95 65
rect 9 23 11 42
rect 16 39 18 42
rect 26 39 28 42
rect 16 38 28 39
rect 16 34 23 38
rect 27 34 28 38
rect 16 33 28 34
rect 23 30 25 33
rect 33 30 35 42
rect 43 39 45 50
rect 53 47 55 50
rect 63 47 65 50
rect 73 47 75 50
rect 53 45 65 47
rect 43 38 57 39
rect 43 34 50 38
rect 54 34 57 38
rect 43 33 57 34
rect 63 35 65 45
rect 69 46 75 47
rect 69 42 70 46
rect 74 42 75 46
rect 69 41 75 42
rect 83 35 85 42
rect 93 39 95 42
rect 93 38 102 39
rect 93 35 97 38
rect 63 34 97 35
rect 101 34 102 38
rect 63 33 102 34
rect 43 30 45 33
rect 55 30 57 33
rect 78 30 80 33
rect 5 22 11 23
rect 5 18 6 22
rect 10 18 11 22
rect 5 17 11 18
rect 55 19 57 24
rect 63 21 69 22
rect 43 12 45 17
rect 23 6 25 11
rect 33 8 35 11
rect 63 17 64 21
rect 68 17 69 21
rect 63 16 69 17
rect 63 8 65 16
rect 33 6 65 8
rect 78 6 80 11
<< ndiffusion >>
rect 18 23 23 30
rect 16 22 23 23
rect 16 18 17 22
rect 21 18 23 22
rect 16 17 23 18
rect 18 11 23 17
rect 25 29 33 30
rect 25 25 27 29
rect 31 25 33 29
rect 25 11 33 25
rect 35 29 43 30
rect 35 25 37 29
rect 41 25 43 29
rect 35 17 43 25
rect 45 24 55 30
rect 57 29 64 30
rect 57 25 59 29
rect 63 25 64 29
rect 57 24 64 25
rect 71 29 78 30
rect 71 25 72 29
rect 76 25 78 29
rect 45 17 53 24
rect 71 22 78 25
rect 35 11 40 17
rect 47 15 53 17
rect 47 11 48 15
rect 52 11 53 15
rect 47 10 53 11
rect 71 18 72 22
rect 76 18 78 22
rect 71 17 78 18
rect 73 11 78 17
rect 80 23 88 30
rect 80 19 82 23
rect 86 19 88 23
rect 80 16 88 19
rect 80 12 82 16
rect 86 12 88 16
rect 80 11 88 12
<< pdiffusion >>
rect 2 69 9 70
rect 2 65 3 69
rect 7 65 9 69
rect 2 62 9 65
rect 2 58 3 62
rect 7 58 9 62
rect 2 42 9 58
rect 11 42 16 70
rect 18 62 26 70
rect 18 58 20 62
rect 24 58 26 62
rect 18 47 26 58
rect 18 43 20 47
rect 24 43 26 47
rect 18 42 26 43
rect 28 42 33 70
rect 35 69 43 70
rect 35 65 37 69
rect 41 65 43 69
rect 35 50 43 65
rect 45 55 53 70
rect 45 51 47 55
rect 51 51 53 55
rect 45 50 53 51
rect 55 68 60 70
rect 55 62 63 68
rect 55 58 57 62
rect 61 58 63 62
rect 55 50 63 58
rect 65 62 73 68
rect 65 58 67 62
rect 71 58 73 62
rect 65 55 73 58
rect 65 51 67 55
rect 71 51 73 55
rect 65 50 73 51
rect 75 61 81 68
rect 75 60 83 61
rect 75 56 77 60
rect 81 56 83 60
rect 75 50 83 56
rect 35 42 41 50
rect 77 42 83 50
rect 85 54 93 61
rect 85 50 87 54
rect 91 50 93 54
rect 85 47 93 50
rect 85 43 87 47
rect 91 43 93 47
rect 85 42 93 43
rect 95 60 102 61
rect 95 56 97 60
rect 101 56 102 60
rect 95 53 102 56
rect 95 49 97 53
rect 101 49 102 53
rect 95 42 102 49
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect -2 69 106 78
rect -2 68 3 69
rect 2 65 3 68
rect 7 68 37 69
rect 7 65 8 68
rect 36 65 37 68
rect 41 68 106 69
rect 41 65 42 68
rect 2 62 8 65
rect 67 62 71 63
rect 2 58 3 62
rect 7 58 8 62
rect 18 58 20 62
rect 24 58 57 62
rect 61 58 63 62
rect 18 48 22 58
rect 67 55 71 58
rect 77 60 81 68
rect 77 55 81 56
rect 97 60 101 68
rect 46 54 47 55
rect 36 51 47 54
rect 51 54 52 55
rect 51 51 67 54
rect 36 50 71 51
rect 87 54 91 55
rect 18 47 24 48
rect 10 43 20 47
rect 10 42 24 43
rect 10 30 14 42
rect 36 38 40 50
rect 87 47 91 50
rect 97 53 101 56
rect 97 48 101 49
rect 22 34 23 38
rect 27 34 40 38
rect 49 42 70 46
rect 74 42 75 46
rect 49 38 55 42
rect 87 38 91 43
rect 49 34 50 38
rect 54 34 55 38
rect 72 34 91 38
rect 97 38 102 39
rect 101 34 102 38
rect 36 30 40 34
rect 10 29 32 30
rect 10 26 27 29
rect 26 25 27 26
rect 31 25 32 29
rect 36 29 64 30
rect 36 25 37 29
rect 41 26 59 29
rect 41 25 42 26
rect 58 25 59 26
rect 63 25 64 29
rect 72 29 76 34
rect 72 22 76 25
rect 5 18 6 22
rect 10 18 17 22
rect 21 21 72 22
rect 21 18 64 21
rect 63 17 64 18
rect 68 18 72 21
rect 68 17 76 18
rect 82 23 86 24
rect 97 23 102 34
rect 82 16 86 19
rect 90 17 102 23
rect 47 12 48 15
rect -2 11 48 12
rect 52 12 53 15
rect 52 11 106 12
rect -2 2 106 11
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
<< ntransistor >>
rect 23 11 25 30
rect 33 11 35 30
rect 43 17 45 30
rect 55 24 57 30
rect 78 11 80 30
<< ptransistor >>
rect 9 42 11 70
rect 16 42 18 70
rect 26 42 28 70
rect 33 42 35 70
rect 43 50 45 70
rect 53 50 55 70
rect 63 50 65 68
rect 73 50 75 68
rect 83 42 85 61
rect 93 42 95 61
<< polycontact >>
rect 23 34 27 38
rect 50 34 54 38
rect 70 42 74 46
rect 97 34 101 38
rect 6 18 10 22
rect 64 17 68 21
<< ndcontact >>
rect 17 18 21 22
rect 27 25 31 29
rect 37 25 41 29
rect 59 25 63 29
rect 72 25 76 29
rect 48 11 52 15
rect 72 18 76 22
rect 82 19 86 23
rect 82 12 86 16
<< pdcontact >>
rect 3 65 7 69
rect 3 58 7 62
rect 20 58 24 62
rect 20 43 24 47
rect 37 65 41 69
rect 47 51 51 55
rect 57 58 61 62
rect 67 58 71 62
rect 67 51 71 55
rect 77 56 81 60
rect 87 50 91 54
rect 87 43 91 47
rect 97 56 101 60
rect 97 49 101 53
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
rect 90 -2 94 2
rect 98 -2 102 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
rect 90 78 94 82
rect 98 78 102 82
<< psubstratepdiff >>
rect 0 2 104 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 104 2
rect 0 -3 104 -2
<< nsubstratendiff >>
rect 0 82 104 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 104 82
rect 0 77 104 78
<< labels >>
rlabel polycontact 8 20 8 20 6 bn
rlabel polysilicon 22 36 22 36 6 an
rlabel polycontact 66 19 66 19 6 bn
rlabel metal1 12 40 12 40 6 z
rlabel metal1 20 28 20 28 6 z
rlabel ndcontact 28 28 28 28 6 z
rlabel metal1 31 36 31 36 6 an
rlabel metal1 20 48 20 48 6 z
rlabel metal1 28 60 28 60 6 z
rlabel metal1 36 60 36 60 6 z
rlabel metal1 52 6 52 6 6 vss
rlabel metal1 52 40 52 40 6 a
rlabel metal1 60 44 60 44 6 a
rlabel metal1 44 60 44 60 6 z
rlabel metal1 52 60 52 60 6 z
rlabel pdcontact 60 60 60 60 6 z
rlabel metal1 52 74 52 74 6 vdd
rlabel metal1 40 20 40 20 6 bn
rlabel metal1 50 28 50 28 6 an
rlabel ndcontact 74 27 74 27 6 bn
rlabel metal1 68 44 68 44 6 a
rlabel metal1 69 56 69 56 6 an
rlabel metal1 53 52 53 52 6 an
rlabel metal1 92 20 92 20 6 b
rlabel metal1 100 28 100 28 6 b
rlabel pdcontact 89 44 89 44 6 bn
<< end >>
