magic
tech scmos
timestamp 1179385954
<< checkpaint >>
rect -22 -25 54 105
<< ab >>
rect 0 0 32 80
<< pwell >>
rect -4 -7 36 36
<< nwell >>
rect -4 36 36 87
<< polysilicon >>
rect 10 70 12 74
rect 20 61 22 65
rect 10 39 12 42
rect 20 39 22 42
rect 9 38 22 39
rect 9 34 17 38
rect 21 34 22 38
rect 9 33 22 34
rect 9 30 11 33
rect 9 13 11 18
<< ndiffusion >>
rect 2 29 9 30
rect 2 25 3 29
rect 7 25 9 29
rect 2 24 9 25
rect 4 18 9 24
rect 11 23 19 30
rect 11 19 13 23
rect 17 19 19 23
rect 11 18 19 19
<< pdiffusion >>
rect 2 69 10 70
rect 2 65 4 69
rect 8 65 10 69
rect 2 62 10 65
rect 2 58 4 62
rect 8 58 10 62
rect 2 42 10 58
rect 12 61 17 70
rect 12 54 20 61
rect 12 50 14 54
rect 18 50 20 54
rect 12 47 20 50
rect 12 43 14 47
rect 18 43 20 47
rect 12 42 20 43
rect 22 60 30 61
rect 22 56 24 60
rect 28 56 30 60
rect 22 53 30 56
rect 22 49 24 53
rect 28 49 30 53
rect 22 42 30 49
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect -2 69 34 78
rect -2 68 4 69
rect 3 65 4 68
rect 8 68 34 69
rect 8 65 9 68
rect 3 62 9 65
rect 3 58 4 62
rect 8 58 9 62
rect 23 60 29 68
rect 23 56 24 60
rect 28 56 29 60
rect 14 54 18 55
rect 14 47 18 50
rect 23 53 29 56
rect 23 49 24 53
rect 28 49 29 53
rect 2 43 14 47
rect 18 43 23 46
rect 2 42 23 43
rect 2 30 6 42
rect 16 34 17 38
rect 21 34 30 38
rect 2 29 7 30
rect 2 25 3 29
rect 26 25 30 34
rect 2 24 7 25
rect 13 23 17 24
rect 13 12 17 19
rect -2 2 34 12
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
<< ntransistor >>
rect 9 18 11 30
<< ptransistor >>
rect 10 42 12 70
rect 20 42 22 61
<< polycontact >>
rect 17 34 21 38
<< ndcontact >>
rect 3 25 7 29
rect 13 19 17 23
<< pdcontact >>
rect 4 65 8 69
rect 4 58 8 62
rect 14 50 18 54
rect 14 43 18 47
rect 24 56 28 60
rect 24 49 28 53
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
<< psubstratepdiff >>
rect 0 2 32 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 32 2
rect 0 -3 32 -2
<< nsubstratendiff >>
rect 0 82 32 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 32 82
rect 0 77 32 78
<< labels >>
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 44 12 44 6 z
rlabel metal1 16 6 16 6 6 vss
rlabel polycontact 20 36 20 36 6 a
rlabel metal1 20 44 20 44 6 z
rlabel metal1 16 74 16 74 6 vdd
rlabel metal1 28 28 28 28 6 a
<< end >>
