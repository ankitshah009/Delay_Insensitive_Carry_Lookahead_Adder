magic
tech scmos
timestamp 1179385680
<< checkpaint >>
rect -22 -25 222 105
<< ab >>
rect 0 0 200 80
<< pwell >>
rect -4 -7 204 36
<< nwell >>
rect -4 36 204 87
<< polysilicon >>
rect 21 70 23 74
rect 31 70 33 74
rect 41 70 43 74
rect 51 70 53 74
rect 61 70 63 74
rect 71 70 73 74
rect 81 70 83 74
rect 91 70 93 74
rect 101 70 103 74
rect 108 70 110 74
rect 121 70 123 74
rect 128 70 130 74
rect 138 70 140 74
rect 145 70 147 74
rect 157 70 159 74
rect 167 70 169 74
rect 177 70 179 74
rect 10 50 12 55
rect 10 39 12 42
rect 21 39 23 42
rect 31 39 33 42
rect 10 38 33 39
rect 10 34 11 38
rect 15 34 18 38
rect 22 37 33 38
rect 22 34 23 37
rect 10 33 23 34
rect 21 30 23 33
rect 31 30 33 37
rect 41 39 43 42
rect 51 39 53 42
rect 41 38 54 39
rect 41 34 42 38
rect 46 34 49 38
rect 53 35 54 38
rect 61 35 63 42
rect 53 34 63 35
rect 41 33 63 34
rect 41 30 43 33
rect 51 30 53 33
rect 61 30 63 33
rect 71 39 73 42
rect 81 39 83 42
rect 91 39 93 42
rect 101 39 103 42
rect 71 38 93 39
rect 71 34 72 38
rect 76 37 93 38
rect 76 34 83 37
rect 71 33 83 34
rect 71 30 73 33
rect 81 30 83 33
rect 91 30 93 37
rect 97 38 103 39
rect 97 34 98 38
rect 102 34 103 38
rect 97 33 103 34
rect 101 30 103 33
rect 108 39 110 42
rect 121 39 123 42
rect 108 38 123 39
rect 108 34 114 38
rect 118 34 123 38
rect 108 33 123 34
rect 108 30 110 33
rect 121 30 123 33
rect 128 39 130 42
rect 138 39 140 42
rect 128 38 140 39
rect 128 34 129 38
rect 133 34 140 38
rect 128 33 140 34
rect 128 30 130 33
rect 138 30 140 33
rect 145 39 147 42
rect 157 39 159 42
rect 167 39 169 42
rect 177 39 179 42
rect 145 38 179 39
rect 145 34 146 38
rect 150 37 179 38
rect 150 34 160 37
rect 145 33 160 34
rect 145 30 147 33
rect 158 30 160 33
rect 168 30 170 37
rect 21 9 23 14
rect 31 9 33 14
rect 41 11 43 16
rect 51 11 53 16
rect 61 8 63 16
rect 71 12 73 16
rect 81 12 83 16
rect 91 12 93 16
rect 101 8 103 16
rect 108 11 110 16
rect 61 6 103 8
rect 121 11 123 16
rect 128 11 130 16
rect 138 11 140 16
rect 145 11 147 16
rect 158 6 160 10
rect 168 6 170 10
<< ndiffusion >>
rect 14 28 21 30
rect 14 24 15 28
rect 19 24 21 28
rect 14 21 21 24
rect 14 17 15 21
rect 19 17 21 21
rect 14 14 21 17
rect 23 29 31 30
rect 23 25 25 29
rect 29 25 31 29
rect 23 22 31 25
rect 23 18 25 22
rect 29 18 31 22
rect 23 14 31 18
rect 33 28 41 30
rect 33 24 35 28
rect 39 24 41 28
rect 33 21 41 24
rect 33 17 35 21
rect 39 17 41 21
rect 33 16 41 17
rect 43 29 51 30
rect 43 25 45 29
rect 49 25 51 29
rect 43 22 51 25
rect 43 18 45 22
rect 49 18 51 22
rect 43 16 51 18
rect 53 21 61 30
rect 53 17 55 21
rect 59 17 61 21
rect 53 16 61 17
rect 63 29 71 30
rect 63 25 65 29
rect 69 25 71 29
rect 63 22 71 25
rect 63 18 65 22
rect 69 18 71 22
rect 63 16 71 18
rect 73 29 81 30
rect 73 25 75 29
rect 79 25 81 29
rect 73 16 81 25
rect 83 22 91 30
rect 83 18 85 22
rect 89 18 91 22
rect 83 16 91 18
rect 93 29 101 30
rect 93 25 95 29
rect 99 25 101 29
rect 93 16 101 25
rect 103 16 108 30
rect 110 16 121 30
rect 123 16 128 30
rect 130 29 138 30
rect 130 25 132 29
rect 136 25 138 29
rect 130 16 138 25
rect 140 16 145 30
rect 147 16 158 30
rect 33 14 39 16
rect 112 12 119 16
rect 112 8 113 12
rect 117 8 119 12
rect 149 15 158 16
rect 149 11 150 15
rect 154 11 158 15
rect 149 10 158 11
rect 160 29 168 30
rect 160 25 162 29
rect 166 25 168 29
rect 160 22 168 25
rect 160 18 162 22
rect 166 18 168 22
rect 160 10 168 18
rect 170 23 178 30
rect 170 19 172 23
rect 176 19 178 23
rect 170 15 178 19
rect 170 11 172 15
rect 176 11 178 15
rect 170 10 178 11
rect 112 7 119 8
<< pdiffusion >>
rect 14 69 21 70
rect 14 65 15 69
rect 19 65 21 69
rect 14 62 21 65
rect 14 58 15 62
rect 19 58 21 62
rect 14 55 21 58
rect 14 51 15 55
rect 19 51 21 55
rect 14 50 21 51
rect 5 48 10 50
rect 3 47 10 48
rect 3 43 4 47
rect 8 43 10 47
rect 3 42 10 43
rect 12 42 21 50
rect 23 54 31 70
rect 23 50 25 54
rect 29 50 31 54
rect 23 47 31 50
rect 23 43 25 47
rect 29 43 31 47
rect 23 42 31 43
rect 33 69 41 70
rect 33 65 35 69
rect 39 65 41 69
rect 33 62 41 65
rect 33 58 35 62
rect 39 58 41 62
rect 33 55 41 58
rect 33 51 35 55
rect 39 51 41 55
rect 33 42 41 51
rect 43 62 51 70
rect 43 58 45 62
rect 49 58 51 62
rect 43 55 51 58
rect 43 51 45 55
rect 49 51 51 55
rect 43 42 51 51
rect 53 69 61 70
rect 53 65 55 69
rect 59 65 61 69
rect 53 62 61 65
rect 53 58 55 62
rect 59 58 61 62
rect 53 42 61 58
rect 63 62 71 70
rect 63 58 65 62
rect 69 58 71 62
rect 63 55 71 58
rect 63 51 65 55
rect 69 51 71 55
rect 63 42 71 51
rect 73 54 81 70
rect 73 50 75 54
rect 79 50 81 54
rect 73 47 81 50
rect 73 43 75 47
rect 79 43 81 47
rect 73 42 81 43
rect 83 62 91 70
rect 83 58 85 62
rect 89 58 91 62
rect 83 55 91 58
rect 83 51 85 55
rect 89 51 91 55
rect 83 42 91 51
rect 93 54 101 70
rect 93 50 95 54
rect 99 50 101 54
rect 93 47 101 50
rect 93 43 95 47
rect 99 43 101 47
rect 93 42 101 43
rect 103 42 108 70
rect 110 69 121 70
rect 110 65 113 69
rect 117 65 121 69
rect 110 42 121 65
rect 123 42 128 70
rect 130 54 138 70
rect 130 50 132 54
rect 136 50 138 54
rect 130 42 138 50
rect 140 42 145 70
rect 147 69 157 70
rect 147 65 150 69
rect 154 65 157 69
rect 147 42 157 65
rect 159 62 167 70
rect 159 58 161 62
rect 165 58 167 62
rect 159 55 167 58
rect 159 51 161 55
rect 165 51 167 55
rect 159 42 167 51
rect 169 69 177 70
rect 169 65 171 69
rect 175 65 177 69
rect 169 62 177 65
rect 169 58 171 62
rect 175 58 177 62
rect 169 42 177 58
rect 179 55 184 70
rect 179 54 186 55
rect 179 50 181 54
rect 185 50 186 54
rect 179 47 186 50
rect 179 43 181 47
rect 185 43 186 47
rect 179 42 186 43
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect 118 78 122 82
rect 126 78 130 82
rect 134 78 138 82
rect 142 78 146 82
rect 150 78 154 82
rect 158 78 162 82
rect 166 78 170 82
rect 174 78 178 82
rect 182 78 186 82
rect 190 78 194 82
rect 198 78 202 82
rect -2 69 202 78
rect -2 68 15 69
rect 4 59 8 68
rect 19 68 35 69
rect 15 62 19 65
rect 15 55 19 58
rect 39 68 55 69
rect 35 62 39 65
rect 59 68 113 69
rect 112 65 113 68
rect 117 68 150 69
rect 117 65 118 68
rect 149 65 150 68
rect 154 68 171 69
rect 154 65 155 68
rect 170 65 171 68
rect 175 68 202 69
rect 175 65 176 68
rect 35 55 39 58
rect 15 50 19 51
rect 25 54 29 55
rect 35 50 39 51
rect 45 62 49 63
rect 45 55 49 58
rect 55 62 59 65
rect 170 62 176 65
rect 55 57 59 58
rect 64 58 65 62
rect 69 58 85 62
rect 89 58 161 62
rect 165 58 166 62
rect 170 58 171 62
rect 175 58 176 62
rect 189 59 193 68
rect 64 55 69 58
rect 85 55 89 58
rect 64 54 65 55
rect 49 51 65 54
rect 45 50 69 51
rect 74 54 79 55
rect 74 50 75 54
rect 161 55 166 58
rect 85 50 89 51
rect 94 50 95 54
rect 99 50 132 54
rect 136 50 158 54
rect 165 54 166 55
rect 165 51 181 54
rect 161 50 181 51
rect 185 50 186 54
rect 25 47 29 50
rect 74 47 79 50
rect 94 47 99 50
rect 3 43 4 47
rect 8 43 25 47
rect 2 38 22 39
rect 2 34 11 38
rect 15 34 18 38
rect 2 33 22 34
rect 25 38 29 43
rect 66 39 70 47
rect 74 43 75 47
rect 79 43 95 47
rect 82 42 99 43
rect 113 42 150 46
rect 66 38 78 39
rect 25 34 42 38
rect 46 34 49 38
rect 53 34 54 38
rect 66 34 72 38
rect 76 34 78 38
rect 2 25 6 33
rect 25 29 29 34
rect 66 33 78 34
rect 45 29 69 30
rect 82 29 86 42
rect 113 38 119 42
rect 146 38 150 42
rect 97 34 98 38
rect 102 34 108 38
rect 113 34 114 38
rect 118 34 119 38
rect 123 34 129 38
rect 133 34 134 38
rect 104 30 108 34
rect 123 30 127 34
rect 146 33 150 34
rect 15 28 19 29
rect 15 21 19 24
rect 4 12 8 21
rect 25 22 29 25
rect 25 17 29 18
rect 35 28 39 29
rect 35 21 39 24
rect 49 26 65 29
rect 45 22 49 25
rect 64 25 65 26
rect 74 25 75 29
rect 79 25 95 29
rect 99 25 100 29
rect 104 26 127 30
rect 154 29 158 50
rect 180 47 186 50
rect 180 43 181 47
rect 185 43 186 47
rect 131 25 132 29
rect 136 25 158 29
rect 162 29 167 30
rect 166 25 167 29
rect 64 22 69 25
rect 162 22 167 25
rect 45 17 49 18
rect 55 21 59 22
rect 64 18 65 22
rect 69 18 85 22
rect 89 18 162 22
rect 166 18 167 22
rect 172 23 176 24
rect 15 12 19 17
rect 35 12 39 17
rect 55 12 59 17
rect 172 15 176 19
rect 149 12 150 15
rect -2 8 113 12
rect 117 11 150 12
rect 154 12 155 15
rect 154 11 172 12
rect 186 12 190 21
rect 176 11 202 12
rect 117 8 202 11
rect -2 2 202 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 122 2
rect 126 -2 130 2
rect 134 -2 138 2
rect 142 -2 146 2
rect 150 -2 154 2
rect 158 -2 162 2
rect 166 -2 170 2
rect 174 -2 178 2
rect 182 -2 186 2
rect 190 -2 194 2
rect 198 -2 202 2
<< ntransistor >>
rect 21 14 23 30
rect 31 14 33 30
rect 41 16 43 30
rect 51 16 53 30
rect 61 16 63 30
rect 71 16 73 30
rect 81 16 83 30
rect 91 16 93 30
rect 101 16 103 30
rect 108 16 110 30
rect 121 16 123 30
rect 128 16 130 30
rect 138 16 140 30
rect 145 16 147 30
rect 158 10 160 30
rect 168 10 170 30
<< ptransistor >>
rect 10 42 12 50
rect 21 42 23 70
rect 31 42 33 70
rect 41 42 43 70
rect 51 42 53 70
rect 61 42 63 70
rect 71 42 73 70
rect 81 42 83 70
rect 91 42 93 70
rect 101 42 103 70
rect 108 42 110 70
rect 121 42 123 70
rect 128 42 130 70
rect 138 42 140 70
rect 145 42 147 70
rect 157 42 159 70
rect 167 42 169 70
rect 177 42 179 70
<< polycontact >>
rect 11 34 15 38
rect 18 34 22 38
rect 42 34 46 38
rect 49 34 53 38
rect 72 34 76 38
rect 98 34 102 38
rect 114 34 118 38
rect 129 34 133 38
rect 146 34 150 38
<< ndcontact >>
rect 15 24 19 28
rect 15 17 19 21
rect 25 25 29 29
rect 25 18 29 22
rect 35 24 39 28
rect 35 17 39 21
rect 45 25 49 29
rect 45 18 49 22
rect 55 17 59 21
rect 65 25 69 29
rect 65 18 69 22
rect 75 25 79 29
rect 85 18 89 22
rect 95 25 99 29
rect 132 25 136 29
rect 113 8 117 12
rect 150 11 154 15
rect 162 25 166 29
rect 162 18 166 22
rect 172 19 176 23
rect 172 11 176 15
<< pdcontact >>
rect 15 65 19 69
rect 15 58 19 62
rect 15 51 19 55
rect 4 43 8 47
rect 25 50 29 54
rect 25 43 29 47
rect 35 65 39 69
rect 35 58 39 62
rect 35 51 39 55
rect 45 58 49 62
rect 45 51 49 55
rect 55 65 59 69
rect 55 58 59 62
rect 65 58 69 62
rect 65 51 69 55
rect 75 50 79 54
rect 75 43 79 47
rect 85 58 89 62
rect 85 51 89 55
rect 95 50 99 54
rect 95 43 99 47
rect 113 65 117 69
rect 132 50 136 54
rect 150 65 154 69
rect 161 58 165 62
rect 161 51 165 55
rect 171 65 175 69
rect 171 58 175 62
rect 181 50 185 54
rect 181 43 185 47
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
rect 90 -2 94 2
rect 98 -2 102 2
rect 106 -2 110 2
rect 114 -2 118 2
rect 122 -2 126 2
rect 130 -2 134 2
rect 138 -2 142 2
rect 146 -2 150 2
rect 154 -2 158 2
rect 162 -2 166 2
rect 170 -2 174 2
rect 178 -2 182 2
rect 186 -2 190 2
rect 194 -2 198 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
rect 90 78 94 82
rect 98 78 102 82
rect 106 78 110 82
rect 114 78 118 82
rect 122 78 126 82
rect 130 78 134 82
rect 138 78 142 82
rect 146 78 150 82
rect 154 78 158 82
rect 162 78 166 82
rect 170 78 174 82
rect 178 78 182 82
rect 186 78 190 82
rect 194 78 198 82
<< psubstratepdiff >>
rect 0 2 200 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 122 2
rect 126 -2 130 2
rect 134 -2 138 2
rect 142 -2 146 2
rect 150 -2 154 2
rect 158 -2 162 2
rect 166 -2 170 2
rect 174 -2 178 2
rect 182 -2 186 2
rect 190 -2 194 2
rect 198 -2 200 2
rect 0 -3 200 -2
<< nsubstratendiff >>
rect 0 82 200 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect 118 78 122 82
rect 126 78 130 82
rect 134 78 138 82
rect 142 78 146 82
rect 150 78 154 82
rect 158 78 162 82
rect 166 78 170 82
rect 174 78 178 82
rect 182 78 186 82
rect 190 78 194 82
rect 198 78 200 82
rect 0 77 200 78
<< labels >>
rlabel polysilicon 47 36 47 36 6 bn
rlabel polycontact 100 36 100 36 6 bn
rlabel polysilicon 134 36 134 36 6 bn
rlabel polycontact 20 36 20 36 6 b
rlabel polycontact 12 36 12 36 6 b
rlabel metal1 4 32 4 32 6 b
rlabel metal1 16 45 16 45 6 bn
rlabel metal1 47 23 47 23 6 n3
rlabel metal1 39 36 39 36 6 bn
rlabel metal1 47 56 47 56 6 n1
rlabel metal1 66 24 66 24 6 n3
rlabel metal1 84 36 84 36 6 z
rlabel metal1 76 36 76 36 6 c
rlabel metal1 92 44 92 44 6 z
rlabel metal1 68 40 68 40 6 c
rlabel pdcontact 76 52 76 52 6 z
rlabel metal1 87 56 87 56 6 n1
rlabel metal1 66 56 66 56 6 n1
rlabel metal1 100 6 100 6 6 vss
rlabel metal1 102 36 102 36 6 bn
rlabel metal1 128 36 128 36 6 bn
rlabel metal1 116 40 116 40 6 a
rlabel metal1 124 44 124 44 6 a
rlabel metal1 132 44 132 44 6 a
rlabel metal1 100 52 100 52 6 z
rlabel metal1 124 52 124 52 6 z
rlabel metal1 132 52 132 52 6 z
rlabel metal1 116 52 116 52 6 z
rlabel metal1 108 52 108 52 6 z
rlabel metal1 100 74 100 74 6 vdd
rlabel metal1 115 20 115 20 6 n3
rlabel metal1 164 24 164 24 6 n3
rlabel polycontact 148 36 148 36 6 a
rlabel metal1 156 36 156 36 6 z
rlabel metal1 140 44 140 44 6 a
rlabel metal1 140 52 140 52 6 z
rlabel metal1 148 52 148 52 6 z
rlabel metal1 163 56 163 56 6 n1
rlabel metal1 173 52 173 52 6 n1
rlabel metal1 183 48 183 48 6 n1
<< end >>
