magic
tech scmos
timestamp 1182250983
<< checkpaint >>
rect -25 -26 89 114
<< ab >>
rect 0 0 64 88
<< pwell >>
rect -7 -8 71 40
<< nwell >>
rect -7 40 71 96
<< polysilicon >>
rect 5 85 14 86
rect 5 81 6 85
rect 10 81 14 85
rect 5 80 14 81
rect 18 80 27 86
rect 37 80 46 86
rect 50 80 59 86
rect 9 77 11 80
rect 21 77 23 80
rect 41 77 43 80
rect 53 77 55 80
rect 9 48 11 51
rect 21 48 23 51
rect 41 48 43 51
rect 53 48 55 51
rect 2 42 11 48
rect 15 47 30 48
rect 15 43 22 47
rect 26 43 30 47
rect 15 42 30 43
rect 34 47 43 48
rect 34 43 38 47
rect 42 43 43 47
rect 34 42 43 43
rect 47 47 62 48
rect 47 43 54 47
rect 58 43 62 47
rect 47 42 62 43
rect 2 32 17 38
rect 21 37 30 38
rect 21 33 22 37
rect 26 33 30 37
rect 21 32 30 33
rect 34 37 49 38
rect 34 33 38 37
rect 42 33 49 37
rect 34 32 49 33
rect 53 37 62 38
rect 53 33 54 37
rect 58 33 62 37
rect 53 32 62 33
rect 9 29 11 32
rect 21 29 23 32
rect 41 29 43 32
rect 53 29 55 32
rect 9 8 11 11
rect 21 8 23 11
rect 41 8 43 11
rect 53 8 55 11
rect 5 7 14 8
rect 5 3 6 7
rect 10 3 14 7
rect 5 2 14 3
rect 18 2 27 8
rect 37 2 46 8
rect 50 2 59 8
<< ndiffusion >>
rect 2 11 9 29
rect 11 24 21 29
rect 11 20 14 24
rect 18 20 21 24
rect 11 17 21 20
rect 11 13 14 17
rect 18 13 21 17
rect 11 11 21 13
rect 23 25 30 29
rect 23 21 25 25
rect 29 21 30 25
rect 23 17 30 21
rect 23 13 25 17
rect 29 13 30 17
rect 23 11 30 13
rect 34 25 41 29
rect 34 21 35 25
rect 39 21 41 25
rect 34 17 41 21
rect 34 13 35 17
rect 39 13 41 17
rect 34 11 41 13
rect 43 26 53 29
rect 43 22 46 26
rect 50 22 53 26
rect 43 18 53 22
rect 43 14 46 18
rect 50 14 53 18
rect 43 11 53 14
rect 55 24 62 29
rect 55 20 57 24
rect 61 20 62 24
rect 55 17 62 20
rect 55 13 57 17
rect 61 13 62 17
rect 55 11 62 13
<< pdiffusion >>
rect 2 51 9 77
rect 11 75 21 77
rect 11 71 14 75
rect 18 71 21 75
rect 11 68 21 71
rect 11 64 14 68
rect 18 64 21 68
rect 11 51 21 64
rect 23 74 30 77
rect 23 70 25 74
rect 29 70 30 74
rect 23 67 30 70
rect 23 63 25 67
rect 29 63 30 67
rect 23 51 30 63
rect 34 75 41 77
rect 34 71 35 75
rect 39 71 41 75
rect 34 51 41 71
rect 43 74 53 77
rect 43 70 46 74
rect 50 70 53 74
rect 43 67 53 70
rect 43 63 46 67
rect 50 63 53 67
rect 43 51 53 63
rect 55 67 62 77
rect 55 63 57 67
rect 61 63 62 67
rect 55 60 62 63
rect 55 56 57 60
rect 61 56 62 60
rect 55 51 62 56
<< metal1 >>
rect -2 86 2 90
rect 30 86 34 90
rect 2 82 6 85
rect -2 81 6 82
rect 10 81 14 85
rect 18 82 30 85
rect 62 86 66 90
rect 34 82 39 85
rect 18 81 39 82
rect 62 81 66 82
rect 14 75 18 81
rect 35 75 39 81
rect 14 68 18 71
rect 14 63 18 64
rect 25 74 29 75
rect 35 70 39 71
rect 46 74 50 75
rect 25 67 29 70
rect 46 67 50 70
rect 29 63 46 66
rect 25 62 50 63
rect 54 67 61 68
rect 54 63 57 67
rect 54 60 61 63
rect 54 59 57 60
rect 22 47 26 59
rect 46 56 57 59
rect 46 55 61 56
rect 22 37 26 43
rect 22 32 26 33
rect 38 47 42 51
rect 38 37 42 43
rect 38 29 42 33
rect 46 26 50 55
rect 54 47 58 51
rect 54 37 58 43
rect 54 29 58 33
rect 14 24 18 25
rect 24 21 25 25
rect 29 21 35 25
rect 39 21 40 25
rect 14 17 18 20
rect 46 18 50 22
rect 24 13 25 17
rect 29 13 35 17
rect 39 13 40 17
rect 46 13 50 14
rect 57 24 61 25
rect 57 17 61 20
rect 14 7 18 13
rect 57 7 61 13
rect -2 6 6 7
rect 2 3 6 6
rect 10 3 14 7
rect 18 6 34 7
rect 18 3 30 6
rect -2 -2 2 2
rect 57 6 66 7
rect 57 3 62 6
rect 30 -2 34 2
rect 62 -2 66 2
<< metal2 >>
rect -2 86 66 90
rect 2 85 30 86
rect 2 82 14 85
rect -2 81 14 82
rect 18 82 30 85
rect 34 82 62 86
rect 18 81 66 82
rect -2 80 66 81
rect -2 7 66 8
rect -2 6 14 7
rect 2 3 14 6
rect 18 6 66 7
rect 18 3 30 6
rect 2 2 30 3
rect 34 2 62 6
rect -2 -2 66 2
<< ntransistor >>
rect 9 11 11 29
rect 21 11 23 29
rect 41 11 43 29
rect 53 11 55 29
<< ptransistor >>
rect 9 51 11 77
rect 21 51 23 77
rect 41 51 43 77
rect 53 51 55 77
<< polycontact >>
rect 6 81 10 85
rect 22 43 26 47
rect 38 43 42 47
rect 54 43 58 47
rect 22 33 26 37
rect 38 33 42 37
rect 54 33 58 37
rect 6 3 10 7
<< ndcontact >>
rect 14 20 18 24
rect 14 13 18 17
rect 25 21 29 25
rect 25 13 29 17
rect 35 21 39 25
rect 35 13 39 17
rect 46 22 50 26
rect 46 14 50 18
rect 57 20 61 24
rect 57 13 61 17
<< pdcontact >>
rect 14 71 18 75
rect 14 64 18 68
rect 25 70 29 74
rect 25 63 29 67
rect 35 71 39 75
rect 46 70 50 74
rect 46 63 50 67
rect 57 63 61 67
rect 57 56 61 60
<< m2contact >>
rect -2 82 2 86
rect 14 81 18 85
rect 30 82 34 86
rect 62 82 66 86
rect -2 2 2 6
rect 14 3 18 7
rect 30 2 34 6
rect 62 2 66 6
<< psubstratepcontact >>
rect -2 2 2 6
rect 30 2 34 6
rect 62 2 66 6
<< nsubstratencontact >>
rect -2 82 2 86
rect 30 82 34 86
rect 62 82 66 86
<< psubstratepdiff >>
rect -3 6 3 7
rect -3 2 -2 6
rect 2 2 3 6
rect 29 6 35 7
rect 29 2 30 6
rect 34 2 35 6
rect 61 6 67 7
rect 61 2 62 6
rect 66 2 67 6
rect -3 0 3 2
rect 29 0 35 2
rect 61 0 67 2
<< nsubstratendiff >>
rect -3 86 3 88
rect 29 86 35 88
rect 61 86 67 88
rect -3 82 -2 86
rect 2 82 3 86
rect -3 81 3 82
rect 29 82 30 86
rect 34 82 35 86
rect 29 81 35 82
rect 61 82 62 86
rect 66 82 67 86
rect 61 81 67 82
<< labels >>
rlabel metal1 24 48 24 48 6 a1
rlabel metal1 40 40 40 40 6 a2
rlabel metal1 48 36 48 36 6 z
rlabel metal1 56 40 56 40 6 b
rlabel metal1 56 64 56 64 6 z
rlabel m2contact 32 4 32 4 6 vss
rlabel m2contact 32 84 32 84 6 vdd
<< end >>
