magic
tech scmos
timestamp 1179385952
<< checkpaint >>
rect -22 -22 54 94
<< ab >>
rect 0 0 32 72
<< pwell >>
rect -4 -4 36 32
<< nwell >>
rect -4 32 36 76
<< polysilicon >>
rect 10 66 12 70
rect 20 57 22 61
rect 10 35 12 38
rect 20 35 22 38
rect 9 34 22 35
rect 9 30 17 34
rect 21 30 22 34
rect 9 29 22 30
rect 9 26 11 29
rect 9 9 11 14
<< ndiffusion >>
rect 2 25 9 26
rect 2 21 3 25
rect 7 21 9 25
rect 2 20 9 21
rect 4 14 9 20
rect 11 19 19 26
rect 11 15 13 19
rect 17 15 19 19
rect 11 14 19 15
<< pdiffusion >>
rect 2 65 10 66
rect 2 61 4 65
rect 8 61 10 65
rect 2 58 10 61
rect 2 54 4 58
rect 8 54 10 58
rect 2 38 10 54
rect 12 57 17 66
rect 12 50 20 57
rect 12 46 14 50
rect 18 46 20 50
rect 12 43 20 46
rect 12 39 14 43
rect 18 39 20 43
rect 12 38 20 39
rect 22 56 30 57
rect 22 52 24 56
rect 28 52 30 56
rect 22 49 30 52
rect 22 45 24 49
rect 28 45 30 49
rect 22 38 30 45
<< metal1 >>
rect -2 68 34 72
rect -2 65 23 68
rect -2 64 4 65
rect 3 61 4 64
rect 8 64 23 65
rect 27 64 34 68
rect 8 61 9 64
rect 3 58 9 61
rect 3 54 4 58
rect 8 54 9 58
rect 23 56 29 64
rect 23 52 24 56
rect 28 52 29 56
rect 14 50 18 51
rect 14 43 18 46
rect 23 49 29 52
rect 23 45 24 49
rect 28 45 29 49
rect 2 39 14 43
rect 18 39 23 42
rect 2 38 23 39
rect 2 26 6 38
rect 16 30 17 34
rect 21 30 30 34
rect 2 25 7 26
rect 2 21 3 25
rect 26 21 30 30
rect 2 20 7 21
rect 13 19 17 20
rect 13 8 17 15
rect -2 4 24 8
rect 28 4 34 8
rect -2 0 34 4
<< ntransistor >>
rect 9 14 11 26
<< ptransistor >>
rect 10 38 12 66
rect 20 38 22 57
<< polycontact >>
rect 17 30 21 34
<< ndcontact >>
rect 3 21 7 25
rect 13 15 17 19
<< pdcontact >>
rect 4 61 8 65
rect 4 54 8 58
rect 14 46 18 50
rect 14 39 18 43
rect 24 52 28 56
rect 24 45 28 49
<< psubstratepcontact >>
rect 24 4 28 8
<< nsubstratencontact >>
rect 23 64 27 68
<< psubstratepdiff >>
rect 23 8 29 24
rect 23 4 24 8
rect 28 4 29 8
rect 23 3 29 4
<< nsubstratendiff >>
rect 21 68 29 69
rect 21 64 23 68
rect 27 64 29 68
rect 21 63 29 64
<< labels >>
rlabel metal1 4 32 4 32 6 z
rlabel metal1 12 40 12 40 6 z
rlabel metal1 16 4 16 4 6 vss
rlabel polycontact 20 32 20 32 6 a
rlabel metal1 20 40 20 40 6 z
rlabel metal1 16 68 16 68 6 vdd
rlabel metal1 28 24 28 24 6 a
<< end >>
