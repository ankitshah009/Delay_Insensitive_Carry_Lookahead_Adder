magic
tech scmos
timestamp 1182081799
<< checkpaint >>
rect -25 -26 89 114
<< ab >>
rect 0 0 64 88
<< pwell >>
rect -7 -8 71 40
<< nwell >>
rect -7 40 71 96
<< polysilicon >>
rect 5 85 14 86
rect 5 81 6 85
rect 10 81 14 85
rect 5 80 14 81
rect 18 80 27 86
rect 37 80 46 86
rect 50 80 59 86
rect 9 77 11 80
rect 21 77 23 80
rect 41 77 43 80
rect 53 77 55 80
rect 9 48 11 51
rect 21 48 23 51
rect 41 48 43 51
rect 53 48 55 51
rect 2 42 11 48
rect 15 47 30 48
rect 15 43 22 47
rect 26 43 30 47
rect 15 42 30 43
rect 34 47 43 48
rect 34 43 38 47
rect 42 43 43 47
rect 34 42 43 43
rect 47 47 62 48
rect 47 43 54 47
rect 58 43 62 47
rect 47 42 62 43
rect 2 32 17 38
rect 21 37 30 38
rect 21 33 22 37
rect 26 33 30 37
rect 21 32 30 33
rect 34 37 49 38
rect 34 33 38 37
rect 42 33 49 37
rect 34 32 49 33
rect 53 37 62 38
rect 53 33 54 37
rect 58 33 62 37
rect 53 32 62 33
rect 9 29 11 32
rect 21 29 23 32
rect 41 29 43 32
rect 53 29 55 32
rect 9 8 11 11
rect 21 8 23 11
rect 41 8 43 11
rect 53 8 55 11
rect 5 7 14 8
rect 5 3 6 7
rect 10 3 14 7
rect 5 2 14 3
rect 18 2 27 8
rect 37 2 46 8
rect 50 2 59 8
<< ndiffusion >>
rect 2 11 9 29
rect 11 24 21 29
rect 11 20 14 24
rect 18 20 21 24
rect 11 17 21 20
rect 11 13 14 17
rect 18 13 21 17
rect 11 11 21 13
rect 23 25 30 29
rect 23 21 25 25
rect 29 21 30 25
rect 23 18 30 21
rect 23 14 25 18
rect 29 14 30 18
rect 23 11 30 14
rect 34 17 41 29
rect 34 13 35 17
rect 39 13 41 17
rect 34 11 41 13
rect 43 11 53 29
rect 55 25 62 29
rect 55 21 57 25
rect 61 21 62 25
rect 55 18 62 21
rect 55 14 57 18
rect 61 14 62 18
rect 55 11 62 14
<< pdiffusion >>
rect 2 51 9 77
rect 11 75 21 77
rect 11 71 14 75
rect 18 71 21 75
rect 11 68 21 71
rect 11 64 14 68
rect 18 64 21 68
rect 11 51 21 64
rect 23 66 30 77
rect 23 62 25 66
rect 29 62 30 66
rect 23 59 30 62
rect 23 55 25 59
rect 29 55 30 59
rect 23 51 30 55
rect 34 75 41 77
rect 34 71 35 75
rect 39 71 41 75
rect 34 68 41 71
rect 34 64 35 68
rect 39 64 41 68
rect 34 51 41 64
rect 43 66 53 77
rect 43 62 46 66
rect 50 62 53 66
rect 43 58 53 62
rect 43 54 46 58
rect 50 54 53 58
rect 43 51 53 54
rect 55 75 62 77
rect 55 71 57 75
rect 61 71 62 75
rect 55 68 62 71
rect 55 64 57 68
rect 61 64 62 68
rect 55 51 62 64
<< metal1 >>
rect -2 86 2 90
rect 30 86 34 90
rect 2 82 6 85
rect -2 81 6 82
rect 10 82 30 85
rect 62 86 66 90
rect 34 82 62 85
rect 10 81 66 82
rect 14 75 18 81
rect 14 68 18 71
rect 35 75 39 81
rect 35 68 39 71
rect 14 63 18 64
rect 22 66 29 67
rect 22 62 25 66
rect 57 75 61 81
rect 57 68 61 71
rect 35 63 39 64
rect 46 66 50 67
rect 22 59 29 62
rect 14 48 18 59
rect 22 55 25 59
rect 57 63 61 64
rect 46 58 50 62
rect 29 55 46 58
rect 22 54 46 55
rect 14 47 26 48
rect 14 44 22 47
rect 22 37 26 43
rect 22 32 26 33
rect 38 47 42 48
rect 38 37 42 43
rect 25 25 29 26
rect 14 24 18 25
rect 14 17 18 20
rect 38 21 42 33
rect 46 26 50 54
rect 54 47 58 59
rect 54 37 58 43
rect 54 32 58 33
rect 46 25 61 26
rect 46 22 57 25
rect 54 21 57 22
rect 25 18 29 21
rect 54 18 61 21
rect 29 14 35 17
rect 25 13 35 14
rect 39 13 40 17
rect 54 14 57 18
rect 54 13 61 14
rect 14 7 18 13
rect -2 6 6 7
rect 2 3 6 6
rect 10 6 34 7
rect 10 3 30 6
rect -2 -2 2 2
rect 30 -2 34 2
rect 62 6 66 7
rect 62 -2 66 2
<< metal2 >>
rect -2 86 66 90
rect 2 82 30 86
rect 34 82 62 86
rect -2 80 66 82
rect -2 6 66 8
rect 2 2 30 6
rect 34 2 62 6
rect -2 -2 66 2
<< ntransistor >>
rect 9 11 11 29
rect 21 11 23 29
rect 41 11 43 29
rect 53 11 55 29
<< ptransistor >>
rect 9 51 11 77
rect 21 51 23 77
rect 41 51 43 77
rect 53 51 55 77
<< polycontact >>
rect 6 81 10 85
rect 22 43 26 47
rect 38 43 42 47
rect 54 43 58 47
rect 22 33 26 37
rect 38 33 42 37
rect 54 33 58 37
rect 6 3 10 7
<< ndcontact >>
rect 14 20 18 24
rect 14 13 18 17
rect 25 21 29 25
rect 25 14 29 18
rect 35 13 39 17
rect 57 21 61 25
rect 57 14 61 18
<< pdcontact >>
rect 14 71 18 75
rect 14 64 18 68
rect 25 62 29 66
rect 25 55 29 59
rect 35 71 39 75
rect 35 64 39 68
rect 46 62 50 66
rect 46 54 50 58
rect 57 71 61 75
rect 57 64 61 68
<< m2contact >>
rect -2 82 2 86
rect 30 82 34 86
rect 62 82 66 86
rect -2 2 2 6
rect 30 2 34 6
rect 62 2 66 6
<< psubstratepcontact >>
rect -2 2 2 6
rect 30 2 34 6
rect 62 2 66 6
<< nsubstratencontact >>
rect -2 82 2 86
rect 30 82 34 86
rect 62 82 66 86
<< psubstratepdiff >>
rect -3 6 3 7
rect -3 2 -2 6
rect 2 2 3 6
rect 29 6 35 7
rect 29 2 30 6
rect 34 2 35 6
rect 61 6 67 7
rect 61 2 62 6
rect 66 2 67 6
rect -3 0 3 2
rect 29 0 35 2
rect 61 0 67 2
<< nsubstratendiff >>
rect -3 86 3 88
rect 29 86 35 88
rect 61 86 67 88
rect -3 82 -2 86
rect 2 82 3 86
rect -3 81 3 82
rect 29 82 30 86
rect 34 82 35 86
rect 29 81 35 82
rect 61 82 62 86
rect 66 82 67 86
rect 61 81 67 82
<< labels >>
rlabel metal1 16 52 16 52 6 a
rlabel metal1 24 40 24 40 6 a
rlabel metal1 32 56 32 56 6 z
rlabel metal1 24 64 24 64 6 z
rlabel metal1 40 32 40 32 6 b
rlabel metal1 48 48 48 48 6 z
rlabel metal1 40 56 40 56 6 z
rlabel metal1 56 20 56 20 6 z
rlabel metal1 56 48 56 48 6 c
rlabel m2contact 32 4 32 4 6 vss
rlabel m2contact 32 84 32 84 6 vdd
<< end >>
