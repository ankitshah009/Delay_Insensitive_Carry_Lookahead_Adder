.subckt nao2o22_x1 i0 i1 i2 i3 nq vdd vss
*   SPICE3 file   created from nao2o22_x1.ext -      technology: scmos
m00 w1     i0     vdd    vdd p w=39u  l=2.3636u ad=195p     pd=49u      as=294p     ps=94u
m01 nq     i1     w1     vdd p w=39u  l=2.3636u ad=195p     pd=49u      as=195p     ps=49u
m02 w2     i3     nq     vdd p w=39u  l=2.3636u ad=195p     pd=49u      as=195p     ps=49u
m03 vdd    i2     w2     vdd p w=39u  l=2.3636u ad=294p     pd=94u      as=195p     ps=49u
m04 nq     i0     w3     vss n w=19u  l=2.3636u ad=119p     pd=37u      as=123.5p   ps=41.5u
m05 w3     i1     nq     vss n w=19u  l=2.3636u ad=123.5p   pd=41.5u    as=119p     ps=37u
m06 vss    i3     w3     vss n w=19u  l=2.3636u ad=95p      pd=29u      as=123.5p   ps=41.5u
m07 w3     i2     vss    vss n w=19u  l=2.3636u ad=123.5p   pd=41.5u    as=95p      ps=29u
C0  nq     i2     0.106f
C1  w2     i3     0.057f
C2  vss    i0     0.010f
C3  w1     vdd    0.019f
C4  w3     i1     0.013f
C5  vdd    i2     0.143f
C6  nq     i1     0.262f
C7  vdd    i1     0.049f
C8  i2     i3     0.361f
C9  w3     nq     0.109f
C10 i3     i1     0.150f
C11 i2     i0     0.057f
C12 vss    i2     0.013f
C13 i1     i0     0.310f
C14 w3     i3     0.029f
C15 nq     vdd    0.069f
C16 vss    i1     0.010f
C17 w3     i0     0.013f
C18 nq     i3     0.283f
C19 vss    w3     0.342f
C20 nq     i0     0.087f
C21 vdd    i3     0.068f
C22 w1     i1     0.057f
C23 vss    nq     0.052f
C24 i2     i1     0.082f
C25 vdd    i0     0.064f
C26 vss    vdd    0.003f
C27 i3     i0     0.082f
C28 w3     i2     0.029f
C29 vss    i3     0.013f
C30 w2     vdd    0.019f
C32 nq     vss    0.016f
C34 i2     vss    0.029f
C35 i3     vss    0.034f
C36 i1     vss    0.029f
C37 i0     vss    0.025f
.ends
