magic
tech scmos
timestamp 1185094634
<< checkpaint >>
rect -22 -22 72 122
<< ab >>
rect 0 0 50 100
<< pwell >>
rect -4 -4 54 48
<< nwell >>
rect -4 48 54 104
<< polysilicon >>
rect 13 83 15 88
rect 25 83 27 88
rect 37 83 39 88
rect 13 53 15 63
rect 25 60 27 63
rect 25 59 33 60
rect 25 55 28 59
rect 32 55 33 59
rect 25 54 33 55
rect 13 52 21 53
rect 13 48 16 52
rect 20 48 21 52
rect 13 47 21 48
rect 13 33 15 47
rect 25 36 27 54
rect 37 53 39 63
rect 37 52 43 53
rect 37 48 38 52
rect 42 48 43 52
rect 37 47 43 48
rect 37 41 39 47
rect 33 39 39 41
rect 33 36 35 39
rect 13 22 15 27
rect 25 22 27 27
rect 33 22 35 27
<< ndiffusion >>
rect 20 33 25 36
rect 5 32 13 33
rect 5 28 6 32
rect 10 28 13 32
rect 5 27 13 28
rect 15 32 25 33
rect 15 28 18 32
rect 22 28 25 32
rect 15 27 25 28
rect 27 27 33 36
rect 35 32 43 36
rect 35 28 38 32
rect 42 28 43 32
rect 35 27 43 28
<< pdiffusion >>
rect 29 92 35 93
rect 29 88 30 92
rect 34 88 35 92
rect 29 83 35 88
rect 5 82 13 83
rect 5 78 6 82
rect 10 78 13 82
rect 5 74 13 78
rect 5 70 6 74
rect 10 70 13 74
rect 5 69 13 70
rect 8 63 13 69
rect 15 82 25 83
rect 15 78 18 82
rect 22 78 25 82
rect 15 63 25 78
rect 27 63 37 83
rect 39 82 47 83
rect 39 78 42 82
rect 46 78 47 82
rect 39 77 47 78
rect 39 63 44 77
<< metal1 >>
rect -2 96 52 100
rect -2 92 8 96
rect 12 92 18 96
rect 22 92 52 96
rect -2 88 30 92
rect 34 88 52 92
rect 6 82 12 83
rect 10 78 12 82
rect 17 78 18 82
rect 22 78 42 82
rect 46 78 47 82
rect 6 74 12 78
rect 10 70 12 74
rect 6 69 12 70
rect 8 43 12 69
rect 18 68 33 73
rect 18 53 22 68
rect 38 63 42 73
rect 16 52 22 53
rect 20 48 22 52
rect 16 47 22 48
rect 28 59 42 63
rect 32 57 42 59
rect 28 47 32 55
rect 38 52 42 53
rect 38 43 42 48
rect 8 37 22 43
rect 6 32 10 33
rect 6 12 10 28
rect 18 32 22 37
rect 18 27 22 28
rect 28 37 42 43
rect 28 27 32 37
rect 38 32 42 33
rect 38 12 42 28
rect -2 8 52 12
rect -2 4 8 8
rect 12 4 18 8
rect 22 4 52 8
rect -2 0 52 4
<< ntransistor >>
rect 13 27 15 33
rect 25 27 27 36
rect 33 27 35 36
<< ptransistor >>
rect 13 63 15 83
rect 25 63 27 83
rect 37 63 39 83
<< polycontact >>
rect 28 55 32 59
rect 16 48 20 52
rect 38 48 42 52
<< ndcontact >>
rect 6 28 10 32
rect 18 28 22 32
rect 38 28 42 32
<< pdcontact >>
rect 30 88 34 92
rect 6 78 10 82
rect 6 70 10 74
rect 18 78 22 82
rect 42 78 46 82
<< psubstratepcontact >>
rect 8 4 12 8
rect 18 4 22 8
<< nsubstratencontact >>
rect 8 92 12 96
rect 18 92 22 96
<< psubstratepdiff >>
rect 7 8 23 9
rect 7 4 8 8
rect 12 4 18 8
rect 22 4 23 8
rect 7 3 23 4
<< nsubstratendiff >>
rect 7 96 23 97
rect 7 92 8 96
rect 12 92 18 96
rect 22 92 23 96
rect 7 91 23 92
<< labels >>
rlabel metal1 20 35 20 35 6 z
rlabel metal1 10 60 10 60 6 z
rlabel metal1 20 60 20 60 6 b
rlabel metal1 25 6 25 6 6 vss
rlabel metal1 30 35 30 35 6 a1
rlabel metal1 30 70 30 70 6 b
rlabel metal1 30 55 30 55 6 a2
rlabel metal1 25 94 25 94 6 vdd
rlabel metal1 40 45 40 45 6 a1
rlabel metal1 40 65 40 65 6 a2
rlabel metal1 32 80 32 80 6 n2
<< end >>
