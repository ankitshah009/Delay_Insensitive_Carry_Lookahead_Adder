magic
tech scmos
timestamp 1179385259
<< checkpaint >>
rect -22 -22 62 94
<< ab >>
rect 0 0 40 72
<< pwell >>
rect -4 -4 44 32
<< nwell >>
rect -4 32 44 76
<< polysilicon >>
rect 29 62 31 67
rect 9 54 11 59
rect 19 54 21 59
rect 29 43 31 46
rect 29 42 35 43
rect 29 38 30 42
rect 34 38 35 42
rect 9 35 11 38
rect 9 34 15 35
rect 9 30 10 34
rect 14 30 15 34
rect 9 29 15 30
rect 19 31 21 38
rect 29 37 35 38
rect 19 30 25 31
rect 12 21 14 29
rect 19 26 20 30
rect 24 26 25 30
rect 19 25 25 26
rect 22 22 24 25
rect 29 22 31 37
rect 12 11 14 15
rect 22 11 24 15
rect 29 11 31 15
<< ndiffusion >>
rect 17 21 22 22
rect 3 15 12 21
rect 14 20 22 21
rect 14 16 16 20
rect 20 16 22 20
rect 14 15 22 16
rect 24 15 29 22
rect 31 15 38 22
rect 3 8 10 15
rect 33 9 38 15
rect 3 4 5 8
rect 9 4 10 8
rect 3 3 10 4
rect 32 8 38 9
rect 32 4 33 8
rect 37 4 38 8
rect 32 3 38 4
<< pdiffusion >>
rect 21 68 27 69
rect 21 64 22 68
rect 26 64 27 68
rect 21 62 27 64
rect 21 61 29 62
rect 23 54 29 61
rect 4 51 9 54
rect 2 50 9 51
rect 2 46 3 50
rect 7 46 9 50
rect 2 43 9 46
rect 2 39 3 43
rect 7 39 9 43
rect 2 38 9 39
rect 11 53 19 54
rect 11 49 13 53
rect 17 49 19 53
rect 11 38 19 49
rect 21 46 29 54
rect 31 59 36 62
rect 31 58 38 59
rect 31 54 33 58
rect 37 54 38 58
rect 31 51 38 54
rect 31 47 33 51
rect 37 47 38 51
rect 31 46 38 47
rect 21 38 27 46
<< metal1 >>
rect -2 68 42 72
rect -2 64 4 68
rect 8 64 12 68
rect 16 64 22 68
rect 26 64 42 68
rect 13 58 37 59
rect 13 55 33 58
rect 13 53 17 55
rect 2 50 7 51
rect 2 46 3 50
rect 33 51 37 54
rect 13 48 17 49
rect 2 43 7 46
rect 26 43 30 51
rect 33 46 37 47
rect 2 39 3 43
rect 2 38 7 39
rect 2 19 6 38
rect 10 37 22 43
rect 26 42 38 43
rect 26 38 30 42
rect 34 38 38 42
rect 26 37 38 38
rect 10 34 14 37
rect 10 29 14 30
rect 19 26 20 30
rect 24 29 25 30
rect 24 26 30 29
rect 19 25 30 26
rect 16 20 20 21
rect 2 16 16 19
rect 26 19 30 25
rect 20 16 22 19
rect 2 13 22 16
rect 26 13 38 19
rect -2 4 5 8
rect 9 4 15 8
rect 19 4 23 8
rect 27 4 33 8
rect 37 4 42 8
rect -2 0 42 4
<< ntransistor >>
rect 12 15 14 21
rect 22 15 24 22
rect 29 15 31 22
<< ptransistor >>
rect 9 38 11 54
rect 19 38 21 54
rect 29 46 31 62
<< polycontact >>
rect 30 38 34 42
rect 10 30 14 34
rect 20 26 24 30
<< ndcontact >>
rect 16 16 20 20
rect 5 4 9 8
rect 33 4 37 8
<< pdcontact >>
rect 22 64 26 68
rect 3 46 7 50
rect 3 39 7 43
rect 13 49 17 53
rect 33 54 37 58
rect 33 47 37 51
<< psubstratepcontact >>
rect 15 4 19 8
rect 23 4 27 8
<< nsubstratencontact >>
rect 4 64 8 68
rect 12 64 16 68
<< psubstratepdiff >>
rect 14 8 28 9
rect 14 4 15 8
rect 19 4 23 8
rect 27 4 28 8
rect 14 3 28 4
<< nsubstratendiff >>
rect 3 68 17 69
rect 3 64 4 68
rect 8 64 12 68
rect 16 64 17 68
rect 3 63 17 64
<< labels >>
rlabel metal1 4 32 4 32 6 z
rlabel metal1 12 16 12 16 6 z
rlabel metal1 12 36 12 36 6 b
rlabel metal1 15 53 15 53 6 n1
rlabel metal1 20 4 20 4 6 vss
rlabel metal1 28 20 28 20 6 a2
rlabel metal1 20 16 20 16 6 z
rlabel metal1 20 40 20 40 6 b
rlabel metal1 28 44 28 44 6 a1
rlabel metal1 20 68 20 68 6 vdd
rlabel metal1 36 16 36 16 6 a2
rlabel metal1 36 40 36 40 6 a1
rlabel metal1 35 52 35 52 6 n1
<< end >>
