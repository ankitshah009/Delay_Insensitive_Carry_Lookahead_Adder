magic
tech scmos
timestamp 1180600617
<< checkpaint >>
rect -22 -22 102 122
<< ab >>
rect 0 0 80 100
<< pwell >>
rect -4 -4 84 48
<< nwell >>
rect -4 48 84 104
<< polysilicon >>
rect 55 94 57 98
rect 67 94 69 98
rect 11 85 13 89
rect 23 86 25 90
rect 33 85 35 89
rect 45 85 47 89
rect 11 53 13 65
rect 23 63 25 66
rect 33 63 35 66
rect 45 63 47 66
rect 19 61 25 63
rect 31 61 35 63
rect 41 61 47 63
rect 19 53 21 61
rect 31 53 33 61
rect 7 52 13 53
rect 7 48 8 52
rect 12 48 13 52
rect 7 47 13 48
rect 17 52 23 53
rect 17 48 18 52
rect 22 48 23 52
rect 17 47 23 48
rect 27 52 33 53
rect 27 48 28 52
rect 32 48 33 52
rect 27 47 33 48
rect 11 34 13 47
rect 19 34 21 47
rect 27 34 29 47
rect 41 43 43 61
rect 55 53 57 56
rect 67 53 69 56
rect 47 52 69 53
rect 47 48 48 52
rect 52 48 69 52
rect 47 47 69 48
rect 37 42 43 43
rect 37 39 38 42
rect 35 38 38 39
rect 42 38 43 42
rect 35 37 43 38
rect 35 34 37 37
rect 55 25 57 47
rect 67 25 69 47
rect 11 11 13 15
rect 19 11 21 15
rect 27 11 29 15
rect 35 11 37 15
rect 55 2 57 6
rect 67 2 69 6
<< ndiffusion >>
rect 3 15 11 34
rect 13 15 19 34
rect 21 15 27 34
rect 29 15 35 34
rect 37 23 43 34
rect 37 22 45 23
rect 37 18 40 22
rect 44 18 45 22
rect 37 17 45 18
rect 37 15 42 17
rect 3 12 9 15
rect 3 8 4 12
rect 8 8 9 12
rect 50 11 55 25
rect 47 10 55 11
rect 3 7 9 8
rect 47 6 48 10
rect 52 6 55 10
rect 57 22 67 25
rect 57 18 60 22
rect 64 18 67 22
rect 57 6 67 18
rect 69 22 77 25
rect 69 18 72 22
rect 76 18 77 22
rect 69 12 77 18
rect 69 8 72 12
rect 76 8 77 12
rect 69 6 77 8
rect 47 5 53 6
<< pdiffusion >>
rect 27 96 33 97
rect 3 92 9 93
rect 3 88 4 92
rect 8 88 9 92
rect 27 92 28 96
rect 32 92 33 96
rect 27 91 33 92
rect 47 96 53 97
rect 47 92 48 96
rect 52 94 53 96
rect 52 92 55 94
rect 47 91 55 92
rect 3 85 9 88
rect 27 86 31 91
rect 15 85 23 86
rect 3 82 11 85
rect 3 78 4 82
rect 8 78 11 82
rect 3 65 11 78
rect 13 82 23 85
rect 13 78 16 82
rect 20 78 23 82
rect 13 66 23 78
rect 25 85 31 86
rect 49 85 55 91
rect 25 66 33 85
rect 35 82 45 85
rect 35 78 38 82
rect 42 78 45 82
rect 35 66 45 78
rect 47 66 55 85
rect 13 65 18 66
rect 49 56 55 66
rect 57 82 67 94
rect 57 78 60 82
rect 64 78 67 82
rect 57 72 67 78
rect 57 68 60 72
rect 64 68 67 72
rect 57 62 67 68
rect 57 58 60 62
rect 64 58 67 62
rect 57 56 67 58
rect 69 92 77 94
rect 69 88 72 92
rect 76 88 77 92
rect 69 82 77 88
rect 69 78 72 82
rect 76 78 77 82
rect 69 72 77 78
rect 69 68 72 72
rect 76 68 77 72
rect 69 62 77 68
rect 69 58 72 62
rect 76 58 77 62
rect 69 56 77 58
<< metal1 >>
rect -2 96 82 100
rect -2 92 28 96
rect 32 92 48 96
rect 52 92 82 96
rect -2 88 4 92
rect 8 88 72 92
rect 76 88 82 92
rect 4 82 8 88
rect 58 82 62 83
rect 72 82 76 88
rect 15 78 16 82
rect 20 78 38 82
rect 42 78 53 82
rect 4 77 8 78
rect 8 52 12 73
rect 8 17 12 48
rect 18 52 22 73
rect 18 17 22 48
rect 28 52 32 73
rect 28 17 32 48
rect 38 42 42 73
rect 49 52 53 78
rect 47 48 48 52
rect 52 48 53 52
rect 38 27 42 38
rect 49 22 53 48
rect 39 18 40 22
rect 44 18 53 22
rect 58 78 60 82
rect 64 78 65 82
rect 58 72 62 78
rect 72 72 76 78
rect 58 68 60 72
rect 64 68 65 72
rect 58 62 62 68
rect 72 62 76 68
rect 58 58 60 62
rect 64 58 65 62
rect 58 22 62 58
rect 72 57 76 58
rect 72 22 76 23
rect 58 18 60 22
rect 64 18 65 22
rect 58 17 62 18
rect 72 12 76 18
rect -2 8 4 12
rect 8 10 72 12
rect 8 8 48 10
rect -2 4 18 8
rect 22 4 34 8
rect 38 6 48 8
rect 52 8 72 10
rect 76 8 82 12
rect 52 6 82 8
rect 38 4 82 6
rect -2 0 82 4
<< ntransistor >>
rect 11 15 13 34
rect 19 15 21 34
rect 27 15 29 34
rect 35 15 37 34
rect 55 6 57 25
rect 67 6 69 25
<< ptransistor >>
rect 11 65 13 85
rect 23 66 25 86
rect 33 66 35 85
rect 45 66 47 85
rect 55 56 57 94
rect 67 56 69 94
<< polycontact >>
rect 8 48 12 52
rect 18 48 22 52
rect 28 48 32 52
rect 48 48 52 52
rect 38 38 42 42
<< ndcontact >>
rect 40 18 44 22
rect 4 8 8 12
rect 48 6 52 10
rect 60 18 64 22
rect 72 18 76 22
rect 72 8 76 12
<< pdcontact >>
rect 4 88 8 92
rect 28 92 32 96
rect 48 92 52 96
rect 4 78 8 82
rect 16 78 20 82
rect 38 78 42 82
rect 60 78 64 82
rect 60 68 64 72
rect 60 58 64 62
rect 72 88 76 92
rect 72 78 76 82
rect 72 68 76 72
rect 72 58 76 62
<< psubstratepcontact >>
rect 18 4 22 8
rect 34 4 38 8
<< psubstratepdiff >>
rect 17 8 39 9
rect 17 4 18 8
rect 22 4 34 8
rect 38 4 39 8
rect 17 3 39 4
<< labels >>
rlabel metal1 10 45 10 45 6 i0
rlabel metal1 20 45 20 45 6 i1
rlabel metal1 30 45 30 45 6 i2
rlabel metal1 40 6 40 6 6 vss
rlabel metal1 40 50 40 50 6 i3
rlabel metal1 40 94 40 94 6 vdd
rlabel metal1 60 50 60 50 6 q
<< end >>
