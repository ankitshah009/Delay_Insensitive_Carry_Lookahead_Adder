magic
tech scmos
timestamp 1179386294
<< checkpaint >>
rect -22 -22 54 94
<< ab >>
rect 0 0 32 72
<< pwell >>
rect -4 -4 36 32
<< nwell >>
rect -4 32 36 76
<< polysilicon >>
rect 10 57 12 62
rect 20 57 22 61
rect 10 35 12 43
rect 9 34 15 35
rect 9 30 10 34
rect 14 30 15 34
rect 9 29 15 30
rect 9 19 11 29
rect 20 28 22 43
rect 20 27 26 28
rect 20 24 21 27
rect 16 23 21 24
rect 25 23 26 27
rect 16 22 26 23
rect 16 19 18 22
rect 9 2 11 7
rect 16 2 18 7
<< ndiffusion >>
rect 2 18 9 19
rect 2 14 3 18
rect 7 14 9 18
rect 2 13 9 14
rect 4 7 9 13
rect 11 7 16 19
rect 18 12 30 19
rect 18 8 25 12
rect 29 8 30 12
rect 18 7 30 8
<< pdiffusion >>
rect 2 58 8 59
rect 2 54 3 58
rect 7 57 8 58
rect 7 54 10 57
rect 2 43 10 54
rect 12 56 20 57
rect 12 52 14 56
rect 18 52 20 56
rect 12 49 20 52
rect 12 45 14 49
rect 18 45 20 49
rect 12 43 20 45
rect 22 56 30 57
rect 22 52 25 56
rect 29 52 30 56
rect 22 49 30 52
rect 22 45 25 49
rect 29 45 30 49
rect 22 43 30 45
<< metal1 >>
rect -2 68 34 72
rect -2 64 16 68
rect 20 64 24 68
rect 28 64 34 68
rect 2 58 8 64
rect 2 54 3 58
rect 7 54 8 58
rect 24 56 30 64
rect 13 52 14 56
rect 18 52 19 56
rect 13 50 19 52
rect 2 49 19 50
rect 2 45 14 49
rect 18 45 19 49
rect 24 52 25 56
rect 29 52 30 56
rect 24 49 30 52
rect 24 45 25 49
rect 29 45 30 49
rect 2 19 6 45
rect 17 38 23 42
rect 10 34 23 38
rect 10 29 14 30
rect 18 23 21 27
rect 25 23 30 27
rect 18 21 30 23
rect 2 18 7 19
rect 2 14 3 18
rect 2 13 7 14
rect 18 13 22 21
rect 25 12 29 13
rect -2 0 34 8
<< ntransistor >>
rect 9 7 11 19
rect 16 7 18 19
<< ptransistor >>
rect 10 43 12 57
rect 20 43 22 57
<< polycontact >>
rect 10 30 14 34
rect 21 23 25 27
<< ndcontact >>
rect 3 14 7 18
rect 25 8 29 12
<< pdcontact >>
rect 3 54 7 58
rect 14 52 18 56
rect 14 45 18 49
rect 25 52 29 56
rect 25 45 29 49
<< nsubstratencontact >>
rect 16 64 20 68
rect 24 64 28 68
<< nsubstratendiff >>
rect 15 68 29 69
rect 15 64 16 68
rect 20 64 24 68
rect 28 64 29 68
rect 15 63 29 64
<< labels >>
rlabel metal1 4 28 4 28 6 z
rlabel polycontact 12 32 12 32 6 b
rlabel metal1 12 48 12 48 6 z
rlabel metal1 16 4 16 4 6 vss
rlabel metal1 20 20 20 20 6 a
rlabel metal1 20 40 20 40 6 b
rlabel metal1 16 68 16 68 6 vdd
rlabel metal1 28 24 28 24 6 a
<< end >>
