.subckt xor2v0x1 a b vdd vss z
*   SPICE3 file   created from xor2v0x1.ext -      technology: scmos
m00 vdd    b      bn     vdd p w=27u  l=2.3636u ad=216p     pd=49.2u    as=147p     ps=68u
m01 an     a      vdd    vdd p w=18u  l=2.3636u ad=72p      pd=26u      as=144p     ps=32.8u
m02 z      bn     an     vdd p w=18u  l=2.3636u ad=75.6p    pd=28u      as=72p      ps=26u
m03 bn     an     z      vdd p w=27u  l=2.3636u ad=147p     pd=68u      as=113.4p   ps=42u
m04 vss    b      bn     vss n w=9u   l=2.3636u ad=77.4p    pd=32.4u    as=57p      ps=32u
m05 an     a      vss    vss n w=9u   l=2.3636u ad=36p      pd=17u      as=77.4p    ps=32.4u
m06 z      b      an     vss n w=9u   l=2.3636u ad=37.2857p pd=17.1429u as=36p      ps=17u
m07 w1     bn     z      vss n w=12u  l=2.3636u ad=30p      pd=17u      as=49.7143p ps=22.8571u
m08 vss    an     w1     vss n w=12u  l=2.3636u ad=103.2p   pd=43.2u    as=30p      ps=17u
C0  vss    bn     0.063f
C1  z      a      0.011f
C2  a      bn     0.199f
C3  z      an     0.376f
C4  vss    b      0.018f
C5  a      b      0.091f
C6  bn     an     0.440f
C7  z      vdd    0.042f
C8  an     b      0.024f
C9  bn     vdd    0.330f
C10 w1     z      0.010f
C11 b      vdd    0.103f
C12 vss    a      0.076f
C13 z      bn     0.226f
C14 vss    an     0.087f
C15 a      an     0.049f
C16 z      b      0.003f
C17 bn     b      0.136f
C18 a      vdd    0.013f
C19 an     vdd    0.046f
C20 vss    z      0.154f
C22 z      vss    0.012f
C23 a      vss    0.030f
C24 bn     vss    0.035f
C25 an     vss    0.029f
C26 b      vss    0.054f
.ends
