magic
tech scmos
timestamp 1179386405
<< checkpaint >>
rect -22 -22 78 94
<< ab >>
rect 0 0 56 72
<< pwell >>
rect -4 -4 60 32
<< nwell >>
rect -4 32 60 76
<< polysilicon >>
rect 14 65 16 70
rect 24 65 26 70
rect 35 57 37 62
rect 45 57 47 61
rect 14 35 16 38
rect 24 35 26 38
rect 35 35 37 38
rect 45 35 47 38
rect 9 34 26 35
rect 9 30 10 34
rect 14 30 26 34
rect 9 29 26 30
rect 24 26 26 29
rect 31 34 47 35
rect 31 30 42 34
rect 46 30 47 34
rect 31 29 47 30
rect 31 26 33 29
rect 24 2 26 7
rect 31 2 33 7
<< ndiffusion >>
rect 17 25 24 26
rect 17 21 18 25
rect 22 21 24 25
rect 17 18 24 21
rect 17 14 18 18
rect 22 14 24 18
rect 17 13 24 14
rect 19 7 24 13
rect 26 7 31 26
rect 33 19 41 26
rect 33 15 35 19
rect 39 15 41 19
rect 33 12 41 15
rect 33 8 35 12
rect 39 8 41 12
rect 33 7 41 8
<< pdiffusion >>
rect 6 64 14 65
rect 6 60 8 64
rect 12 60 14 64
rect 6 57 14 60
rect 6 53 8 57
rect 12 53 14 57
rect 6 38 14 53
rect 16 50 24 65
rect 16 46 18 50
rect 22 46 24 50
rect 16 43 24 46
rect 16 39 18 43
rect 22 39 24 43
rect 16 38 24 39
rect 26 64 33 65
rect 26 60 28 64
rect 32 60 33 64
rect 26 57 33 60
rect 26 53 28 57
rect 32 53 35 57
rect 26 38 35 53
rect 37 50 45 57
rect 37 46 39 50
rect 43 46 45 50
rect 37 43 45 46
rect 37 39 39 43
rect 43 39 45 43
rect 37 38 45 39
rect 47 56 54 57
rect 47 52 49 56
rect 53 52 54 56
rect 47 49 54 52
rect 47 45 49 49
rect 53 45 54 49
rect 47 38 54 45
<< metal1 >>
rect -2 68 58 72
rect -2 64 40 68
rect 44 64 48 68
rect 52 64 58 68
rect 8 57 12 60
rect 8 52 12 53
rect 28 57 32 60
rect 28 52 32 53
rect 49 56 53 64
rect 18 50 22 51
rect 18 43 22 46
rect 2 35 6 43
rect 39 50 43 51
rect 39 43 43 46
rect 49 49 53 52
rect 49 44 53 45
rect 22 39 39 42
rect 18 38 43 39
rect 2 34 14 35
rect 2 30 10 34
rect 2 29 14 30
rect 18 25 22 38
rect 41 30 42 34
rect 46 30 54 34
rect 50 21 54 30
rect 18 18 22 21
rect 18 13 22 14
rect 35 19 39 20
rect 35 12 39 15
rect -2 4 4 8
rect 8 4 48 8
rect 52 4 58 8
rect -2 0 58 4
<< ntransistor >>
rect 24 7 26 26
rect 31 7 33 26
<< ptransistor >>
rect 14 38 16 65
rect 24 38 26 65
rect 35 38 37 57
rect 45 38 47 57
<< polycontact >>
rect 10 30 14 34
rect 42 30 46 34
<< ndcontact >>
rect 18 21 22 25
rect 18 14 22 18
rect 35 15 39 19
rect 35 8 39 12
<< pdcontact >>
rect 8 60 12 64
rect 8 53 12 57
rect 18 46 22 50
rect 18 39 22 43
rect 28 60 32 64
rect 28 53 32 57
rect 39 46 43 50
rect 39 39 43 43
rect 49 52 53 56
rect 49 45 53 49
<< psubstratepcontact >>
rect 4 4 8 8
rect 48 4 52 8
<< nsubstratencontact >>
rect 40 64 44 68
rect 48 64 52 68
<< psubstratepdiff >>
rect 3 8 9 24
rect 3 4 4 8
rect 8 4 9 8
rect 47 8 53 24
rect 3 3 9 4
rect 47 4 48 8
rect 52 4 53 8
rect 47 3 53 4
<< nsubstratendiff >>
rect 39 68 53 69
rect 39 64 40 68
rect 44 64 48 68
rect 52 64 53 68
rect 39 63 53 64
<< labels >>
rlabel metal1 4 36 4 36 6 b
rlabel polycontact 12 32 12 32 6 b
rlabel metal1 20 32 20 32 6 z
rlabel metal1 28 4 28 4 6 vss
rlabel metal1 36 40 36 40 6 z
rlabel metal1 28 40 28 40 6 z
rlabel metal1 28 68 28 68 6 vdd
rlabel polycontact 44 32 44 32 6 a
rlabel metal1 52 24 52 24 6 a
<< end >>
