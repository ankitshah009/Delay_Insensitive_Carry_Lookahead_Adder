magic
tech scmos
timestamp 1179385539
<< checkpaint >>
rect -22 -25 62 105
<< ab >>
rect 0 0 40 80
<< pwell >>
rect -4 -7 44 36
<< nwell >>
rect -4 36 44 87
<< polysilicon >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 9 38 11 42
rect 19 38 21 42
rect 29 39 31 42
rect 26 38 32 39
rect 9 37 22 38
rect 9 33 17 37
rect 21 33 22 37
rect 26 34 27 38
rect 31 34 32 38
rect 26 33 32 34
rect 9 32 22 33
rect 9 29 11 32
rect 19 29 21 32
rect 29 29 31 33
rect 9 10 11 15
rect 19 10 21 15
rect 29 10 31 15
<< ndiffusion >>
rect 2 28 9 29
rect 2 24 3 28
rect 7 24 9 28
rect 2 20 9 24
rect 2 16 3 20
rect 7 16 9 20
rect 2 15 9 16
rect 11 22 19 29
rect 11 18 13 22
rect 17 18 19 22
rect 11 15 19 18
rect 21 20 29 29
rect 21 16 23 20
rect 27 16 29 20
rect 21 15 29 16
rect 31 28 38 29
rect 31 24 33 28
rect 37 24 38 28
rect 31 21 38 24
rect 31 17 33 21
rect 37 17 38 21
rect 31 15 38 17
<< pdiffusion >>
rect 2 69 9 70
rect 2 65 3 69
rect 7 65 9 69
rect 2 62 9 65
rect 2 58 3 62
rect 7 58 9 62
rect 2 42 9 58
rect 11 62 19 70
rect 11 58 13 62
rect 17 58 19 62
rect 11 55 19 58
rect 11 51 13 55
rect 17 51 19 55
rect 11 42 19 51
rect 21 69 29 70
rect 21 65 23 69
rect 27 65 29 69
rect 21 62 29 65
rect 21 58 23 62
rect 27 58 29 62
rect 21 42 29 58
rect 31 62 36 70
rect 31 61 38 62
rect 31 57 33 61
rect 37 57 38 61
rect 31 54 38 57
rect 31 50 33 54
rect 37 50 38 54
rect 31 49 38 50
rect 31 42 36 49
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect -2 69 42 78
rect -2 68 3 69
rect 2 65 3 68
rect 7 68 23 69
rect 7 65 8 68
rect 2 62 8 65
rect 22 65 23 68
rect 27 68 42 69
rect 27 65 28 68
rect 2 58 3 62
rect 7 58 8 62
rect 13 62 17 63
rect 22 62 28 65
rect 22 58 23 62
rect 27 58 28 62
rect 33 61 38 62
rect 13 55 17 58
rect 2 51 13 54
rect 2 50 17 51
rect 37 57 38 61
rect 33 54 38 57
rect 37 50 38 54
rect 2 37 6 50
rect 33 49 38 50
rect 17 42 31 46
rect 26 38 31 42
rect 17 37 21 38
rect 2 33 14 37
rect 3 28 7 29
rect 3 20 7 24
rect 10 23 14 33
rect 26 34 27 38
rect 26 33 31 34
rect 17 30 21 33
rect 34 30 38 49
rect 17 28 38 30
rect 17 26 33 28
rect 37 26 38 28
rect 10 22 17 23
rect 10 18 13 22
rect 33 21 37 24
rect 10 17 17 18
rect 23 20 27 21
rect 3 12 7 16
rect 33 16 37 17
rect 23 12 27 16
rect -2 2 42 12
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
<< ntransistor >>
rect 9 15 11 29
rect 19 15 21 29
rect 29 15 31 29
<< ptransistor >>
rect 9 42 11 70
rect 19 42 21 70
rect 29 42 31 70
<< polycontact >>
rect 17 33 21 37
rect 27 34 31 38
<< ndcontact >>
rect 3 24 7 28
rect 3 16 7 20
rect 13 18 17 22
rect 23 16 27 20
rect 33 24 37 28
rect 33 17 37 21
<< pdcontact >>
rect 3 65 7 69
rect 3 58 7 62
rect 13 58 17 62
rect 13 51 17 55
rect 23 65 27 69
rect 23 58 27 62
rect 33 57 37 61
rect 33 50 37 54
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
<< psubstratepdiff >>
rect 0 2 40 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 40 2
rect 0 -3 40 -2
<< nsubstratendiff >>
rect 0 82 40 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 40 82
rect 0 77 40 78
<< labels >>
rlabel polysilicon 15 35 15 35 6 an
rlabel metal1 4 40 4 40 6 z
rlabel metal1 12 24 12 24 6 z
rlabel metal1 12 52 12 52 6 z
rlabel metal1 20 6 20 6 6 vss
rlabel metal1 19 32 19 32 6 an
rlabel metal1 28 40 28 40 6 a
rlabel metal1 20 44 20 44 6 a
rlabel metal1 20 74 20 74 6 vdd
rlabel metal1 35 23 35 23 6 an
rlabel metal1 36 44 36 44 6 an
<< end >>
