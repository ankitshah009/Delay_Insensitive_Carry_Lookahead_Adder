.subckt bf1_w05 a vdd vss z
*   SPICE3 file   created from bf1_w05.ext -      technology: scmos
m00 vdd    a      an     vdd p w=9u   l=2.3636u ad=88.5p    pd=46u      as=75p      ps=38u
m01 z      an     vdd    vdd p w=9u   l=2.3636u ad=63p      pd=34u      as=88.5p    ps=46u
m02 z      an     vss    vss n w=6u   l=2.3636u ad=54p      pd=30u      as=72p      ps=40u
m03 vss    a      an     vss n w=6u   l=2.3636u ad=72p      pd=40u      as=54p      ps=30u
C0  vss    an     0.154f
C1  z      a      0.030f
C2  vss    vdd    0.011f
C3  an     vdd    0.136f
C4  vss    z      0.044f
C5  vss    a      0.002f
C6  z      an     0.024f
C7  z      vdd    0.047f
C8  an     a      0.193f
C9  a      vdd    0.079f
C11 z      vss    0.017f
C12 an     vss    0.029f
C13 a      vss    0.036f
.ends
