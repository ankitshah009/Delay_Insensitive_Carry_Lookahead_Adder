magic
tech scmos
timestamp 1179387175
<< checkpaint >>
rect -22 -25 86 105
<< ab >>
rect 0 0 64 80
<< pwell >>
rect -4 -7 68 36
<< nwell >>
rect -4 36 68 87
<< polysilicon >>
rect 9 63 11 68
rect 19 63 21 68
rect 29 63 31 68
rect 36 63 38 68
rect 46 59 48 64
rect 53 59 55 64
rect 9 39 11 43
rect 19 39 21 43
rect 9 38 21 39
rect 9 34 16 38
rect 20 34 21 38
rect 29 34 31 43
rect 36 40 38 43
rect 46 40 48 43
rect 36 38 48 40
rect 53 40 55 43
rect 53 39 62 40
rect 53 38 57 39
rect 38 37 48 38
rect 9 33 21 34
rect 28 33 34 34
rect 9 30 11 33
rect 28 29 29 33
rect 33 29 34 33
rect 28 28 34 29
rect 38 33 41 37
rect 45 33 48 37
rect 56 35 57 38
rect 61 35 62 39
rect 56 34 62 35
rect 38 32 48 33
rect 28 25 30 28
rect 38 25 40 32
rect 28 10 30 15
rect 38 10 40 15
rect 9 6 11 10
<< ndiffusion >>
rect 2 29 9 30
rect 2 25 3 29
rect 7 25 9 29
rect 2 22 9 25
rect 2 18 3 22
rect 7 18 9 22
rect 2 17 9 18
rect 4 10 9 17
rect 11 25 26 30
rect 11 23 28 25
rect 11 19 13 23
rect 17 19 28 23
rect 11 15 28 19
rect 30 24 38 25
rect 30 20 32 24
rect 36 20 38 24
rect 30 15 38 20
rect 40 20 48 25
rect 40 16 42 20
rect 46 16 48 20
rect 40 15 48 16
rect 11 11 13 15
rect 17 11 21 15
rect 25 11 26 15
rect 11 10 26 11
<< pdiffusion >>
rect 2 62 9 63
rect 2 58 3 62
rect 7 58 9 62
rect 2 55 9 58
rect 2 51 3 55
rect 7 51 9 55
rect 2 43 9 51
rect 11 55 19 63
rect 11 51 13 55
rect 17 51 19 55
rect 11 48 19 51
rect 11 44 13 48
rect 17 44 19 48
rect 11 43 19 44
rect 21 62 29 63
rect 21 58 23 62
rect 27 58 29 62
rect 21 43 29 58
rect 31 43 36 63
rect 38 59 43 63
rect 38 54 46 59
rect 38 50 40 54
rect 44 50 46 54
rect 38 43 46 50
rect 48 43 53 59
rect 55 58 62 59
rect 55 54 57 58
rect 61 54 62 58
rect 55 43 62 54
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect -2 68 66 78
rect 2 62 8 68
rect 2 58 3 62
rect 7 58 8 62
rect 22 62 28 68
rect 22 58 23 62
rect 27 58 28 62
rect 57 58 61 68
rect 2 55 8 58
rect 2 51 3 55
rect 7 51 8 55
rect 13 55 17 56
rect 13 48 17 51
rect 2 44 13 47
rect 2 42 17 44
rect 21 50 40 54
rect 44 50 45 54
rect 57 53 61 54
rect 2 30 6 42
rect 21 38 25 50
rect 58 46 62 47
rect 15 34 16 38
rect 20 34 25 38
rect 2 29 7 30
rect 2 25 3 29
rect 2 22 7 25
rect 21 24 25 34
rect 29 42 62 46
rect 29 33 33 42
rect 56 39 62 42
rect 29 28 33 29
rect 41 37 47 38
rect 45 33 47 37
rect 56 35 57 39
rect 61 35 62 39
rect 58 33 62 35
rect 41 31 47 33
rect 41 25 54 31
rect 2 18 3 22
rect 2 17 7 18
rect 13 23 17 24
rect 21 20 32 24
rect 36 20 37 24
rect 42 20 46 21
rect 13 15 17 19
rect -2 11 13 12
rect 21 15 25 16
rect 17 11 21 12
rect 42 12 46 16
rect 25 11 66 12
rect -2 2 66 11
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
<< ntransistor >>
rect 9 10 11 30
rect 28 15 30 25
rect 38 15 40 25
<< ptransistor >>
rect 9 43 11 63
rect 19 43 21 63
rect 29 43 31 63
rect 36 43 38 63
rect 46 43 48 59
rect 53 43 55 59
<< polycontact >>
rect 16 34 20 38
rect 29 29 33 33
rect 41 33 45 37
rect 57 35 61 39
<< ndcontact >>
rect 3 25 7 29
rect 3 18 7 22
rect 13 19 17 23
rect 32 20 36 24
rect 42 16 46 20
rect 13 11 17 15
rect 21 11 25 15
<< pdcontact >>
rect 3 58 7 62
rect 3 51 7 55
rect 13 51 17 55
rect 13 44 17 48
rect 23 58 27 62
rect 40 50 44 54
rect 57 54 61 58
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
<< psubstratepdiff >>
rect 0 2 64 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 64 2
rect 0 -3 64 -2
<< nsubstratendiff >>
rect 0 82 64 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 64 82
rect 0 77 64 78
<< labels >>
rlabel polysilicon 15 36 15 36 6 zn
rlabel metal1 4 32 4 32 6 z
rlabel metal1 12 44 12 44 6 z
rlabel metal1 32 6 32 6 6 vss
rlabel metal1 29 22 29 22 6 zn
rlabel metal1 20 36 20 36 6 zn
rlabel metal1 36 44 36 44 6 a
rlabel metal1 32 74 32 74 6 vdd
rlabel metal1 44 32 44 32 6 b
rlabel metal1 44 44 44 44 6 a
rlabel metal1 33 52 33 52 6 zn
rlabel metal1 52 28 52 28 6 b
rlabel metal1 52 44 52 44 6 a
rlabel metal1 60 40 60 40 6 a
<< end >>
