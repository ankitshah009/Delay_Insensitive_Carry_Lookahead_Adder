magic
tech scmos
timestamp 1180639982
<< checkpaint >>
rect -24 -26 64 126
<< ab >>
rect 0 0 40 100
<< pwell >>
rect -4 -6 44 49
<< nwell >>
rect -4 49 44 106
<< polysilicon >>
rect 15 83 17 88
rect 27 83 29 88
rect 15 50 17 63
rect 27 50 29 63
rect 15 49 23 50
rect 15 45 18 49
rect 22 45 23 49
rect 15 44 23 45
rect 27 49 33 50
rect 27 45 28 49
rect 32 45 33 49
rect 27 44 33 45
rect 15 33 17 44
rect 27 33 29 44
rect 15 18 17 23
rect 27 18 29 23
<< ndiffusion >>
rect 7 32 15 33
rect 7 28 8 32
rect 12 28 15 32
rect 7 27 15 28
rect 10 23 15 27
rect 17 23 27 33
rect 29 32 37 33
rect 29 28 32 32
rect 36 28 37 32
rect 29 27 37 28
rect 29 23 34 27
rect 19 22 25 23
rect 19 18 20 22
rect 24 18 25 22
rect 19 17 25 18
<< pdiffusion >>
rect 10 77 15 83
rect 7 76 15 77
rect 7 72 8 76
rect 12 72 15 76
rect 7 68 15 72
rect 7 64 8 68
rect 12 64 15 68
rect 7 63 15 64
rect 17 82 27 83
rect 17 78 20 82
rect 24 78 27 82
rect 17 63 27 78
rect 29 82 37 83
rect 29 78 32 82
rect 36 78 37 82
rect 29 74 37 78
rect 29 70 32 74
rect 36 70 37 74
rect 29 69 37 70
rect 29 63 34 69
<< metal1 >>
rect -2 88 42 100
rect 20 82 24 88
rect 20 77 24 78
rect 32 82 36 83
rect 8 76 12 77
rect 32 74 36 78
rect 8 68 12 72
rect 8 32 12 64
rect 18 70 32 72
rect 18 68 36 70
rect 18 49 22 68
rect 18 32 22 45
rect 28 49 32 63
rect 28 37 32 45
rect 18 28 32 32
rect 36 28 37 32
rect 8 27 12 28
rect 20 22 24 23
rect 20 12 24 18
rect -2 0 42 12
<< ntransistor >>
rect 15 23 17 33
rect 27 23 29 33
<< ptransistor >>
rect 15 63 17 83
rect 27 63 29 83
<< polycontact >>
rect 18 45 22 49
rect 28 45 32 49
<< ndcontact >>
rect 8 28 12 32
rect 32 28 36 32
rect 20 18 24 22
<< pdcontact >>
rect 8 72 12 76
rect 8 64 12 68
rect 20 78 24 82
rect 32 78 36 82
rect 32 70 36 74
<< psubstratepcontact >>
rect 8 4 12 8
rect 18 4 22 8
<< nsubstratencontact >>
rect 8 92 12 96
rect 18 92 22 96
<< psubstratepdiff >>
rect 7 8 23 9
rect 7 4 8 8
rect 12 4 18 8
rect 22 4 23 8
rect 7 3 23 4
<< nsubstratendiff >>
rect 7 96 23 97
rect 7 92 8 96
rect 12 92 18 96
rect 22 92 23 96
rect 7 91 23 92
<< labels >>
rlabel polycontact 19 47 19 47 6 an
rlabel metal1 10 50 10 50 6 z
rlabel metal1 10 50 10 50 6 z
rlabel metal1 20 6 20 6 6 vss
rlabel metal1 20 6 20 6 6 vss
rlabel metal1 20 50 20 50 6 an
rlabel metal1 20 94 20 94 6 vdd
rlabel metal1 20 94 20 94 6 vdd
rlabel metal1 27 30 27 30 6 an
rlabel metal1 30 50 30 50 6 a
rlabel metal1 30 50 30 50 6 a
rlabel metal1 34 75 34 75 6 an
<< end >>
