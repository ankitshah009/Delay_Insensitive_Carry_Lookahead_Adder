magic
tech scmos
timestamp 1179385393
<< checkpaint >>
rect -22 -22 78 94
<< ab >>
rect 0 0 56 72
<< pwell >>
rect -4 -4 60 32
<< nwell >>
rect -4 32 60 76
<< polysilicon >>
rect 9 54 11 59
rect 19 54 21 59
rect 30 55 32 60
rect 40 55 42 60
rect 9 29 11 46
rect 19 43 21 46
rect 19 42 25 43
rect 19 38 20 42
rect 24 38 25 42
rect 19 37 25 38
rect 9 28 15 29
rect 9 24 10 28
rect 14 24 15 28
rect 9 23 15 24
rect 12 20 14 23
rect 19 20 21 37
rect 30 29 32 46
rect 40 43 42 46
rect 39 42 47 43
rect 39 38 42 42
rect 46 38 47 42
rect 39 37 47 38
rect 25 28 34 29
rect 25 24 26 28
rect 30 24 34 28
rect 25 23 34 24
rect 32 20 34 23
rect 39 20 41 37
rect 12 8 14 13
rect 19 8 21 13
rect 32 8 34 13
rect 39 8 41 13
<< ndiffusion >>
rect 5 19 12 20
rect 5 15 6 19
rect 10 15 12 19
rect 5 13 12 15
rect 14 13 19 20
rect 21 18 32 20
rect 21 14 26 18
rect 30 14 32 18
rect 21 13 32 14
rect 34 13 39 20
rect 41 19 48 20
rect 41 15 43 19
rect 47 15 48 19
rect 41 13 48 15
<< pdiffusion >>
rect 23 54 30 55
rect 2 53 9 54
rect 2 49 3 53
rect 7 49 9 53
rect 2 46 9 49
rect 11 51 19 54
rect 11 47 13 51
rect 17 47 19 51
rect 11 46 19 47
rect 21 53 30 54
rect 21 49 24 53
rect 28 49 30 53
rect 21 46 30 49
rect 32 51 40 55
rect 32 47 34 51
rect 38 47 40 51
rect 32 46 40 47
rect 42 53 50 55
rect 42 49 45 53
rect 49 49 50 53
rect 42 46 50 49
<< metal1 >>
rect -2 68 58 72
rect -2 64 4 68
rect 8 64 12 68
rect 16 64 58 68
rect 3 53 7 64
rect 24 53 28 64
rect 3 48 7 49
rect 10 51 17 52
rect 10 47 13 51
rect 45 53 49 64
rect 24 48 28 49
rect 34 51 38 52
rect 10 46 17 47
rect 45 48 49 49
rect 10 43 14 46
rect 2 39 14 43
rect 34 42 38 47
rect 2 15 6 39
rect 19 38 20 42
rect 24 38 38 42
rect 41 42 54 43
rect 41 38 42 42
rect 46 38 54 42
rect 10 28 14 35
rect 26 28 30 35
rect 34 34 38 38
rect 34 30 47 34
rect 14 24 22 27
rect 10 23 22 24
rect 10 15 14 19
rect 2 13 14 15
rect 18 13 22 23
rect 30 24 38 27
rect 26 21 38 24
rect 43 19 47 30
rect 50 21 54 38
rect 25 14 26 18
rect 30 14 31 18
rect 43 14 47 15
rect 25 8 31 14
rect -2 4 48 8
rect 52 4 58 8
rect -2 0 58 4
<< ntransistor >>
rect 12 13 14 20
rect 19 13 21 20
rect 32 13 34 20
rect 39 13 41 20
<< ptransistor >>
rect 9 46 11 54
rect 19 46 21 54
rect 30 46 32 55
rect 40 46 42 55
<< polycontact >>
rect 20 38 24 42
rect 10 24 14 28
rect 42 38 46 42
rect 26 24 30 28
<< ndcontact >>
rect 6 15 10 19
rect 26 14 30 18
rect 43 15 47 19
<< pdcontact >>
rect 3 49 7 53
rect 13 47 17 51
rect 24 49 28 53
rect 34 47 38 51
rect 45 49 49 53
<< psubstratepcontact >>
rect 48 4 52 8
<< nsubstratencontact >>
rect 4 64 8 68
rect 12 64 16 68
<< psubstratepdiff >>
rect 47 8 53 9
rect 47 4 48 8
rect 52 4 53 8
rect 47 3 53 4
<< nsubstratendiff >>
rect 3 68 17 69
rect 3 64 4 68
rect 8 64 12 68
rect 16 64 17 68
rect 3 63 17 64
<< labels >>
rlabel polycontact 22 40 22 40 6 an
rlabel metal1 4 28 4 28 6 z
rlabel metal1 20 20 20 20 6 b
rlabel metal1 12 16 12 16 6 z
rlabel metal1 12 32 12 32 6 b
rlabel metal1 12 48 12 48 6 z
rlabel metal1 28 4 28 4 6 vss
rlabel metal1 28 28 28 28 6 a1
rlabel metal1 36 24 36 24 6 a1
rlabel metal1 28 40 28 40 6 an
rlabel metal1 28 68 28 68 6 vdd
rlabel metal1 45 24 45 24 6 an
rlabel metal1 52 32 52 32 6 a2
rlabel polycontact 44 40 44 40 6 a2
<< end >>
