magic
tech scmos
timestamp 1179385387
<< checkpaint >>
rect -22 -25 166 105
<< ab >>
rect 0 0 144 80
<< pwell >>
rect -4 -7 148 36
<< nwell >>
rect -4 36 148 87
<< polysilicon >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 39 70 41 74
rect 49 70 51 74
rect 59 70 61 74
rect 69 70 71 74
rect 79 70 81 74
rect 89 70 91 74
rect 99 70 101 74
rect 109 70 111 74
rect 119 70 121 74
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 9 38 31 39
rect 9 34 10 38
rect 14 37 31 38
rect 14 34 21 37
rect 9 33 21 34
rect 19 27 21 33
rect 29 27 31 37
rect 39 39 41 42
rect 49 39 51 42
rect 59 39 61 42
rect 39 38 61 39
rect 39 34 44 38
rect 48 34 56 38
rect 60 34 61 38
rect 39 33 61 34
rect 39 30 41 33
rect 49 30 51 33
rect 59 30 61 33
rect 69 39 71 42
rect 79 39 81 42
rect 89 39 91 42
rect 69 38 91 39
rect 69 34 76 38
rect 80 34 84 38
rect 88 34 91 38
rect 69 33 91 34
rect 69 30 71 33
rect 79 30 81 33
rect 89 30 91 33
rect 99 39 101 42
rect 109 39 111 42
rect 119 39 121 42
rect 99 38 121 39
rect 99 37 109 38
rect 99 30 101 37
rect 108 34 109 37
rect 113 34 116 38
rect 120 34 121 38
rect 108 33 121 34
rect 109 30 111 33
rect 119 30 121 33
rect 19 11 21 16
rect 29 11 31 16
rect 39 7 41 12
rect 49 7 51 12
rect 59 7 61 12
rect 69 7 71 12
rect 79 7 81 12
rect 89 7 91 12
rect 99 7 101 12
rect 109 7 111 12
rect 119 7 121 12
<< ndiffusion >>
rect 34 27 39 30
rect 12 26 19 27
rect 12 22 13 26
rect 17 22 19 26
rect 12 21 19 22
rect 14 16 19 21
rect 21 21 29 27
rect 21 17 23 21
rect 27 17 29 21
rect 21 16 29 17
rect 31 26 39 27
rect 31 22 33 26
rect 37 22 39 26
rect 31 16 39 22
rect 34 12 39 16
rect 41 21 49 30
rect 41 17 43 21
rect 47 17 49 21
rect 41 12 49 17
rect 51 29 59 30
rect 51 25 53 29
rect 57 25 59 29
rect 51 12 59 25
rect 61 28 69 30
rect 61 24 63 28
rect 67 24 69 28
rect 61 21 69 24
rect 61 17 63 21
rect 67 17 69 21
rect 61 12 69 17
rect 71 29 79 30
rect 71 25 73 29
rect 77 25 79 29
rect 71 12 79 25
rect 81 21 89 30
rect 81 17 83 21
rect 87 17 89 21
rect 81 12 89 17
rect 91 29 99 30
rect 91 25 93 29
rect 97 25 99 29
rect 91 22 99 25
rect 91 18 93 22
rect 97 18 99 22
rect 91 12 99 18
rect 101 17 109 30
rect 101 13 103 17
rect 107 13 109 17
rect 101 12 109 13
rect 111 28 119 30
rect 111 24 113 28
rect 117 24 119 28
rect 111 21 119 24
rect 111 17 113 21
rect 117 17 119 21
rect 111 12 119 17
rect 121 25 128 30
rect 121 21 123 25
rect 127 21 128 25
rect 121 17 128 21
rect 121 13 123 17
rect 127 13 128 17
rect 121 12 128 13
<< pdiffusion >>
rect 4 55 9 70
rect 2 54 9 55
rect 2 50 3 54
rect 7 50 9 54
rect 2 47 9 50
rect 2 43 3 47
rect 7 43 9 47
rect 2 42 9 43
rect 11 62 19 70
rect 11 58 13 62
rect 17 58 19 62
rect 11 55 19 58
rect 11 51 13 55
rect 17 51 19 55
rect 11 42 19 51
rect 21 54 29 70
rect 21 50 23 54
rect 27 50 29 54
rect 21 47 29 50
rect 21 43 23 47
rect 27 43 29 47
rect 21 42 29 43
rect 31 62 39 70
rect 31 58 33 62
rect 37 58 39 62
rect 31 55 39 58
rect 31 51 33 55
rect 37 51 39 55
rect 31 42 39 51
rect 41 69 49 70
rect 41 65 43 69
rect 47 65 49 69
rect 41 62 49 65
rect 41 58 43 62
rect 47 58 49 62
rect 41 42 49 58
rect 51 54 59 70
rect 51 50 53 54
rect 57 50 59 54
rect 51 47 59 50
rect 51 43 53 47
rect 57 43 59 47
rect 51 42 59 43
rect 61 69 69 70
rect 61 65 63 69
rect 67 65 69 69
rect 61 62 69 65
rect 61 58 63 62
rect 67 58 69 62
rect 61 42 69 58
rect 71 54 79 70
rect 71 50 73 54
rect 77 50 79 54
rect 71 47 79 50
rect 71 43 73 47
rect 77 43 79 47
rect 71 42 79 43
rect 81 69 89 70
rect 81 65 83 69
rect 87 65 89 69
rect 81 62 89 65
rect 81 58 83 62
rect 87 58 89 62
rect 81 42 89 58
rect 91 54 99 70
rect 91 50 93 54
rect 97 50 99 54
rect 91 47 99 50
rect 91 43 93 47
rect 97 43 99 47
rect 91 42 99 43
rect 101 69 109 70
rect 101 65 103 69
rect 107 65 109 69
rect 101 62 109 65
rect 101 58 103 62
rect 107 58 109 62
rect 101 42 109 58
rect 111 62 119 70
rect 111 58 113 62
rect 117 58 119 62
rect 111 55 119 58
rect 111 51 113 55
rect 117 51 119 55
rect 111 42 119 51
rect 121 69 128 70
rect 121 65 123 69
rect 127 65 128 69
rect 121 62 128 65
rect 121 58 123 62
rect 127 58 128 62
rect 121 42 128 58
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect 118 78 122 82
rect 126 78 130 82
rect 134 78 138 82
rect 142 78 146 82
rect -2 69 146 78
rect -2 68 43 69
rect 42 65 43 68
rect 47 68 63 69
rect 47 65 48 68
rect 2 54 7 63
rect 42 62 48 65
rect 2 50 3 54
rect 12 58 13 62
rect 17 58 33 62
rect 37 58 38 62
rect 42 58 43 62
rect 47 58 48 62
rect 62 65 63 68
rect 67 68 83 69
rect 67 65 68 68
rect 62 62 68 65
rect 62 58 63 62
rect 67 58 68 62
rect 82 65 83 68
rect 87 68 103 69
rect 87 65 88 68
rect 82 62 88 65
rect 82 58 83 62
rect 87 58 88 62
rect 102 65 103 68
rect 107 68 123 69
rect 107 65 108 68
rect 102 62 108 65
rect 122 65 123 68
rect 127 68 146 69
rect 127 65 128 68
rect 102 58 103 62
rect 107 58 108 62
rect 113 62 117 63
rect 122 62 128 65
rect 122 58 123 62
rect 127 58 128 62
rect 12 55 18 58
rect 12 51 13 55
rect 17 51 18 55
rect 32 55 38 58
rect 2 47 7 50
rect 2 43 3 47
rect 22 50 23 54
rect 27 50 28 54
rect 32 51 33 55
rect 37 54 38 55
rect 113 55 117 58
rect 37 51 53 54
rect 32 50 53 51
rect 57 50 73 54
rect 77 50 93 54
rect 97 51 113 54
rect 97 50 117 51
rect 22 47 28 50
rect 22 46 23 47
rect 7 43 23 46
rect 27 46 28 47
rect 53 47 57 50
rect 27 43 30 46
rect 2 42 30 43
rect 2 34 10 38
rect 14 34 15 38
rect 2 17 6 34
rect 26 30 30 42
rect 41 38 47 46
rect 53 42 57 43
rect 73 47 77 50
rect 93 47 97 50
rect 73 42 77 43
rect 81 38 87 46
rect 93 42 97 43
rect 122 38 126 55
rect 41 34 44 38
rect 48 34 56 38
rect 60 34 63 38
rect 73 34 76 38
rect 80 34 84 38
rect 88 34 95 38
rect 105 34 109 38
rect 113 34 116 38
rect 120 34 126 38
rect 13 29 58 30
rect 13 26 53 29
rect 37 25 53 26
rect 57 25 58 29
rect 63 28 67 29
rect 37 22 38 25
rect 13 21 17 22
rect 23 21 27 22
rect 33 17 38 22
rect 72 25 73 29
rect 77 25 93 29
rect 97 28 117 29
rect 97 25 113 28
rect 63 21 67 24
rect 93 22 97 25
rect 42 17 43 21
rect 47 17 63 21
rect 67 17 83 21
rect 87 17 88 21
rect 113 21 117 24
rect 93 17 97 18
rect 103 17 107 18
rect 23 12 27 17
rect 113 16 117 17
rect 123 25 127 26
rect 123 17 127 21
rect 103 12 107 13
rect 123 12 127 13
rect -2 2 146 12
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 122 2
rect 126 -2 130 2
rect 134 -2 138 2
rect 142 -2 146 2
<< ntransistor >>
rect 19 16 21 27
rect 29 16 31 27
rect 39 12 41 30
rect 49 12 51 30
rect 59 12 61 30
rect 69 12 71 30
rect 79 12 81 30
rect 89 12 91 30
rect 99 12 101 30
rect 109 12 111 30
rect 119 12 121 30
<< ptransistor >>
rect 9 42 11 70
rect 19 42 21 70
rect 29 42 31 70
rect 39 42 41 70
rect 49 42 51 70
rect 59 42 61 70
rect 69 42 71 70
rect 79 42 81 70
rect 89 42 91 70
rect 99 42 101 70
rect 109 42 111 70
rect 119 42 121 70
<< polycontact >>
rect 10 34 14 38
rect 44 34 48 38
rect 56 34 60 38
rect 76 34 80 38
rect 84 34 88 38
rect 109 34 113 38
rect 116 34 120 38
<< ndcontact >>
rect 13 22 17 26
rect 23 17 27 21
rect 33 22 37 26
rect 43 17 47 21
rect 53 25 57 29
rect 63 24 67 28
rect 63 17 67 21
rect 73 25 77 29
rect 83 17 87 21
rect 93 25 97 29
rect 93 18 97 22
rect 103 13 107 17
rect 113 24 117 28
rect 113 17 117 21
rect 123 21 127 25
rect 123 13 127 17
<< pdcontact >>
rect 3 50 7 54
rect 3 43 7 47
rect 13 58 17 62
rect 13 51 17 55
rect 23 50 27 54
rect 23 43 27 47
rect 33 58 37 62
rect 33 51 37 55
rect 43 65 47 69
rect 43 58 47 62
rect 53 50 57 54
rect 53 43 57 47
rect 63 65 67 69
rect 63 58 67 62
rect 73 50 77 54
rect 73 43 77 47
rect 83 65 87 69
rect 83 58 87 62
rect 93 50 97 54
rect 93 43 97 47
rect 103 65 107 69
rect 103 58 107 62
rect 113 58 117 62
rect 113 51 117 55
rect 123 65 127 69
rect 123 58 127 62
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
rect 90 -2 94 2
rect 98 -2 102 2
rect 106 -2 110 2
rect 114 -2 118 2
rect 122 -2 126 2
rect 130 -2 134 2
rect 138 -2 142 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
rect 90 78 94 82
rect 98 78 102 82
rect 106 78 110 82
rect 114 78 118 82
rect 122 78 126 82
rect 130 78 134 82
rect 138 78 142 82
<< psubstratepdiff >>
rect 0 2 144 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 122 2
rect 126 -2 130 2
rect 134 -2 138 2
rect 142 -2 144 2
rect 0 -3 144 -2
<< nsubstratendiff >>
rect 0 82 144 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect 118 78 122 82
rect 126 78 130 82
rect 134 78 138 82
rect 142 78 144 82
rect 0 77 144 78
<< labels >>
rlabel metal1 20 28 20 28 6 z
rlabel metal1 4 24 4 24 6 b
rlabel polycontact 12 36 12 36 6 b
rlabel metal1 12 44 12 44 6 z
rlabel metal1 20 44 20 44 6 z
rlabel metal1 15 56 15 56 6 n3
rlabel metal1 4 56 4 56 6 z
rlabel ndcontact 36 24 36 24 6 z
rlabel metal1 44 28 44 28 6 z
rlabel metal1 52 28 52 28 6 z
rlabel metal1 28 32 28 32 6 z
rlabel metal1 44 40 44 40 6 a3
rlabel metal1 52 36 52 36 6 a3
rlabel metal1 35 56 35 56 6 n3
rlabel metal1 25 60 25 60 6 n3
rlabel metal1 72 6 72 6 6 vss
rlabel metal1 65 23 65 23 6 n2
rlabel metal1 60 36 60 36 6 a3
rlabel metal1 76 36 76 36 6 a2
rlabel metal1 84 40 84 40 6 a2
rlabel metal1 75 48 75 48 6 n3
rlabel metal1 55 48 55 48 6 n3
rlabel metal1 72 74 72 74 6 vdd
rlabel ndcontact 65 19 65 19 6 n2
rlabel metal1 95 23 95 23 6 n1
rlabel metal1 108 36 108 36 6 a1
rlabel metal1 92 36 92 36 6 a2
rlabel metal1 95 48 95 48 6 n3
rlabel metal1 115 22 115 22 6 n1
rlabel ndcontact 94 27 94 27 6 n1
rlabel metal1 116 36 116 36 6 a1
rlabel metal1 124 48 124 48 6 a1
rlabel metal1 115 56 115 56 6 n3
rlabel pdcontact 74 52 74 52 6 n3
<< end >>
