magic
tech scmos
timestamp 1182081807
<< checkpaint >>
rect -25 -26 89 114
<< ab >>
rect 0 0 64 88
<< pwell >>
rect -7 -8 71 40
<< nwell >>
rect -7 40 71 96
<< polysilicon >>
rect 5 80 14 86
rect 18 80 27 86
rect 37 80 46 86
rect 50 80 59 86
rect 9 77 11 80
rect 21 77 23 80
rect 41 77 43 80
rect 53 77 55 80
rect 9 48 11 51
rect 21 48 23 51
rect 41 48 43 51
rect 53 48 55 51
rect 2 47 11 48
rect 2 43 6 47
rect 10 43 11 47
rect 2 42 11 43
rect 15 47 30 48
rect 15 43 22 47
rect 26 43 30 47
rect 15 42 30 43
rect 34 47 43 48
rect 34 43 38 47
rect 42 43 43 47
rect 34 42 43 43
rect 47 47 62 48
rect 47 43 54 47
rect 58 43 62 47
rect 47 42 62 43
rect 2 32 17 38
rect 21 37 30 38
rect 21 33 22 37
rect 26 33 30 37
rect 21 32 30 33
rect 34 37 49 38
rect 34 33 38 37
rect 42 33 49 37
rect 34 32 49 33
rect 53 32 62 38
rect 9 29 11 32
rect 21 29 23 32
rect 41 29 43 32
rect 53 29 55 32
rect 9 8 11 11
rect 21 8 23 11
rect 41 8 43 11
rect 53 8 55 11
rect 5 7 14 8
rect 5 3 6 7
rect 10 3 14 7
rect 5 2 14 3
rect 18 2 27 8
rect 37 2 46 8
rect 50 7 59 8
rect 50 3 54 7
rect 58 3 59 7
rect 50 2 59 3
<< ndiffusion >>
rect 2 11 9 29
rect 11 24 21 29
rect 11 20 14 24
rect 18 20 21 24
rect 11 16 21 20
rect 11 12 14 16
rect 18 12 21 16
rect 11 11 21 12
rect 23 26 30 29
rect 23 22 25 26
rect 29 22 30 26
rect 23 18 30 22
rect 23 14 25 18
rect 29 14 30 18
rect 23 11 30 14
rect 34 26 41 29
rect 34 22 35 26
rect 39 22 41 26
rect 34 18 41 22
rect 34 14 35 18
rect 39 14 41 18
rect 34 11 41 14
rect 43 24 53 29
rect 43 20 46 24
rect 50 20 53 24
rect 43 17 53 20
rect 43 13 46 17
rect 50 13 53 17
rect 43 11 53 13
rect 55 11 62 29
<< pdiffusion >>
rect 2 75 9 77
rect 2 71 3 75
rect 7 71 9 75
rect 2 68 9 71
rect 2 64 3 68
rect 7 64 9 68
rect 2 51 9 64
rect 11 66 21 77
rect 11 62 14 66
rect 18 62 21 66
rect 11 59 21 62
rect 11 55 14 59
rect 18 55 21 59
rect 11 51 21 55
rect 23 75 30 77
rect 23 71 25 75
rect 29 71 30 75
rect 23 51 30 71
rect 34 75 41 77
rect 34 71 35 75
rect 39 71 41 75
rect 34 68 41 71
rect 34 64 35 68
rect 39 64 41 68
rect 34 51 41 64
rect 43 66 53 77
rect 43 62 46 66
rect 50 62 53 66
rect 43 58 53 62
rect 43 54 46 58
rect 50 54 53 58
rect 43 51 53 54
rect 55 75 62 77
rect 55 71 57 75
rect 61 71 62 75
rect 55 68 62 71
rect 55 64 57 68
rect 61 64 62 68
rect 55 51 62 64
<< metal1 >>
rect -2 86 2 90
rect 30 86 34 90
rect 2 82 30 85
rect -2 81 34 82
rect 62 86 66 90
rect 62 81 66 82
rect 3 75 7 81
rect 3 68 7 71
rect 25 75 29 81
rect 25 70 29 71
rect 35 75 61 76
rect 39 72 57 75
rect 35 68 39 71
rect 3 63 7 64
rect 14 66 35 67
rect 18 64 35 66
rect 57 68 61 71
rect 18 63 39 64
rect 46 66 50 67
rect 14 59 18 62
rect 57 63 61 64
rect 46 59 50 62
rect 14 54 18 55
rect 22 50 26 59
rect 5 47 26 50
rect 5 43 6 47
rect 10 46 22 47
rect 10 43 11 46
rect 22 37 26 43
rect 22 32 26 33
rect 30 58 50 59
rect 30 55 46 58
rect 30 26 34 55
rect 46 53 50 54
rect 38 47 42 51
rect 38 42 42 43
rect 53 43 54 47
rect 58 43 59 47
rect 53 42 59 43
rect 38 38 59 42
rect 38 37 42 38
rect 38 29 42 33
rect 14 24 18 25
rect 24 22 25 26
rect 29 22 35 26
rect 39 22 40 26
rect 46 24 50 25
rect 14 16 18 20
rect 30 18 34 22
rect 24 14 25 18
rect 29 14 35 18
rect 39 14 40 18
rect 46 17 50 20
rect 14 7 18 12
rect 46 7 50 13
rect -2 6 6 7
rect 2 3 6 6
rect 10 6 54 7
rect 10 3 30 6
rect -2 -2 2 2
rect 34 3 54 6
rect 58 6 66 7
rect 58 3 62 6
rect 30 -2 34 2
rect 62 -2 66 2
<< metal2 >>
rect -2 86 66 90
rect 2 82 30 86
rect 34 82 62 86
rect -2 80 66 82
rect -2 6 66 8
rect 2 2 30 6
rect 34 2 62 6
rect -2 -2 66 2
<< ntransistor >>
rect 9 11 11 29
rect 21 11 23 29
rect 41 11 43 29
rect 53 11 55 29
<< ptransistor >>
rect 9 51 11 77
rect 21 51 23 77
rect 41 51 43 77
rect 53 51 55 77
<< polycontact >>
rect 6 43 10 47
rect 22 43 26 47
rect 38 43 42 47
rect 54 43 58 47
rect 22 33 26 37
rect 38 33 42 37
rect 6 3 10 7
rect 54 3 58 7
<< ndcontact >>
rect 14 20 18 24
rect 14 12 18 16
rect 25 22 29 26
rect 25 14 29 18
rect 35 22 39 26
rect 35 14 39 18
rect 46 20 50 24
rect 46 13 50 17
<< pdcontact >>
rect 3 71 7 75
rect 3 64 7 68
rect 14 62 18 66
rect 14 55 18 59
rect 25 71 29 75
rect 35 71 39 75
rect 35 64 39 68
rect 46 62 50 66
rect 46 54 50 58
rect 57 71 61 75
rect 57 64 61 68
<< m2contact >>
rect -2 82 2 86
rect 30 82 34 86
rect 62 82 66 86
rect -2 2 2 6
rect 30 2 34 6
rect 62 2 66 6
<< psubstratepcontact >>
rect -2 2 2 6
rect 30 2 34 6
rect 62 2 66 6
<< nsubstratencontact >>
rect -2 82 2 86
rect 30 82 34 86
rect 62 82 66 86
<< psubstratepdiff >>
rect -3 6 3 7
rect -3 2 -2 6
rect 2 2 3 6
rect 29 6 35 7
rect 29 2 30 6
rect 34 2 35 6
rect 61 6 67 7
rect 61 2 62 6
rect 66 2 67 6
rect -3 0 3 2
rect 29 0 35 2
rect 61 0 67 2
<< nsubstratendiff >>
rect -3 86 3 88
rect 29 86 35 88
rect 61 86 67 88
rect -3 82 -2 86
rect 2 82 3 86
rect -3 81 3 82
rect 29 82 30 86
rect 34 82 35 86
rect 29 81 35 82
rect 61 82 62 86
rect 66 82 67 86
rect 61 81 67 82
<< labels >>
rlabel metal1 8 48 8 48 6 a
rlabel metal1 24 48 24 48 6 a
rlabel metal1 16 48 16 48 6 a
rlabel metal1 32 36 32 36 6 z
rlabel metal1 40 40 40 40 6 b
rlabel metal1 48 40 48 40 6 b
rlabel metal1 56 40 56 40 6 b
rlabel metal1 48 60 48 60 6 z
rlabel m2contact 32 4 32 4 6 vss
rlabel m2contact 32 84 32 84 6 vdd
<< end >>
