magic
tech scmos
timestamp 1185039065
<< checkpaint >>
rect -22 -24 192 124
<< ab >>
rect 0 0 170 100
<< pwell >>
rect -2 -4 172 49
<< nwell >>
rect -2 49 172 104
<< polysilicon >>
rect 11 95 13 98
rect 23 95 25 98
rect 47 95 49 98
rect 59 95 61 98
rect 71 95 73 98
rect 83 95 85 98
rect 109 95 111 98
rect 121 95 123 98
rect 133 95 135 98
rect 145 95 147 98
rect 157 75 159 78
rect 11 53 13 55
rect 7 52 13 53
rect 7 48 8 52
rect 12 48 13 52
rect 7 47 13 48
rect 11 25 13 47
rect 23 53 25 55
rect 47 53 49 55
rect 59 53 61 55
rect 71 53 73 55
rect 83 53 85 55
rect 23 52 33 53
rect 23 48 28 52
rect 32 48 33 52
rect 23 47 33 48
rect 47 52 53 53
rect 47 48 48 52
rect 52 48 53 52
rect 47 47 53 48
rect 57 52 63 53
rect 57 48 58 52
rect 62 48 63 52
rect 57 47 63 48
rect 67 52 73 53
rect 67 48 68 52
rect 72 48 73 52
rect 67 47 73 48
rect 77 52 85 53
rect 77 48 78 52
rect 82 51 85 52
rect 82 48 83 51
rect 77 47 83 48
rect 23 25 25 47
rect 51 25 53 47
rect 59 25 61 47
rect 71 25 73 47
rect 79 25 81 47
rect 109 43 111 55
rect 121 43 123 55
rect 107 42 113 43
rect 107 38 108 42
rect 112 38 113 42
rect 107 37 113 38
rect 121 42 127 43
rect 121 38 122 42
rect 126 38 127 42
rect 121 37 127 38
rect 133 41 135 55
rect 145 43 147 55
rect 145 42 153 43
rect 145 41 148 42
rect 133 39 148 41
rect 109 29 111 37
rect 109 27 115 29
rect 113 25 115 27
rect 121 25 123 37
rect 133 25 135 39
rect 145 38 148 39
rect 152 38 153 42
rect 145 37 153 38
rect 145 25 147 37
rect 157 33 159 55
rect 151 32 159 33
rect 151 28 152 32
rect 156 28 159 32
rect 151 27 159 28
rect 157 25 159 27
rect 157 12 159 15
rect 11 2 13 5
rect 23 2 25 5
rect 51 2 53 5
rect 59 2 61 5
rect 71 2 73 5
rect 79 2 81 5
rect 113 2 115 5
rect 121 2 123 5
rect 133 2 135 5
rect 145 2 147 5
<< ndiffusion >>
rect 137 32 143 33
rect 137 28 138 32
rect 142 28 143 32
rect 137 25 143 28
rect 3 12 11 25
rect 3 8 4 12
rect 8 8 11 12
rect 3 5 11 8
rect 13 5 23 25
rect 25 22 33 25
rect 25 18 28 22
rect 32 18 33 22
rect 25 5 33 18
rect 43 12 51 25
rect 43 8 44 12
rect 48 8 51 12
rect 43 5 51 8
rect 53 5 59 25
rect 61 22 71 25
rect 61 18 64 22
rect 68 18 71 22
rect 61 5 71 18
rect 73 5 79 25
rect 81 12 89 25
rect 81 8 84 12
rect 88 8 89 12
rect 81 5 89 8
rect 105 22 113 25
rect 105 18 106 22
rect 110 18 113 22
rect 105 5 113 18
rect 115 5 121 25
rect 123 12 133 25
rect 123 8 126 12
rect 130 8 133 12
rect 123 5 133 8
rect 135 5 145 25
rect 147 15 157 25
rect 159 22 167 25
rect 159 18 162 22
rect 166 18 167 22
rect 159 15 167 18
rect 147 12 155 15
rect 147 8 150 12
rect 154 8 155 12
rect 147 5 155 8
<< pdiffusion >>
rect 3 82 11 95
rect 3 78 4 82
rect 8 78 11 82
rect 3 72 11 78
rect 3 68 4 72
rect 8 68 11 72
rect 3 55 11 68
rect 13 72 23 95
rect 13 68 16 72
rect 20 68 23 72
rect 13 55 23 68
rect 25 82 33 95
rect 25 78 28 82
rect 32 78 33 82
rect 25 72 33 78
rect 25 68 28 72
rect 32 68 33 72
rect 25 55 33 68
rect 39 82 47 95
rect 39 78 40 82
rect 44 78 47 82
rect 39 55 47 78
rect 49 72 59 95
rect 49 68 52 72
rect 56 68 59 72
rect 49 55 59 68
rect 61 82 71 95
rect 61 78 64 82
rect 68 78 71 82
rect 61 72 71 78
rect 61 68 64 72
rect 68 68 71 72
rect 61 55 71 68
rect 73 72 83 95
rect 73 68 76 72
rect 80 68 83 72
rect 73 55 83 68
rect 85 82 93 95
rect 85 78 88 82
rect 92 78 93 82
rect 85 55 93 78
rect 101 92 109 95
rect 101 88 102 92
rect 106 88 109 92
rect 101 82 109 88
rect 101 78 102 82
rect 106 78 109 82
rect 101 55 109 78
rect 111 82 121 95
rect 111 78 114 82
rect 118 78 121 82
rect 111 55 121 78
rect 123 92 133 95
rect 123 88 126 92
rect 130 88 133 92
rect 123 82 133 88
rect 123 78 126 82
rect 130 78 133 82
rect 123 55 133 78
rect 135 82 145 95
rect 135 78 138 82
rect 142 78 145 82
rect 135 72 145 78
rect 135 68 138 72
rect 142 68 145 72
rect 135 62 145 68
rect 135 58 138 62
rect 142 58 145 62
rect 135 55 145 58
rect 147 92 155 95
rect 147 88 150 92
rect 154 88 155 92
rect 147 82 155 88
rect 147 78 150 82
rect 154 78 155 82
rect 147 75 155 78
rect 147 72 157 75
rect 147 68 150 72
rect 154 68 157 72
rect 147 55 157 68
rect 159 72 167 75
rect 159 68 162 72
rect 166 68 167 72
rect 159 60 167 68
rect 159 56 162 60
rect 166 56 167 60
rect 159 55 167 56
<< metal1 >>
rect -2 94 172 101
rect -2 92 162 94
rect -2 88 102 92
rect 106 88 126 92
rect 130 88 150 92
rect 154 90 162 92
rect 166 90 172 94
rect 154 88 172 90
rect -2 87 172 88
rect 3 82 9 83
rect 27 82 33 83
rect 3 78 4 82
rect 8 78 28 82
rect 32 78 33 82
rect 3 77 9 78
rect 27 77 33 78
rect 39 82 45 83
rect 63 82 69 83
rect 87 82 93 83
rect 39 78 40 82
rect 44 78 64 82
rect 68 78 88 82
rect 92 78 93 82
rect 39 77 45 78
rect 63 77 69 78
rect 87 77 93 78
rect 101 82 107 87
rect 101 78 102 82
rect 106 78 107 82
rect 101 77 107 78
rect 113 82 119 83
rect 113 78 114 82
rect 118 78 119 82
rect 113 77 119 78
rect 125 82 131 87
rect 125 78 126 82
rect 130 78 131 82
rect 125 77 131 78
rect 137 82 143 83
rect 137 78 138 82
rect 142 78 143 82
rect 4 73 8 77
rect 28 73 32 77
rect 64 73 68 77
rect 3 72 9 73
rect 3 68 4 72
rect 8 68 9 72
rect 3 67 9 68
rect 15 72 21 73
rect 27 72 33 73
rect 51 72 57 73
rect 15 68 16 72
rect 20 68 22 72
rect 15 67 22 68
rect 27 68 28 72
rect 32 68 52 72
rect 56 68 57 72
rect 27 67 33 68
rect 51 67 57 68
rect 63 72 69 73
rect 63 68 64 72
rect 68 68 69 72
rect 63 67 69 68
rect 75 72 81 73
rect 114 72 118 77
rect 137 72 143 78
rect 75 68 76 72
rect 80 68 118 72
rect 75 67 81 68
rect 7 52 13 62
rect 7 48 8 52
rect 12 48 13 52
rect 7 18 13 48
rect 18 22 22 67
rect 27 52 33 62
rect 27 48 28 52
rect 32 48 33 52
rect 27 28 33 48
rect 47 52 53 62
rect 47 48 48 52
rect 52 48 53 52
rect 47 28 53 48
rect 57 52 63 62
rect 57 48 58 52
rect 62 48 63 52
rect 57 28 63 48
rect 67 52 73 62
rect 67 48 68 52
rect 72 48 73 52
rect 67 28 73 48
rect 77 52 83 62
rect 77 48 78 52
rect 82 48 83 52
rect 77 28 83 48
rect 107 42 113 62
rect 127 43 133 72
rect 107 38 108 42
rect 112 38 113 42
rect 107 28 113 38
rect 121 42 133 43
rect 121 38 122 42
rect 126 38 133 42
rect 121 37 133 38
rect 127 28 133 37
rect 137 68 138 72
rect 142 68 143 72
rect 137 62 143 68
rect 149 82 155 87
rect 149 78 150 82
rect 154 78 155 82
rect 149 72 155 78
rect 149 68 150 72
rect 154 68 155 72
rect 149 67 155 68
rect 161 72 167 73
rect 161 68 162 72
rect 166 68 167 72
rect 161 67 167 68
rect 137 58 138 62
rect 142 58 143 62
rect 162 61 166 67
rect 137 32 143 58
rect 161 60 167 61
rect 161 56 162 60
rect 166 56 167 60
rect 161 55 167 56
rect 147 42 153 43
rect 162 42 166 55
rect 147 38 148 42
rect 152 38 166 42
rect 147 37 153 38
rect 137 28 138 32
rect 142 28 143 32
rect 137 27 143 28
rect 151 32 157 33
rect 151 28 152 32
rect 156 28 157 32
rect 151 27 157 28
rect 27 22 33 23
rect 63 22 69 23
rect 105 22 111 23
rect 152 22 156 27
rect 162 23 166 38
rect 18 18 28 22
rect 32 18 64 22
rect 68 18 106 22
rect 110 18 156 22
rect 161 22 167 23
rect 161 18 162 22
rect 166 18 167 22
rect 27 17 33 18
rect 63 17 69 18
rect 105 17 111 18
rect 161 17 167 18
rect -2 12 172 13
rect -2 8 4 12
rect 8 8 44 12
rect 48 8 84 12
rect 88 8 126 12
rect 130 8 150 12
rect 154 8 172 12
rect -2 -1 172 8
<< ntransistor >>
rect 11 5 13 25
rect 23 5 25 25
rect 51 5 53 25
rect 59 5 61 25
rect 71 5 73 25
rect 79 5 81 25
rect 113 5 115 25
rect 121 5 123 25
rect 133 5 135 25
rect 145 5 147 25
rect 157 15 159 25
<< ptransistor >>
rect 11 55 13 95
rect 23 55 25 95
rect 47 55 49 95
rect 59 55 61 95
rect 71 55 73 95
rect 83 55 85 95
rect 109 55 111 95
rect 121 55 123 95
rect 133 55 135 95
rect 145 55 147 95
rect 157 55 159 75
<< polycontact >>
rect 8 48 12 52
rect 28 48 32 52
rect 48 48 52 52
rect 58 48 62 52
rect 68 48 72 52
rect 78 48 82 52
rect 108 38 112 42
rect 122 38 126 42
rect 148 38 152 42
rect 152 28 156 32
<< ndcontact >>
rect 138 28 142 32
rect 4 8 8 12
rect 28 18 32 22
rect 44 8 48 12
rect 64 18 68 22
rect 84 8 88 12
rect 106 18 110 22
rect 126 8 130 12
rect 162 18 166 22
rect 150 8 154 12
<< pdcontact >>
rect 4 78 8 82
rect 4 68 8 72
rect 16 68 20 72
rect 28 78 32 82
rect 28 68 32 72
rect 40 78 44 82
rect 52 68 56 72
rect 64 78 68 82
rect 64 68 68 72
rect 76 68 80 72
rect 88 78 92 82
rect 102 88 106 92
rect 102 78 106 82
rect 114 78 118 82
rect 126 88 130 92
rect 126 78 130 82
rect 138 78 142 82
rect 138 68 142 72
rect 138 58 142 62
rect 150 88 154 92
rect 150 78 154 82
rect 150 68 154 72
rect 162 68 166 72
rect 162 56 166 60
<< nsubstratencontact >>
rect 162 90 166 94
<< nsubstratendiff >>
rect 161 94 167 95
rect 161 90 162 94
rect 166 90 167 94
rect 161 83 167 90
<< labels >>
rlabel metal1 10 40 10 40 6 i7
rlabel metal1 10 40 10 40 6 i7
rlabel metal1 30 45 30 45 6 i6
rlabel metal1 30 45 30 45 6 i6
rlabel metal1 60 45 60 45 6 i4
rlabel metal1 50 45 50 45 6 i5
rlabel metal1 60 45 60 45 6 i4
rlabel metal1 50 45 50 45 6 i5
rlabel metal1 85 6 85 6 6 vss
rlabel metal1 85 6 85 6 6 vss
rlabel metal1 70 45 70 45 6 i3
rlabel metal1 70 45 70 45 6 i3
rlabel metal1 80 45 80 45 6 i2
rlabel metal1 80 45 80 45 6 i2
rlabel metal1 85 94 85 94 6 vdd
rlabel metal1 85 94 85 94 6 vdd
rlabel metal1 130 50 130 50 6 i0
rlabel metal1 110 45 110 45 6 i1
rlabel metal1 110 45 110 45 6 i1
rlabel metal1 130 50 130 50 6 i0
rlabel metal1 140 55 140 55 6 nq
rlabel metal1 140 55 140 55 6 nq
<< end >>
