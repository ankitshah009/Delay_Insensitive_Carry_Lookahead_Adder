magic
tech scmos
timestamp 1179386169
<< checkpaint >>
rect -22 -22 78 94
<< ab >>
rect 0 0 56 72
<< pwell >>
rect -4 -4 60 32
<< nwell >>
rect -4 32 60 76
<< polysilicon >>
rect 9 59 11 64
rect 22 59 24 64
rect 32 59 34 64
rect 44 57 46 61
rect 9 33 11 47
rect 22 43 24 47
rect 16 42 24 43
rect 16 38 17 42
rect 21 38 24 42
rect 16 37 24 38
rect 9 32 15 33
rect 9 28 10 32
rect 14 28 15 32
rect 9 27 15 28
rect 22 27 24 37
rect 32 36 34 47
rect 44 42 46 45
rect 41 41 47 42
rect 41 37 42 41
rect 46 37 47 41
rect 41 36 47 37
rect 32 34 37 36
rect 35 32 37 34
rect 35 31 41 32
rect 35 27 36 31
rect 40 27 41 31
rect 9 22 11 27
rect 22 25 30 27
rect 28 22 30 25
rect 35 26 41 27
rect 35 22 37 26
rect 45 22 47 36
rect 9 11 11 16
rect 28 7 30 12
rect 35 7 37 12
rect 45 11 47 16
<< ndiffusion >>
rect 2 21 9 22
rect 2 17 3 21
rect 7 17 9 21
rect 2 16 9 17
rect 11 16 17 22
rect 23 20 28 22
rect 13 10 17 16
rect 21 19 28 20
rect 21 15 22 19
rect 26 15 28 19
rect 21 14 28 15
rect 23 12 28 14
rect 30 12 35 22
rect 37 21 45 22
rect 37 17 39 21
rect 43 17 45 21
rect 37 16 45 17
rect 47 21 54 22
rect 47 17 49 21
rect 53 17 54 21
rect 47 16 54 17
rect 37 12 43 16
rect 13 8 19 10
rect 13 4 14 8
rect 18 4 19 8
rect 13 3 19 4
<< pdiffusion >>
rect 4 53 9 59
rect 2 52 9 53
rect 2 48 3 52
rect 7 48 9 52
rect 2 47 9 48
rect 11 58 22 59
rect 11 54 15 58
rect 19 54 22 58
rect 11 47 22 54
rect 24 53 32 59
rect 24 49 26 53
rect 30 49 32 53
rect 24 47 32 49
rect 34 58 42 59
rect 34 54 36 58
rect 40 57 42 58
rect 40 54 44 57
rect 34 47 44 54
rect 36 45 44 47
rect 46 51 51 57
rect 46 50 53 51
rect 46 46 48 50
rect 52 46 53 50
rect 46 45 53 46
<< metal1 >>
rect -2 68 58 72
rect -2 64 41 68
rect 45 64 48 68
rect 52 64 58 68
rect 15 58 19 64
rect 15 53 19 54
rect 26 53 30 59
rect 35 58 41 64
rect 35 54 36 58
rect 40 54 41 58
rect 3 52 7 53
rect 3 42 7 48
rect 2 38 17 42
rect 21 38 22 42
rect 2 22 6 38
rect 10 32 22 35
rect 14 29 22 32
rect 2 21 7 22
rect 2 17 3 21
rect 2 16 7 17
rect 10 13 14 28
rect 18 15 22 19
rect 26 15 30 49
rect 34 43 38 51
rect 47 46 48 50
rect 52 46 54 50
rect 34 41 47 43
rect 34 37 42 41
rect 46 37 47 41
rect 50 31 54 46
rect 35 27 36 31
rect 40 27 54 31
rect 50 22 54 27
rect 18 13 30 15
rect 39 21 43 22
rect 39 8 43 17
rect 49 21 54 22
rect 53 17 54 21
rect 49 16 54 17
rect -2 4 4 8
rect 8 4 14 8
rect 18 4 48 8
rect 52 4 58 8
rect -2 0 58 4
<< ntransistor >>
rect 9 16 11 22
rect 28 12 30 22
rect 35 12 37 22
rect 45 16 47 22
<< ptransistor >>
rect 9 47 11 59
rect 22 47 24 59
rect 32 47 34 59
rect 44 45 46 57
<< polycontact >>
rect 17 38 21 42
rect 10 28 14 32
rect 42 37 46 41
rect 36 27 40 31
<< ndcontact >>
rect 3 17 7 21
rect 22 15 26 19
rect 39 17 43 21
rect 49 17 53 21
rect 14 4 18 8
<< pdcontact >>
rect 3 48 7 52
rect 15 54 19 58
rect 26 49 30 53
rect 36 54 40 58
rect 48 46 52 50
<< psubstratepcontact >>
rect 4 4 8 8
rect 48 4 52 8
<< nsubstratencontact >>
rect 41 64 45 68
rect 48 64 52 68
<< psubstratepdiff >>
rect 3 8 9 9
rect 3 4 4 8
rect 8 4 9 8
rect 3 3 9 4
rect 47 8 53 9
rect 47 4 48 8
rect 52 4 53 8
rect 47 3 53 4
<< nsubstratendiff >>
rect 40 68 53 69
rect 40 64 41 68
rect 45 64 48 68
rect 52 64 53 68
rect 40 63 53 64
<< labels >>
rlabel polycontact 20 40 20 40 6 bn
rlabel polycontact 38 29 38 29 6 an
rlabel metal1 5 45 5 45 6 bn
rlabel metal1 4 29 4 29 6 bn
rlabel metal1 20 16 20 16 6 z
rlabel metal1 12 24 12 24 6 b
rlabel metal1 20 32 20 32 6 b
rlabel metal1 12 40 12 40 6 bn
rlabel metal1 28 4 28 4 6 vss
rlabel metal1 28 36 28 36 6 z
rlabel metal1 36 44 36 44 6 a
rlabel metal1 28 68 28 68 6 vdd
rlabel metal1 44 29 44 29 6 an
rlabel polycontact 44 40 44 40 6 a
rlabel metal1 52 33 52 33 6 an
rlabel pdcontact 50 48 50 48 6 an
<< end >>
