.subckt nao2o22_x4 i0 i1 i2 i3 nq vdd vss
*   SPICE3 file   created from nao2o22_x4.ext -      technology: scmos
m00 w1     i0     vdd    vdd p w=20u  l=2.3636u ad=100p     pd=30u      as=156.571p ps=48.5714u
m01 w2     i1     w1     vdd p w=20u  l=2.3636u ad=100p     pd=30u      as=100p     ps=30u
m02 w3     i3     w2     vdd p w=20u  l=2.3636u ad=100p     pd=30u      as=100p     ps=30u
m03 vdd    i2     w3     vdd p w=20u  l=2.3636u ad=156.571p pd=48.5714u as=100p     ps=30u
m04 vdd    w2     w4     vdd p w=20u  l=2.3636u ad=156.571p pd=48.5714u as=160p     ps=56u
m05 nq     w4     vdd    vdd p w=40u  l=2.3636u ad=200p     pd=50u      as=313.143p ps=97.1429u
m06 vdd    w4     nq     vdd p w=40u  l=2.3636u ad=313.143p pd=97.1429u as=200p     ps=50u
m07 w2     i0     w5     vss n w=10u  l=2.3636u ad=74p      pd=28u      as=65p      ps=28u
m08 w5     i1     w2     vss n w=10u  l=2.3636u ad=65p      pd=28u      as=74p      ps=28u
m09 vss    i3     w5     vss n w=10u  l=2.3636u ad=69.7143p pd=24.5714u as=65p      ps=28u
m10 w5     i2     vss    vss n w=10u  l=2.3636u ad=65p      pd=28u      as=69.7143p ps=24.5714u
m11 vss    w2     w4     vss n w=10u  l=2.3636u ad=69.7143p pd=24.5714u as=80p      ps=36u
m12 nq     w4     vss    vss n w=20u  l=2.3636u ad=100p     pd=30u      as=139.429p ps=49.1429u
m13 vss    w4     nq     vss n w=20u  l=2.3636u ad=139.429p pd=49.1429u as=100p     ps=30u
C0  w5     i0     0.018f
C1  w2     i2     0.194f
C2  w3     i3     0.016f
C3  vss    vdd    0.005f
C4  vss    nq     0.130f
C5  w4     i2     0.117f
C6  w2     i1     0.345f
C7  nq     vdd    0.231f
C8  vss    w2     0.050f
C9  w1     i0     0.009f
C10 w2     vdd    0.415f
C11 w4     i1     0.019f
C12 i2     i3     0.425f
C13 nq     w2     0.103f
C14 vss    w4     0.120f
C15 i2     i0     0.054f
C16 w4     vdd    0.031f
C17 i3     i1     0.152f
C18 nq     w4     0.132f
C19 w5     i2     0.038f
C20 vss    i3     0.015f
C21 i1     i0     0.432f
C22 i3     vdd    0.017f
C23 w2     w4     0.339f
C24 w5     i1     0.017f
C25 w3     i2     0.004f
C26 vss    i0     0.011f
C27 i0     vdd    0.065f
C28 vss    w5     0.409f
C29 w2     i3     0.355f
C30 w5     nq     0.006f
C31 w4     i3     0.056f
C32 w1     i1     0.035f
C33 w2     i0     0.093f
C34 w5     w2     0.117f
C35 i2     i1     0.079f
C36 w3     w2     0.019f
C37 w5     w4     0.032f
C38 vss    i2     0.015f
C39 i2     vdd    0.027f
C40 i3     i0     0.079f
C41 vss    i1     0.011f
C42 w5     i3     0.036f
C43 nq     i2     0.039f
C44 i1     vdd    0.042f
C46 nq     vss    0.018f
C47 w2     vss    0.051f
C48 w4     vss    0.069f
C49 i2     vss    0.040f
C50 i3     vss    0.050f
C51 i1     vss    0.043f
C52 i0     vss    0.035f
.ends
