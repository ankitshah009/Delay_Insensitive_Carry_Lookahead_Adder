magic
tech scmos
timestamp 1179385277
<< checkpaint >>
rect -22 -22 94 94
<< ab >>
rect 0 0 72 72
<< pwell >>
rect -4 -4 76 32
<< nwell >>
rect -4 32 76 76
<< polysilicon >>
rect 9 66 11 70
rect 19 66 21 70
rect 29 66 31 70
rect 39 66 41 70
rect 51 66 53 70
rect 61 66 63 70
rect 9 36 11 39
rect 9 35 15 36
rect 9 31 10 35
rect 14 31 15 35
rect 9 30 15 31
rect 19 35 21 39
rect 29 35 31 39
rect 19 34 31 35
rect 39 36 41 39
rect 51 36 53 39
rect 61 36 63 39
rect 39 34 54 36
rect 19 30 26 34
rect 30 30 31 34
rect 41 30 42 34
rect 46 30 54 34
rect 58 35 64 36
rect 58 31 59 35
rect 63 31 64 35
rect 58 30 64 31
rect 19 29 31 30
rect 20 25 22 29
rect 35 25 37 30
rect 41 29 54 30
rect 42 25 44 29
rect 52 25 54 29
rect 59 25 61 30
rect 20 5 22 10
rect 35 4 37 12
rect 42 8 44 12
rect 52 8 54 12
rect 59 4 61 12
rect 35 2 61 4
<< ndiffusion >>
rect 15 19 20 25
rect 13 18 20 19
rect 13 14 14 18
rect 18 14 20 18
rect 13 13 20 14
rect 15 10 20 13
rect 22 12 35 25
rect 37 12 42 25
rect 44 18 52 25
rect 44 14 46 18
rect 50 14 52 18
rect 44 12 52 14
rect 54 12 59 25
rect 61 12 69 25
rect 22 11 33 12
rect 22 10 26 11
rect 24 7 26 10
rect 30 7 33 11
rect 24 6 33 7
rect 63 8 69 12
rect 63 4 64 8
rect 68 4 69 8
rect 63 3 69 4
<< pdiffusion >>
rect 43 68 49 69
rect 43 66 44 68
rect 2 65 9 66
rect 2 61 3 65
rect 7 61 9 65
rect 2 58 9 61
rect 2 54 3 58
rect 7 54 9 58
rect 2 39 9 54
rect 11 59 19 66
rect 11 55 13 59
rect 17 55 19 59
rect 11 39 19 55
rect 21 50 29 66
rect 21 46 23 50
rect 27 46 29 50
rect 21 39 29 46
rect 31 58 39 66
rect 31 54 33 58
rect 37 54 39 58
rect 31 51 39 54
rect 31 47 33 51
rect 37 47 39 51
rect 31 39 39 47
rect 41 64 44 66
rect 48 66 49 68
rect 48 64 51 66
rect 41 39 51 64
rect 53 58 61 66
rect 53 54 55 58
rect 59 54 61 58
rect 53 51 61 54
rect 53 47 55 51
rect 59 47 61 51
rect 53 39 61 47
rect 63 65 70 66
rect 63 61 65 65
rect 69 61 70 65
rect 63 57 70 61
rect 63 53 65 57
rect 69 53 70 57
rect 63 39 70 53
<< metal1 >>
rect -2 68 74 72
rect -2 65 44 68
rect -2 64 3 65
rect 2 61 3 64
rect 7 64 44 65
rect 48 65 74 68
rect 48 64 65 65
rect 7 61 8 64
rect 2 58 8 61
rect 69 64 74 65
rect 2 54 3 58
rect 7 54 8 58
rect 12 55 13 59
rect 17 58 59 59
rect 17 55 33 58
rect 37 55 55 58
rect 33 51 37 54
rect 55 51 59 54
rect 65 57 69 61
rect 65 52 69 53
rect 2 50 28 51
rect 2 46 23 50
rect 27 46 28 50
rect 33 46 37 47
rect 2 18 6 46
rect 42 42 46 51
rect 55 46 59 47
rect 10 38 63 42
rect 10 35 14 38
rect 57 35 63 38
rect 10 30 14 31
rect 25 30 26 34
rect 30 30 31 34
rect 25 26 31 30
rect 17 22 31 26
rect 41 30 42 34
rect 46 30 47 34
rect 57 31 59 35
rect 57 30 63 31
rect 41 26 47 30
rect 41 22 55 26
rect 2 14 14 18
rect 18 14 46 18
rect 50 14 55 18
rect 25 8 26 11
rect -2 4 4 8
rect 8 7 26 8
rect 30 8 31 11
rect 30 7 64 8
rect 8 4 64 7
rect 68 4 74 8
rect -2 0 74 4
<< ntransistor >>
rect 20 10 22 25
rect 35 12 37 25
rect 42 12 44 25
rect 52 12 54 25
rect 59 12 61 25
<< ptransistor >>
rect 9 39 11 66
rect 19 39 21 66
rect 29 39 31 66
rect 39 39 41 66
rect 51 39 53 66
rect 61 39 63 66
<< polycontact >>
rect 10 31 14 35
rect 26 30 30 34
rect 42 30 46 34
rect 59 31 63 35
<< ndcontact >>
rect 14 14 18 18
rect 46 14 50 18
rect 26 7 30 11
rect 64 4 68 8
<< pdcontact >>
rect 3 61 7 65
rect 3 54 7 58
rect 13 55 17 59
rect 23 46 27 50
rect 33 54 37 58
rect 33 47 37 51
rect 44 64 48 68
rect 55 54 59 58
rect 55 47 59 51
rect 65 61 69 65
rect 65 53 69 57
<< psubstratepcontact >>
rect 4 4 8 8
<< psubstratepdiff >>
rect 3 8 9 24
rect 3 4 4 8
rect 8 4 9 8
rect 3 3 9 4
<< labels >>
rlabel metal1 4 36 4 36 6 z
rlabel metal1 20 16 20 16 6 z
rlabel metal1 12 16 12 16 6 z
rlabel metal1 20 24 20 24 6 b
rlabel metal1 20 40 20 40 6 a1
rlabel metal1 12 48 12 48 6 z
rlabel metal1 20 48 20 48 6 z
rlabel metal1 36 4 36 4 6 vss
rlabel metal1 36 16 36 16 6 z
rlabel metal1 28 16 28 16 6 z
rlabel metal1 28 28 28 28 6 b
rlabel metal1 28 40 28 40 6 a1
rlabel metal1 36 40 36 40 6 a1
rlabel metal1 35 52 35 52 6 n1
rlabel metal1 36 68 36 68 6 vdd
rlabel metal1 52 16 52 16 6 z
rlabel metal1 44 16 44 16 6 z
rlabel metal1 52 24 52 24 6 a2
rlabel metal1 44 28 44 28 6 a2
rlabel metal1 52 40 52 40 6 a1
rlabel metal1 44 44 44 44 6 a1
rlabel metal1 60 36 60 36 6 a1
rlabel metal1 57 52 57 52 6 n1
rlabel pdcontact 35 57 35 57 6 n1
<< end >>
