magic
tech scmos
timestamp 1179386634
<< checkpaint >>
rect -22 -22 78 94
<< ab >>
rect 0 0 56 72
<< pwell >>
rect -4 -4 60 32
<< nwell >>
rect -4 32 60 76
<< polysilicon >>
rect 9 59 11 64
rect 19 59 21 64
rect 29 59 31 64
rect 39 59 41 64
rect 9 34 11 49
rect 19 44 21 49
rect 16 43 24 44
rect 16 39 17 43
rect 21 39 24 43
rect 16 38 24 39
rect 9 33 15 34
rect 9 29 10 33
rect 14 30 15 33
rect 14 29 17 30
rect 9 28 17 29
rect 15 25 17 28
rect 22 25 24 38
rect 29 43 31 49
rect 29 42 35 43
rect 29 38 30 42
rect 34 38 35 42
rect 29 37 35 38
rect 29 25 31 37
rect 39 34 41 49
rect 39 33 47 34
rect 39 30 42 33
rect 36 29 42 30
rect 46 29 47 33
rect 36 28 47 29
rect 36 25 38 28
rect 15 8 17 13
rect 22 8 24 13
rect 29 8 31 13
rect 36 8 38 13
<< ndiffusion >>
rect 10 19 15 25
rect 8 18 15 19
rect 8 14 9 18
rect 13 14 15 18
rect 8 13 15 14
rect 17 13 22 25
rect 24 13 29 25
rect 31 13 36 25
rect 38 18 49 25
rect 38 14 43 18
rect 47 14 49 18
rect 38 13 49 14
<< pdiffusion >>
rect 2 58 9 59
rect 2 54 3 58
rect 7 54 9 58
rect 2 49 9 54
rect 11 55 19 59
rect 11 51 13 55
rect 17 51 19 55
rect 11 49 19 51
rect 21 58 29 59
rect 21 54 23 58
rect 27 54 29 58
rect 21 49 29 54
rect 31 55 39 59
rect 31 51 33 55
rect 37 51 39 55
rect 31 49 39 51
rect 41 58 49 59
rect 41 54 44 58
rect 48 54 49 58
rect 41 49 49 54
<< metal1 >>
rect -2 68 58 72
rect -2 64 48 68
rect 52 64 58 68
rect 2 58 8 64
rect 2 54 3 58
rect 7 54 8 58
rect 22 58 28 64
rect 13 55 17 56
rect 22 54 23 58
rect 27 54 28 58
rect 33 55 38 59
rect 13 50 17 51
rect 37 51 38 55
rect 43 58 49 64
rect 43 54 44 58
rect 48 54 49 58
rect 33 50 38 51
rect 2 46 38 50
rect 2 18 6 46
rect 42 43 46 51
rect 16 39 17 43
rect 21 39 22 43
rect 10 33 14 35
rect 18 34 22 39
rect 25 38 30 42
rect 34 38 46 43
rect 18 29 30 34
rect 34 29 38 38
rect 42 33 46 35
rect 10 25 14 29
rect 10 21 22 25
rect 2 14 9 18
rect 13 14 14 18
rect 2 13 6 14
rect 18 13 22 21
rect 26 13 30 29
rect 42 25 46 29
rect 34 21 46 25
rect 34 13 38 21
rect 42 14 43 18
rect 47 14 48 18
rect 42 8 48 14
rect -2 4 4 8
rect 8 4 47 8
rect 51 4 58 8
rect -2 0 58 4
<< ntransistor >>
rect 15 13 17 25
rect 22 13 24 25
rect 29 13 31 25
rect 36 13 38 25
<< ptransistor >>
rect 9 49 11 59
rect 19 49 21 59
rect 29 49 31 59
rect 39 49 41 59
<< polycontact >>
rect 17 39 21 43
rect 10 29 14 33
rect 30 38 34 42
rect 42 29 46 33
<< ndcontact >>
rect 9 14 13 18
rect 43 14 47 18
<< pdcontact >>
rect 3 54 7 58
rect 13 51 17 55
rect 23 54 27 58
rect 33 51 37 55
rect 44 54 48 58
<< psubstratepcontact >>
rect 4 4 8 8
rect 47 4 51 8
<< nsubstratencontact >>
rect 48 64 52 68
<< psubstratepdiff >>
rect 3 8 9 9
rect 45 8 53 9
rect 3 4 4 8
rect 8 4 9 8
rect 3 3 9 4
rect 45 4 47 8
rect 51 4 53 8
rect 45 3 53 4
<< nsubstratendiff >>
rect 47 68 53 69
rect 47 64 48 68
rect 52 64 53 68
rect 47 63 53 64
<< labels >>
rlabel metal1 4 28 4 28 6 z
rlabel metal1 12 28 12 28 6 d
rlabel metal1 12 48 12 48 6 z
rlabel metal1 28 4 28 4 6 vss
rlabel metal1 20 16 20 16 6 d
rlabel metal1 28 20 28 20 6 c
rlabel metal1 20 32 20 32 6 c
rlabel metal1 28 40 28 40 6 b
rlabel metal1 20 48 20 48 6 z
rlabel metal1 28 48 28 48 6 z
rlabel metal1 28 68 28 68 6 vdd
rlabel metal1 36 16 36 16 6 a
rlabel metal1 44 28 44 28 6 a
rlabel metal1 36 32 36 32 6 b
rlabel metal1 44 48 44 48 6 b
rlabel metal1 36 56 36 56 6 z
<< end >>
