magic
tech scmos
timestamp 1179386976
<< checkpaint >>
rect -22 -22 94 94
<< ab >>
rect 0 0 72 72
<< pwell >>
rect -4 -4 76 32
<< nwell >>
rect -4 32 76 76
<< polysilicon >>
rect 9 60 11 65
rect 21 56 23 61
rect 9 33 11 48
rect 44 54 46 59
rect 54 54 56 59
rect 61 54 63 59
rect 21 43 23 46
rect 15 42 23 43
rect 44 42 46 46
rect 15 38 16 42
rect 20 40 23 42
rect 40 40 46 42
rect 20 38 21 40
rect 15 37 21 38
rect 9 32 15 33
rect 9 28 10 32
rect 14 28 15 32
rect 9 27 15 28
rect 9 24 11 27
rect 19 25 21 37
rect 40 35 42 40
rect 54 35 56 38
rect 25 34 42 35
rect 25 30 26 34
rect 30 33 42 34
rect 30 30 31 33
rect 25 29 31 30
rect 40 26 42 33
rect 49 34 56 35
rect 49 30 50 34
rect 54 30 56 34
rect 49 29 56 30
rect 61 35 63 38
rect 61 34 67 35
rect 61 30 62 34
rect 66 30 67 34
rect 61 29 67 30
rect 50 26 52 29
rect 19 22 22 25
rect 20 19 22 22
rect 61 19 63 29
rect 9 13 11 18
rect 40 14 42 19
rect 50 14 52 19
rect 20 8 22 13
rect 61 7 63 12
<< ndiffusion >>
rect 33 25 40 26
rect 2 23 9 24
rect 2 19 3 23
rect 7 19 9 23
rect 2 18 9 19
rect 11 19 17 24
rect 33 21 34 25
rect 38 21 40 25
rect 33 19 40 21
rect 42 25 50 26
rect 42 21 44 25
rect 48 21 50 25
rect 42 19 50 21
rect 52 19 59 26
rect 11 18 20 19
rect 13 14 14 18
rect 18 14 20 18
rect 13 13 20 14
rect 22 18 29 19
rect 22 14 24 18
rect 28 14 29 18
rect 54 17 61 19
rect 22 13 29 14
rect 54 13 55 17
rect 59 13 61 17
rect 54 12 61 13
rect 63 18 70 19
rect 63 14 65 18
rect 69 14 70 18
rect 63 12 70 14
<< pdiffusion >>
rect 13 68 19 69
rect 13 64 14 68
rect 18 64 19 68
rect 13 60 19 64
rect 35 68 42 69
rect 35 64 37 68
rect 41 64 42 68
rect 2 59 9 60
rect 2 55 3 59
rect 7 55 9 59
rect 2 54 9 55
rect 4 48 9 54
rect 11 56 19 60
rect 11 48 21 56
rect 13 46 21 48
rect 23 52 28 56
rect 35 54 42 64
rect 23 51 31 52
rect 23 47 26 51
rect 30 47 31 51
rect 23 46 31 47
rect 35 46 44 54
rect 46 51 54 54
rect 46 47 48 51
rect 52 47 54 51
rect 46 46 54 47
rect 49 38 54 46
rect 56 38 61 54
rect 63 53 70 54
rect 63 49 65 53
rect 69 49 70 53
rect 63 38 70 49
<< metal1 >>
rect -2 68 74 72
rect -2 64 14 68
rect 18 64 26 68
rect 30 64 37 68
rect 41 64 56 68
rect 60 64 64 68
rect 68 64 74 68
rect 2 55 3 59
rect 7 55 62 59
rect 2 24 6 55
rect 26 51 30 52
rect 10 42 14 51
rect 10 38 16 42
rect 20 38 23 42
rect 26 34 30 47
rect 10 32 23 34
rect 14 30 23 32
rect 2 23 7 24
rect 2 19 3 23
rect 10 21 14 28
rect 26 26 30 30
rect 24 22 30 26
rect 34 47 48 51
rect 52 47 54 51
rect 34 45 54 47
rect 34 25 38 45
rect 58 42 62 55
rect 65 53 69 64
rect 65 48 69 49
rect 50 38 62 42
rect 50 34 54 38
rect 66 35 70 43
rect 50 29 54 30
rect 58 34 70 35
rect 58 30 62 34
rect 66 30 70 34
rect 58 29 70 30
rect 2 18 7 19
rect 24 18 28 22
rect 13 14 14 18
rect 18 14 19 18
rect 13 8 19 14
rect 24 13 28 14
rect 43 21 44 25
rect 48 21 69 25
rect 34 13 38 21
rect 65 18 69 21
rect 54 13 55 17
rect 59 13 60 17
rect 65 13 69 14
rect 54 8 60 13
rect -2 4 34 8
rect 38 4 42 8
rect 46 4 74 8
rect -2 0 74 4
<< ntransistor >>
rect 9 18 11 24
rect 40 19 42 26
rect 50 19 52 26
rect 20 13 22 19
rect 61 12 63 19
<< ptransistor >>
rect 9 48 11 60
rect 21 46 23 56
rect 44 46 46 54
rect 54 38 56 54
rect 61 38 63 54
<< polycontact >>
rect 16 38 20 42
rect 10 28 14 32
rect 26 30 30 34
rect 50 30 54 34
rect 62 30 66 34
<< ndcontact >>
rect 3 19 7 23
rect 34 21 38 25
rect 44 21 48 25
rect 14 14 18 18
rect 24 14 28 18
rect 55 13 59 17
rect 65 14 69 18
<< pdcontact >>
rect 14 64 18 68
rect 37 64 41 68
rect 3 55 7 59
rect 26 47 30 51
rect 48 47 52 51
rect 65 49 69 53
<< psubstratepcontact >>
rect 34 4 38 8
rect 42 4 46 8
<< nsubstratencontact >>
rect 26 64 30 68
rect 56 64 60 68
rect 64 64 68 68
<< psubstratepdiff >>
rect 33 8 47 9
rect 33 4 34 8
rect 38 4 42 8
rect 46 4 47 8
rect 33 3 47 4
<< nsubstratendiff >>
rect 25 68 31 69
rect 25 64 26 68
rect 30 64 31 68
rect 25 63 31 64
rect 55 68 69 69
rect 55 64 56 68
rect 60 64 64 68
rect 68 64 69 68
rect 55 63 69 64
<< labels >>
rlabel polycontact 28 32 28 32 6 bn
rlabel polycontact 52 32 52 32 6 a2n
rlabel metal1 12 24 12 24 6 a2
rlabel metal1 12 48 12 48 6 b
rlabel metal1 4 38 4 38 6 a2n
rlabel metal1 26 19 26 19 6 bn
rlabel metal1 20 32 20 32 6 a2
rlabel metal1 28 37 28 37 6 bn
rlabel metal1 20 40 20 40 6 b
rlabel metal1 36 4 36 4 6 vss
rlabel metal1 36 32 36 32 6 z
rlabel metal1 52 35 52 35 6 a2n
rlabel metal1 44 48 44 48 6 z
rlabel metal1 52 48 52 48 6 z
rlabel metal1 36 68 36 68 6 vdd
rlabel metal1 67 19 67 19 6 n1
rlabel metal1 56 23 56 23 6 n1
rlabel metal1 60 32 60 32 6 a1
rlabel metal1 68 36 68 36 6 a1
rlabel metal1 32 57 32 57 6 a2n
<< end >>
