magic
tech scmos
timestamp 1185038965
<< checkpaint >>
rect -22 -24 52 124
<< ab >>
rect 0 0 30 100
<< pwell >>
rect -2 -4 32 49
<< nwell >>
rect -2 49 32 104
<< polysilicon >>
rect 13 75 15 78
rect 13 43 15 55
rect 7 42 15 43
rect 7 38 8 42
rect 12 38 15 42
rect 7 37 15 38
rect 13 25 15 37
rect 13 12 15 15
<< ndiffusion >>
rect 3 15 13 25
rect 15 22 23 25
rect 15 18 18 22
rect 22 18 23 22
rect 15 15 23 18
rect 3 12 11 15
rect 3 8 6 12
rect 10 8 11 12
rect 3 7 11 8
<< pdiffusion >>
rect 3 92 11 93
rect 3 88 6 92
rect 10 88 11 92
rect 3 75 11 88
rect 3 55 13 75
rect 15 72 23 75
rect 15 68 18 72
rect 22 68 23 72
rect 15 62 23 68
rect 15 58 18 62
rect 22 58 23 62
rect 15 55 23 58
<< metal1 >>
rect -2 96 32 101
rect -2 92 18 96
rect 22 92 32 96
rect -2 88 6 92
rect 10 88 32 92
rect -2 87 32 88
rect 7 42 13 82
rect 7 38 8 42
rect 12 38 13 42
rect 7 18 13 38
rect 17 72 23 82
rect 17 68 18 72
rect 22 68 23 72
rect 17 62 23 68
rect 17 58 18 62
rect 22 58 23 62
rect 17 22 23 58
rect 17 18 18 22
rect 22 18 23 22
rect 17 17 23 18
rect -2 12 32 13
rect -2 8 6 12
rect 10 8 32 12
rect -2 -1 32 8
<< ntransistor >>
rect 13 15 15 25
<< ptransistor >>
rect 13 55 15 75
<< polycontact >>
rect 8 38 12 42
<< ndcontact >>
rect 18 18 22 22
rect 6 8 10 12
<< pdcontact >>
rect 6 88 10 92
rect 18 68 22 72
rect 18 58 22 62
<< nsubstratencontact >>
rect 18 92 22 96
<< nsubstratendiff >>
rect 17 96 23 97
rect 17 92 18 96
rect 22 92 23 96
rect 17 85 23 92
<< labels >>
rlabel metal1 15 6 15 6 6 vss
rlabel metal1 15 6 15 6 6 vss
rlabel metal1 10 50 10 50 6 i
rlabel metal1 10 50 10 50 6 i
rlabel metal1 15 94 15 94 6 vdd
rlabel metal1 15 94 15 94 6 vdd
rlabel metal1 20 50 20 50 6 nq
rlabel metal1 20 50 20 50 6 nq
<< end >>
