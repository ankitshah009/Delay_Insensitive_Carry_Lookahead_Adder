magic
tech scmos
timestamp 1179385295
<< checkpaint >>
rect -22 -22 78 94
<< ab >>
rect 0 0 56 72
<< pwell >>
rect -4 -4 60 32
<< nwell >>
rect -4 32 60 76
<< polysilicon >>
rect 9 66 11 70
rect 19 66 21 70
rect 29 66 31 70
rect 41 66 43 70
rect 9 29 11 39
rect 19 36 21 39
rect 19 35 25 36
rect 19 31 20 35
rect 24 31 25 35
rect 19 30 25 31
rect 29 35 31 39
rect 29 34 35 35
rect 29 30 30 34
rect 34 30 35 34
rect 9 28 15 29
rect 9 24 10 28
rect 14 24 15 28
rect 9 23 15 24
rect 12 19 14 23
rect 20 19 22 30
rect 29 29 35 30
rect 30 19 32 29
rect 41 28 43 39
rect 41 27 47 28
rect 41 24 42 27
rect 38 23 42 24
rect 46 23 47 27
rect 38 22 47 23
rect 38 19 40 22
rect 12 2 14 7
rect 20 2 22 7
rect 30 2 32 7
rect 38 2 40 7
<< ndiffusion >>
rect 3 8 12 19
rect 3 4 5 8
rect 9 7 12 8
rect 14 7 20 19
rect 22 17 30 19
rect 22 13 24 17
rect 28 13 30 17
rect 22 7 30 13
rect 32 7 38 19
rect 40 12 48 19
rect 40 8 42 12
rect 46 8 48 12
rect 40 7 48 8
rect 9 4 10 7
rect 3 3 10 4
<< pdiffusion >>
rect 4 59 9 66
rect 2 58 9 59
rect 2 54 3 58
rect 7 54 9 58
rect 2 53 9 54
rect 4 39 9 53
rect 11 51 19 66
rect 11 47 13 51
rect 17 47 19 51
rect 11 39 19 47
rect 21 58 29 66
rect 21 54 23 58
rect 27 54 29 58
rect 21 39 29 54
rect 31 65 41 66
rect 31 61 34 65
rect 38 61 41 65
rect 31 39 41 61
rect 43 59 48 66
rect 43 58 50 59
rect 43 54 45 58
rect 49 54 50 58
rect 43 53 50 54
rect 43 39 48 53
<< metal1 >>
rect -2 65 58 72
rect -2 64 34 65
rect 33 61 34 64
rect 38 64 58 65
rect 38 61 39 64
rect 2 54 3 58
rect 7 54 23 58
rect 27 54 45 58
rect 49 54 50 58
rect 2 47 13 51
rect 17 47 18 51
rect 2 19 6 47
rect 26 43 30 51
rect 10 28 14 43
rect 18 37 30 43
rect 34 46 47 50
rect 20 35 24 37
rect 20 30 24 31
rect 29 30 30 34
rect 34 29 38 46
rect 42 27 46 35
rect 14 24 22 27
rect 10 23 22 24
rect 18 21 22 23
rect 26 25 30 27
rect 26 23 42 25
rect 26 21 46 23
rect 2 17 14 19
rect 2 13 24 17
rect 28 13 29 17
rect 34 13 38 21
rect 42 12 46 13
rect -2 4 5 8
rect 9 4 58 8
rect -2 0 58 4
<< ntransistor >>
rect 12 7 14 19
rect 20 7 22 19
rect 30 7 32 19
rect 38 7 40 19
<< ptransistor >>
rect 9 39 11 66
rect 19 39 21 66
rect 29 39 31 66
rect 41 39 43 66
<< polycontact >>
rect 20 31 24 35
rect 30 30 34 34
rect 10 24 14 28
rect 42 23 46 27
<< ndcontact >>
rect 5 4 9 8
rect 24 13 28 17
rect 42 8 46 12
<< pdcontact >>
rect 3 54 7 58
rect 13 47 17 51
rect 23 54 27 58
rect 34 61 38 65
rect 45 54 49 58
<< labels >>
rlabel metal1 4 32 4 32 6 z
rlabel metal1 12 16 12 16 6 z
rlabel metal1 20 24 20 24 6 b1
rlabel metal1 20 40 20 40 6 b2
rlabel metal1 12 36 12 36 6 b1
rlabel metal1 28 4 28 4 6 vss
rlabel metal1 36 16 36 16 6 a1
rlabel metal1 28 24 28 24 6 a1
rlabel metal1 36 36 36 36 6 a2
rlabel metal1 28 44 28 44 6 b2
rlabel metal1 28 68 28 68 6 vdd
rlabel metal1 44 28 44 28 6 a1
rlabel metal1 44 48 44 48 6 a2
rlabel pdcontact 26 56 26 56 6 n3
<< end >>
