magic
tech scmos
timestamp 1185038988
<< checkpaint >>
rect -22 -24 62 124
<< ab >>
rect 0 0 40 100
<< pwell >>
rect -2 -4 42 49
<< nwell >>
rect -2 49 42 104
<< polysilicon >>
rect 13 85 15 88
rect 25 85 27 88
rect 13 63 15 65
rect 7 62 15 63
rect 7 58 8 62
rect 12 58 15 62
rect 7 57 15 58
rect 13 35 15 57
rect 25 43 27 65
rect 25 42 33 43
rect 25 39 28 42
rect 21 38 28 39
rect 32 38 33 42
rect 21 37 33 38
rect 21 35 23 37
rect 13 12 15 15
rect 21 12 23 15
<< ndiffusion >>
rect 5 15 13 35
rect 15 15 21 35
rect 23 22 31 35
rect 23 18 26 22
rect 30 18 31 22
rect 23 15 31 18
rect 5 12 11 15
rect 5 8 6 12
rect 10 8 11 12
rect 5 7 11 8
<< pdiffusion >>
rect 5 92 11 93
rect 5 88 6 92
rect 10 88 11 92
rect 29 92 35 93
rect 29 88 30 92
rect 34 88 35 92
rect 5 85 11 88
rect 29 85 35 88
rect 5 65 13 85
rect 15 82 25 85
rect 15 78 18 82
rect 22 78 25 82
rect 15 72 25 78
rect 15 68 18 72
rect 22 68 25 72
rect 15 65 25 68
rect 27 65 35 85
<< metal1 >>
rect -2 92 42 101
rect -2 88 6 92
rect 10 88 30 92
rect 34 88 42 92
rect -2 87 42 88
rect 17 82 23 83
rect 7 62 13 82
rect 7 58 8 62
rect 12 58 13 62
rect 7 18 13 58
rect 17 78 18 82
rect 22 78 23 82
rect 17 72 23 78
rect 17 68 18 72
rect 22 68 23 72
rect 17 23 23 68
rect 27 42 33 82
rect 27 38 28 42
rect 32 38 33 42
rect 27 28 33 38
rect 17 22 31 23
rect 17 18 26 22
rect 30 18 31 22
rect 17 17 31 18
rect -2 12 42 13
rect -2 8 6 12
rect 10 8 42 12
rect -2 4 23 8
rect 27 4 42 8
rect -2 -1 42 4
<< ntransistor >>
rect 13 15 15 35
rect 21 15 23 35
<< ptransistor >>
rect 13 65 15 85
rect 25 65 27 85
<< polycontact >>
rect 8 58 12 62
rect 28 38 32 42
<< ndcontact >>
rect 26 18 30 22
rect 6 8 10 12
<< pdcontact >>
rect 6 88 10 92
rect 30 88 34 92
rect 18 78 22 82
rect 18 68 22 72
<< psubstratepcontact >>
rect 23 4 27 8
<< psubstratepdiff >>
rect 22 8 35 9
rect 22 4 23 8
rect 27 4 35 8
rect 22 3 35 4
<< labels >>
rlabel metal1 10 50 10 50 6 i0
rlabel metal1 10 50 10 50 6 i0
rlabel metal1 20 6 20 6 6 vss
rlabel metal1 20 6 20 6 6 vss
rlabel metal1 20 50 20 50 6 nq
rlabel metal1 20 50 20 50 6 nq
rlabel metal1 30 55 30 55 6 i1
rlabel metal1 30 55 30 55 6 i1
rlabel metal1 20 94 20 94 6 vdd
rlabel metal1 20 94 20 94 6 vdd
<< end >>
