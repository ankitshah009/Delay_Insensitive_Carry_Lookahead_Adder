magic
tech scmos
timestamp 1179387308
<< checkpaint >>
rect -22 -25 86 105
<< ab >>
rect 0 0 64 80
<< pwell >>
rect -4 -7 68 36
<< nwell >>
rect -4 36 68 87
<< polysilicon >>
rect 9 70 11 74
rect 28 70 30 74
rect 35 70 37 74
rect 42 70 44 74
rect 49 70 51 74
rect 9 39 11 42
rect 28 39 30 42
rect 9 38 15 39
rect 9 34 10 38
rect 14 34 15 38
rect 9 33 15 34
rect 19 38 30 39
rect 19 34 20 38
rect 24 37 30 38
rect 24 34 25 37
rect 19 33 25 34
rect 9 24 11 33
rect 20 22 22 33
rect 35 31 37 42
rect 30 30 37 31
rect 30 26 32 30
rect 36 26 37 30
rect 30 25 37 26
rect 42 31 44 42
rect 49 39 51 42
rect 49 38 59 39
rect 49 37 54 38
rect 52 34 54 37
rect 58 34 59 38
rect 52 33 59 34
rect 42 30 48 31
rect 42 26 43 30
rect 47 26 48 30
rect 42 25 48 26
rect 30 22 32 25
rect 42 22 44 25
rect 52 22 54 33
rect 9 6 11 10
rect 20 9 22 14
rect 30 9 32 14
rect 42 9 44 14
rect 52 9 54 14
<< ndiffusion >>
rect 2 23 9 24
rect 2 19 3 23
rect 7 19 9 23
rect 2 18 9 19
rect 4 10 9 18
rect 11 22 18 24
rect 11 18 13 22
rect 17 18 20 22
rect 11 15 20 18
rect 11 11 13 15
rect 17 14 20 15
rect 22 21 30 22
rect 22 17 24 21
rect 28 17 30 21
rect 22 14 30 17
rect 32 14 42 22
rect 44 21 52 22
rect 44 17 46 21
rect 50 17 52 21
rect 44 14 52 17
rect 54 14 62 22
rect 17 11 18 14
rect 11 10 18 11
rect 34 12 40 14
rect 34 8 35 12
rect 39 8 40 12
rect 56 12 62 14
rect 34 7 40 8
rect 56 8 57 12
rect 61 8 62 12
rect 56 7 62 8
<< pdiffusion >>
rect 13 70 19 72
rect 4 56 9 70
rect 2 55 9 56
rect 2 51 3 55
rect 7 51 9 55
rect 2 50 9 51
rect 4 42 9 50
rect 11 66 14 70
rect 18 66 19 70
rect 11 59 19 66
rect 11 42 17 59
rect 23 55 28 70
rect 21 54 28 55
rect 21 50 22 54
rect 26 50 28 54
rect 21 49 28 50
rect 23 42 28 49
rect 30 42 35 70
rect 37 42 42 70
rect 44 42 49 70
rect 51 69 59 70
rect 51 65 53 69
rect 57 65 59 69
rect 51 62 59 65
rect 51 58 53 62
rect 57 58 59 62
rect 51 42 59 58
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect -2 70 66 78
rect -2 68 14 70
rect 13 66 14 68
rect 18 69 66 70
rect 18 68 53 69
rect 18 66 19 68
rect 52 65 53 68
rect 57 68 66 69
rect 57 65 58 68
rect 2 57 14 63
rect 2 55 7 57
rect 2 51 3 55
rect 2 50 7 51
rect 11 50 22 54
rect 26 50 27 54
rect 2 24 6 50
rect 11 39 15 50
rect 34 46 38 63
rect 52 62 58 65
rect 52 58 53 62
rect 57 58 58 62
rect 10 38 15 39
rect 14 34 15 38
rect 19 42 38 46
rect 42 46 46 55
rect 42 42 59 46
rect 19 38 25 42
rect 53 38 59 42
rect 19 34 20 38
rect 24 34 25 38
rect 32 34 47 38
rect 53 34 54 38
rect 58 34 59 38
rect 10 33 15 34
rect 11 30 15 33
rect 32 30 38 34
rect 11 26 27 30
rect 2 23 7 24
rect 2 19 3 23
rect 2 17 7 19
rect 12 18 13 22
rect 17 18 18 22
rect 12 15 18 18
rect 23 21 27 26
rect 36 26 38 30
rect 42 26 43 30
rect 47 26 62 30
rect 32 25 38 26
rect 23 17 24 21
rect 28 17 46 21
rect 50 17 51 21
rect 58 17 62 26
rect 12 12 13 15
rect -2 11 13 12
rect 17 12 18 15
rect 17 11 35 12
rect -2 8 35 11
rect 39 8 57 12
rect 61 8 66 12
rect -2 2 66 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
<< ntransistor >>
rect 9 10 11 24
rect 20 14 22 22
rect 30 14 32 22
rect 42 14 44 22
rect 52 14 54 22
<< ptransistor >>
rect 9 42 11 70
rect 28 42 30 70
rect 35 42 37 70
rect 42 42 44 70
rect 49 42 51 70
<< polycontact >>
rect 10 34 14 38
rect 20 34 24 38
rect 32 26 36 30
rect 54 34 58 38
rect 43 26 47 30
<< ndcontact >>
rect 3 19 7 23
rect 13 18 17 22
rect 13 11 17 15
rect 24 17 28 21
rect 46 17 50 21
rect 35 8 39 12
rect 57 8 61 12
<< pdcontact >>
rect 3 51 7 55
rect 14 66 18 70
rect 22 50 26 54
rect 53 65 57 69
rect 53 58 57 62
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
<< psubstratepdiff >>
rect 0 2 64 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 64 2
rect 0 -3 64 -2
<< nsubstratendiff >>
rect 0 82 64 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 64 82
rect 0 77 64 78
<< labels >>
rlabel polycontact 12 36 12 36 6 zn
rlabel metal1 4 40 4 40 6 z
rlabel metal1 13 40 13 40 6 zn
rlabel metal1 12 60 12 60 6 z
rlabel metal1 32 6 32 6 6 vss
rlabel metal1 36 32 36 32 6 c
rlabel metal1 28 44 28 44 6 d
rlabel metal1 19 52 19 52 6 zn
rlabel metal1 36 56 36 56 6 d
rlabel metal1 32 74 32 74 6 vdd
rlabel metal1 37 19 37 19 6 zn
rlabel metal1 44 36 44 36 6 c
rlabel metal1 44 52 44 52 6 a
rlabel metal1 52 28 52 28 6 b
rlabel metal1 60 20 60 20 6 b
rlabel metal1 52 44 52 44 6 a
<< end >>
