magic
tech scmos
timestamp 1180600619
<< checkpaint >>
rect -22 -22 72 122
<< ab >>
rect 0 0 50 100
<< pwell >>
rect -4 -4 54 48
<< nwell >>
rect -4 48 54 104
<< polysilicon >>
rect 17 94 19 98
rect 25 94 27 98
rect 37 76 39 80
rect 17 43 19 55
rect 13 42 21 43
rect 13 38 16 42
rect 20 38 21 42
rect 13 37 21 38
rect 25 41 27 55
rect 37 53 39 56
rect 31 52 39 53
rect 31 48 32 52
rect 36 48 39 52
rect 31 47 39 48
rect 41 42 47 43
rect 41 41 42 42
rect 25 39 42 41
rect 13 25 15 37
rect 25 25 27 39
rect 41 38 42 39
rect 46 38 47 42
rect 41 37 47 38
rect 31 32 39 33
rect 31 28 32 32
rect 36 28 39 32
rect 31 27 39 28
rect 37 24 39 27
rect 13 11 15 15
rect 25 11 27 15
rect 37 10 39 14
<< ndiffusion >>
rect 5 15 13 25
rect 15 22 25 25
rect 15 18 18 22
rect 22 18 25 22
rect 15 15 25 18
rect 27 24 32 25
rect 27 15 37 24
rect 5 12 11 15
rect 5 8 6 12
rect 10 8 11 12
rect 29 14 37 15
rect 39 22 47 24
rect 39 18 42 22
rect 46 18 47 22
rect 39 14 47 18
rect 29 12 35 14
rect 5 7 11 8
rect 29 8 30 12
rect 34 8 35 12
rect 29 7 35 8
<< pdiffusion >>
rect 12 85 17 94
rect 5 82 17 85
rect 5 78 6 82
rect 10 78 17 82
rect 5 72 17 78
rect 5 68 6 72
rect 10 68 17 72
rect 5 62 17 68
rect 5 58 6 62
rect 10 58 17 62
rect 5 55 17 58
rect 19 55 25 94
rect 27 92 35 94
rect 27 88 30 92
rect 34 88 35 92
rect 27 76 35 88
rect 27 56 37 76
rect 39 72 47 76
rect 39 68 42 72
rect 46 68 47 72
rect 39 62 47 68
rect 39 58 42 62
rect 46 58 47 62
rect 39 56 47 58
rect 27 55 32 56
<< metal1 >>
rect -2 96 52 100
rect -2 92 42 96
rect 46 92 52 96
rect -2 88 30 92
rect 34 88 52 92
rect 8 82 12 83
rect 5 78 6 82
rect 10 78 12 82
rect 8 72 12 78
rect 5 68 6 72
rect 10 68 12 72
rect 8 62 12 68
rect 5 58 6 62
rect 10 58 12 62
rect 8 52 12 58
rect 4 47 12 52
rect 4 33 8 47
rect 18 42 22 83
rect 15 38 16 42
rect 20 38 22 42
rect 4 28 12 33
rect 8 22 12 28
rect 18 27 22 38
rect 8 18 18 22
rect 22 18 23 22
rect 8 17 12 18
rect 28 17 32 83
rect 42 72 46 73
rect 42 62 46 68
rect 36 48 37 52
rect 42 42 46 58
rect 36 28 37 32
rect 42 22 46 38
rect 42 17 46 18
rect -2 8 6 12
rect 10 8 30 12
rect 34 8 52 12
rect -2 0 52 8
<< ntransistor >>
rect 13 15 15 25
rect 25 15 27 25
rect 37 14 39 24
<< ptransistor >>
rect 17 55 19 94
rect 25 55 27 94
rect 37 56 39 76
<< polycontact >>
rect 16 38 20 42
rect 32 48 36 52
rect 42 38 46 42
rect 32 28 36 32
<< ndcontact >>
rect 18 18 22 22
rect 6 8 10 12
rect 42 18 46 22
rect 30 8 34 12
<< pdcontact >>
rect 6 78 10 82
rect 6 68 10 72
rect 6 58 10 62
rect 30 88 34 92
rect 42 68 46 72
rect 42 58 46 62
<< nsubstratencontact >>
rect 42 92 46 96
<< nsubstratendiff >>
rect 41 96 47 97
rect 41 92 42 96
rect 46 92 47 96
rect 41 86 47 92
<< labels >>
rlabel ndcontact 20 20 20 20 6 q
rlabel metal1 10 25 10 25 6 q
rlabel metal1 10 65 10 65 6 q
rlabel metal1 20 55 20 55 6 i0
rlabel metal1 25 6 25 6 6 vss
rlabel metal1 30 50 30 50 6 i1
rlabel metal1 25 94 25 94 6 vdd
<< end >>
