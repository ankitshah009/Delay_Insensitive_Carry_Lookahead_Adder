magic
tech scmos
timestamp 1180640008
<< checkpaint >>
rect -24 -26 94 126
<< ab >>
rect 0 0 70 100
<< pwell >>
rect -4 -6 74 49
<< nwell >>
rect -4 49 74 106
<< polysilicon >>
rect 13 94 15 98
rect 25 94 27 98
rect 33 94 35 98
rect 45 94 47 98
rect 57 94 59 98
rect 13 52 15 55
rect 25 52 27 55
rect 13 51 27 52
rect 13 47 18 51
rect 22 47 27 51
rect 13 46 27 47
rect 13 35 15 46
rect 25 35 27 46
rect 33 52 35 55
rect 45 52 47 55
rect 57 52 59 55
rect 33 51 41 52
rect 33 47 36 51
rect 40 47 41 51
rect 33 46 41 47
rect 45 51 53 52
rect 45 47 48 51
rect 52 47 53 51
rect 45 46 53 47
rect 57 51 63 52
rect 57 47 58 51
rect 62 47 63 51
rect 57 46 63 47
rect 33 35 35 46
rect 45 35 47 46
rect 57 35 59 46
rect 13 12 15 17
rect 25 12 27 17
rect 33 12 35 17
rect 45 12 47 17
rect 57 12 59 17
<< ndiffusion >>
rect 8 31 13 35
rect 5 30 13 31
rect 5 26 6 30
rect 10 26 13 30
rect 5 22 13 26
rect 5 18 6 22
rect 10 18 13 22
rect 5 17 13 18
rect 15 17 25 35
rect 27 17 33 35
rect 35 32 45 35
rect 35 28 38 32
rect 42 28 45 32
rect 35 17 45 28
rect 47 32 57 35
rect 47 28 50 32
rect 54 28 57 32
rect 47 22 57 28
rect 47 18 50 22
rect 54 18 57 22
rect 47 17 57 18
rect 59 32 67 35
rect 59 28 62 32
rect 66 28 67 32
rect 59 22 67 28
rect 59 18 62 22
rect 66 18 67 22
rect 59 17 67 18
rect 17 12 23 17
rect 17 8 18 12
rect 22 8 23 12
rect 17 7 23 8
<< pdiffusion >>
rect 8 83 13 94
rect 5 82 13 83
rect 5 78 6 82
rect 10 78 13 82
rect 5 74 13 78
rect 5 70 6 74
rect 10 70 13 74
rect 5 69 13 70
rect 8 55 13 69
rect 15 92 25 94
rect 15 88 18 92
rect 22 88 25 92
rect 15 82 25 88
rect 15 78 18 82
rect 22 78 25 82
rect 15 55 25 78
rect 27 55 33 94
rect 35 72 45 94
rect 35 68 38 72
rect 42 68 45 72
rect 35 62 45 68
rect 35 58 38 62
rect 42 58 45 62
rect 35 55 45 58
rect 47 82 57 94
rect 47 78 50 82
rect 54 78 57 82
rect 47 55 57 78
rect 59 92 67 94
rect 59 88 62 92
rect 66 88 67 92
rect 59 82 67 88
rect 59 78 62 82
rect 66 78 67 82
rect 59 55 67 78
<< metal1 >>
rect -2 92 72 100
rect -2 88 18 92
rect 22 88 62 92
rect 66 88 72 92
rect 6 82 10 83
rect 6 74 10 78
rect 18 82 22 88
rect 62 82 66 88
rect 18 77 22 78
rect 28 78 50 82
rect 54 78 55 82
rect 28 72 32 78
rect 62 77 66 78
rect 10 70 32 72
rect 6 68 32 70
rect 38 72 42 73
rect 38 63 42 68
rect 8 52 12 63
rect 28 62 42 63
rect 28 58 38 62
rect 28 57 42 58
rect 47 68 63 72
rect 8 51 23 52
rect 8 47 18 51
rect 22 47 23 51
rect 8 46 23 47
rect 8 37 12 46
rect 28 32 32 57
rect 36 51 42 53
rect 40 47 42 51
rect 47 51 53 68
rect 47 47 48 51
rect 52 47 53 51
rect 58 51 62 63
rect 36 42 42 47
rect 58 42 62 47
rect 36 37 62 42
rect 50 32 55 33
rect 5 26 6 30
rect 10 26 11 30
rect 28 28 38 32
rect 42 28 43 32
rect 28 27 43 28
rect 54 28 55 32
rect 5 22 11 26
rect 50 22 55 28
rect 5 18 6 22
rect 10 18 50 22
rect 54 18 55 22
rect 62 32 66 33
rect 62 22 66 28
rect 62 12 66 18
rect -2 8 18 12
rect 22 8 72 12
rect -2 0 72 8
<< ntransistor >>
rect 13 17 15 35
rect 25 17 27 35
rect 33 17 35 35
rect 45 17 47 35
rect 57 17 59 35
<< ptransistor >>
rect 13 55 15 94
rect 25 55 27 94
rect 33 55 35 94
rect 45 55 47 94
rect 57 55 59 94
<< polycontact >>
rect 18 47 22 51
rect 36 47 40 51
rect 48 47 52 51
rect 58 47 62 51
<< ndcontact >>
rect 6 26 10 30
rect 6 18 10 22
rect 38 28 42 32
rect 50 28 54 32
rect 50 18 54 22
rect 62 28 66 32
rect 62 18 66 22
rect 18 8 22 12
<< pdcontact >>
rect 6 78 10 82
rect 6 70 10 74
rect 18 88 22 92
rect 18 78 22 82
rect 38 68 42 72
rect 38 58 42 62
rect 50 78 54 82
rect 62 88 66 92
rect 62 78 66 82
<< psubstratepcontact >>
rect 48 4 52 8
rect 58 4 62 8
<< psubstratepdiff >>
rect 47 8 63 9
rect 47 4 48 8
rect 52 4 58 8
rect 62 4 63 8
rect 47 3 63 4
<< labels >>
rlabel metal1 8 24 8 24 6 n4
rlabel metal1 8 75 8 75 6 n2
rlabel metal1 10 50 10 50 6 a
rlabel metal1 10 50 10 50 6 a
rlabel polycontact 20 50 20 50 6 a
rlabel polycontact 20 50 20 50 6 a
rlabel metal1 35 6 35 6 6 vss
rlabel metal1 35 6 35 6 6 vss
rlabel metal1 30 45 30 45 6 z
rlabel metal1 30 45 30 45 6 z
rlabel metal1 35 94 35 94 6 vdd
rlabel metal1 35 94 35 94 6 vdd
rlabel metal1 52 25 52 25 6 n4
rlabel metal1 30 20 30 20 6 n4
rlabel ndcontact 40 30 40 30 6 z
rlabel ndcontact 40 30 40 30 6 z
rlabel metal1 50 40 50 40 6 b
rlabel metal1 50 40 50 40 6 b
rlabel metal1 40 45 40 45 6 b
rlabel metal1 40 45 40 45 6 b
rlabel metal1 50 60 50 60 6 c
rlabel metal1 50 60 50 60 6 c
rlabel metal1 40 65 40 65 6 z
rlabel metal1 40 65 40 65 6 z
rlabel metal1 41 80 41 80 6 n2
rlabel polycontact 60 50 60 50 6 b
rlabel polycontact 60 50 60 50 6 b
rlabel metal1 60 70 60 70 6 c
rlabel metal1 60 70 60 70 6 c
<< end >>
