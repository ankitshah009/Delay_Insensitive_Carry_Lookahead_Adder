magic
tech scmos
timestamp 1179385349
<< checkpaint >>
rect -22 -25 78 105
<< ab >>
rect 0 0 56 80
<< pwell >>
rect -4 -7 60 36
<< nwell >>
rect -4 36 60 87
<< polysilicon >>
rect 31 66 33 71
rect 41 66 43 71
rect 9 61 11 65
rect 19 61 21 65
rect 31 47 33 50
rect 30 46 37 47
rect 9 39 11 45
rect 19 42 21 45
rect 30 42 32 46
rect 36 42 37 46
rect 19 41 26 42
rect 9 38 15 39
rect 9 34 10 38
rect 14 34 15 38
rect 19 37 21 41
rect 25 37 26 41
rect 19 36 26 37
rect 30 41 37 42
rect 9 33 15 34
rect 13 24 15 33
rect 23 28 25 36
rect 30 28 32 41
rect 41 37 43 50
rect 41 36 47 37
rect 41 33 42 36
rect 37 32 42 33
rect 46 32 47 36
rect 37 31 47 32
rect 37 28 39 31
rect 13 13 15 18
rect 23 13 25 18
rect 30 13 32 18
rect 37 13 39 18
<< ndiffusion >>
rect 18 24 23 28
rect 3 18 13 24
rect 15 23 23 24
rect 15 19 17 23
rect 21 19 23 23
rect 15 18 23 19
rect 25 18 30 28
rect 32 18 37 28
rect 39 23 50 28
rect 39 19 44 23
rect 48 19 50 23
rect 39 18 50 19
rect 3 12 10 18
rect 3 8 5 12
rect 9 8 10 12
rect 3 7 10 8
<< pdiffusion >>
rect 23 72 29 73
rect 23 68 24 72
rect 28 68 29 72
rect 23 66 29 68
rect 23 61 31 66
rect 4 58 9 61
rect 2 57 9 58
rect 2 53 3 57
rect 7 53 9 57
rect 2 50 9 53
rect 2 46 3 50
rect 7 46 9 50
rect 2 45 9 46
rect 11 60 19 61
rect 11 56 13 60
rect 17 56 19 60
rect 11 45 19 56
rect 21 50 31 61
rect 33 62 41 66
rect 33 58 35 62
rect 39 58 41 62
rect 33 55 41 58
rect 33 51 35 55
rect 39 51 41 55
rect 33 50 41 51
rect 43 65 50 66
rect 43 61 45 65
rect 49 61 50 65
rect 43 50 50 61
rect 21 45 26 50
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect -2 72 58 78
rect -2 68 24 72
rect 28 68 58 72
rect 45 65 49 68
rect 2 57 7 63
rect 2 53 3 57
rect 13 62 39 63
rect 13 60 35 62
rect 17 59 35 60
rect 13 55 17 56
rect 45 60 49 61
rect 35 55 39 58
rect 2 50 7 53
rect 2 46 3 50
rect 21 50 31 54
rect 35 50 39 51
rect 21 47 25 50
rect 2 45 7 46
rect 2 23 6 45
rect 18 41 25 47
rect 42 46 47 55
rect 31 42 32 46
rect 36 42 47 46
rect 10 38 14 39
rect 25 37 31 38
rect 21 34 31 37
rect 41 36 47 38
rect 10 30 14 34
rect 41 32 42 36
rect 46 32 47 36
rect 41 30 47 32
rect 10 26 31 30
rect 35 26 47 30
rect 2 19 17 23
rect 21 19 22 23
rect 35 22 39 26
rect 2 17 15 19
rect 25 18 39 22
rect 43 19 44 23
rect 48 19 49 23
rect 43 12 49 19
rect -2 8 5 12
rect 9 8 58 12
rect -2 2 58 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
<< ntransistor >>
rect 13 18 15 24
rect 23 18 25 28
rect 30 18 32 28
rect 37 18 39 28
<< ptransistor >>
rect 9 45 11 61
rect 19 45 21 61
rect 31 50 33 66
rect 41 50 43 66
<< polycontact >>
rect 32 42 36 46
rect 10 34 14 38
rect 21 37 25 41
rect 42 32 46 36
<< ndcontact >>
rect 17 19 21 23
rect 44 19 48 23
rect 5 8 9 12
<< pdcontact >>
rect 24 68 28 72
rect 3 53 7 57
rect 3 46 7 50
rect 13 56 17 60
rect 35 58 39 62
rect 35 51 39 55
rect 45 61 49 65
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
<< psubstratepdiff >>
rect 0 2 56 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 56 2
rect 0 -3 56 -2
<< nsubstratendiff >>
rect 0 82 56 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 56 82
rect 0 77 56 78
<< labels >>
rlabel metal1 4 40 4 40 6 z
rlabel metal1 12 20 12 20 6 z
rlabel polycontact 12 36 12 36 6 b
rlabel metal1 28 6 28 6 6 vss
rlabel metal1 20 28 20 28 6 b
rlabel metal1 28 20 28 20 6 a1
rlabel metal1 28 28 28 28 6 b
rlabel metal1 20 44 20 44 6 a3
rlabel metal1 28 36 28 36 6 a3
rlabel metal1 28 52 28 52 6 a3
rlabel metal1 28 74 28 74 6 vdd
rlabel metal1 36 20 36 20 6 a1
rlabel metal1 44 32 44 32 6 a1
rlabel metal1 36 44 36 44 6 a2
rlabel metal1 44 48 44 48 6 a2
rlabel metal1 37 56 37 56 6 n3
rlabel metal1 26 61 26 61 6 n3
<< end >>
