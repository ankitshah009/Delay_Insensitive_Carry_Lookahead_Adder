magic
tech scmos
timestamp 1185039016
<< checkpaint >>
rect -22 -24 92 124
<< ab >>
rect 0 0 70 100
<< pwell >>
rect -2 -4 72 49
<< nwell >>
rect -2 49 72 104
<< polysilicon >>
rect 23 95 25 98
rect 33 95 35 98
rect 45 95 47 98
rect 57 95 59 98
rect 11 85 13 88
rect 11 41 13 65
rect 23 53 25 55
rect 17 52 25 53
rect 17 48 18 52
rect 22 51 25 52
rect 22 48 23 51
rect 17 47 23 48
rect 33 43 35 55
rect 45 53 47 55
rect 57 53 59 55
rect 45 52 53 53
rect 45 51 48 52
rect 47 48 48 51
rect 52 48 53 52
rect 47 47 53 48
rect 57 52 63 53
rect 57 48 58 52
rect 62 48 63 52
rect 57 47 63 48
rect 27 42 35 43
rect 27 41 28 42
rect 11 39 28 41
rect 11 25 13 39
rect 27 38 28 39
rect 32 41 35 42
rect 32 39 47 41
rect 32 38 33 39
rect 27 37 33 38
rect 17 32 23 33
rect 17 28 18 32
rect 22 29 23 32
rect 29 32 35 33
rect 22 28 25 29
rect 17 27 25 28
rect 29 28 30 32
rect 34 28 35 32
rect 29 27 35 28
rect 23 25 25 27
rect 33 25 35 27
rect 45 25 47 39
rect 57 32 63 33
rect 57 28 58 32
rect 62 28 63 32
rect 57 27 63 28
rect 57 25 59 27
rect 11 12 13 15
rect 23 2 25 5
rect 33 2 35 5
rect 45 2 47 5
rect 57 2 59 5
<< ndiffusion >>
rect 3 22 11 25
rect 3 18 4 22
rect 8 18 11 22
rect 3 15 11 18
rect 13 15 23 25
rect 15 12 23 15
rect 15 8 16 12
rect 20 8 23 12
rect 15 5 23 8
rect 25 5 33 25
rect 35 22 45 25
rect 35 18 38 22
rect 42 18 45 22
rect 35 5 45 18
rect 47 5 57 25
rect 59 12 67 25
rect 59 8 62 12
rect 66 8 67 12
rect 59 5 67 8
<< pdiffusion >>
rect 15 92 23 95
rect 15 88 16 92
rect 20 88 23 92
rect 15 85 23 88
rect 3 82 11 85
rect 3 78 4 82
rect 8 78 11 82
rect 3 72 11 78
rect 3 68 4 72
rect 8 68 11 72
rect 3 65 11 68
rect 13 65 23 85
rect 15 55 23 65
rect 25 55 33 95
rect 35 72 45 95
rect 35 68 38 72
rect 42 68 45 72
rect 35 62 45 68
rect 35 58 38 62
rect 42 58 45 62
rect 35 55 45 58
rect 47 55 57 95
rect 59 92 67 95
rect 59 88 62 92
rect 66 88 67 92
rect 59 55 67 88
<< metal1 >>
rect -2 92 72 101
rect -2 88 16 92
rect 20 88 62 92
rect 66 88 72 92
rect -2 87 72 88
rect 3 82 9 83
rect 3 78 4 82
rect 8 78 52 82
rect 3 77 9 78
rect 4 73 8 77
rect 3 72 9 73
rect 37 72 43 73
rect 3 68 4 72
rect 8 68 9 72
rect 3 67 9 68
rect 4 23 8 67
rect 17 52 23 72
rect 17 48 18 52
rect 22 48 23 52
rect 17 32 23 48
rect 27 42 33 72
rect 27 38 28 42
rect 32 38 33 42
rect 27 37 33 38
rect 37 68 38 72
rect 42 68 43 72
rect 37 62 43 68
rect 37 58 38 62
rect 42 58 43 62
rect 37 43 43 58
rect 48 53 52 78
rect 47 52 53 53
rect 47 48 48 52
rect 52 48 53 52
rect 47 47 53 48
rect 57 52 63 82
rect 57 48 58 52
rect 62 48 63 52
rect 37 37 45 43
rect 39 33 45 37
rect 17 28 18 32
rect 22 28 23 32
rect 17 27 23 28
rect 29 32 35 33
rect 29 28 30 32
rect 34 28 35 32
rect 29 27 35 28
rect 39 27 52 33
rect 57 32 63 48
rect 57 28 58 32
rect 62 28 63 32
rect 3 22 9 23
rect 29 22 33 27
rect 39 23 45 27
rect 3 18 4 22
rect 8 18 33 22
rect 37 22 45 23
rect 37 18 38 22
rect 42 18 45 22
rect 57 18 63 28
rect 3 17 9 18
rect 37 17 45 18
rect -2 12 72 13
rect -2 8 16 12
rect 20 8 62 12
rect 66 8 72 12
rect -2 -1 72 8
<< ntransistor >>
rect 11 15 13 25
rect 23 5 25 25
rect 33 5 35 25
rect 45 5 47 25
rect 57 5 59 25
<< ptransistor >>
rect 11 65 13 85
rect 23 55 25 95
rect 33 55 35 95
rect 45 55 47 95
rect 57 55 59 95
<< polycontact >>
rect 18 48 22 52
rect 48 48 52 52
rect 58 48 62 52
rect 28 38 32 42
rect 18 28 22 32
rect 30 28 34 32
rect 58 28 62 32
<< ndcontact >>
rect 4 18 8 22
rect 16 8 20 12
rect 38 18 42 22
rect 62 8 66 12
<< pdcontact >>
rect 16 88 20 92
rect 4 78 8 82
rect 4 68 8 72
rect 38 68 42 72
rect 38 58 42 62
rect 62 88 66 92
<< labels >>
rlabel polycontact 20 50 20 50 6 i0
rlabel polycontact 20 50 20 50 6 i0
rlabel metal1 30 55 30 55 6 cmd
rlabel metal1 30 55 30 55 6 cmd
rlabel metal1 35 6 35 6 6 vss
rlabel metal1 35 6 35 6 6 vss
rlabel ndcontact 40 20 40 20 6 nq
rlabel ndcontact 40 20 40 20 6 nq
rlabel metal1 50 30 50 30 6 nq
rlabel metal1 50 30 50 30 6 nq
rlabel metal1 40 55 40 55 6 nq
rlabel metal1 40 55 40 55 6 nq
rlabel metal1 35 94 35 94 6 vdd
rlabel metal1 35 94 35 94 6 vdd
rlabel polycontact 60 50 60 50 6 i1
rlabel polycontact 60 50 60 50 6 i1
<< end >>
