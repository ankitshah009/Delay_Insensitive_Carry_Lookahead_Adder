magic
tech scmos
timestamp 1179386007
<< checkpaint >>
rect -22 -25 54 105
<< ab >>
rect 0 0 32 80
<< pwell >>
rect -4 -7 36 36
<< nwell >>
rect -4 36 36 87
<< polysilicon >>
rect 10 66 12 71
rect 20 58 22 63
rect 10 39 12 42
rect 20 39 22 42
rect 9 38 23 39
rect 9 34 18 38
rect 22 34 23 38
rect 9 33 23 34
rect 9 30 11 33
rect 9 10 11 15
<< ndiffusion >>
rect 2 29 9 30
rect 2 25 3 29
rect 7 25 9 29
rect 2 22 9 25
rect 2 18 3 22
rect 7 18 9 22
rect 2 17 9 18
rect 4 15 9 17
rect 11 28 19 30
rect 11 24 13 28
rect 17 24 19 28
rect 11 20 19 24
rect 11 16 13 20
rect 17 16 19 20
rect 11 15 19 16
<< pdiffusion >>
rect 2 65 10 66
rect 2 61 4 65
rect 8 61 10 65
rect 2 57 10 61
rect 2 53 4 57
rect 8 53 10 57
rect 2 42 10 53
rect 12 58 17 66
rect 12 54 20 58
rect 12 50 14 54
rect 18 50 20 54
rect 12 47 20 50
rect 12 43 14 47
rect 18 43 20 47
rect 12 42 20 43
rect 22 57 30 58
rect 22 53 24 57
rect 28 53 30 57
rect 22 42 30 53
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect -2 68 34 78
rect 4 65 8 68
rect 4 57 8 61
rect 24 57 28 68
rect 4 52 8 53
rect 13 50 14 54
rect 18 50 19 54
rect 24 52 28 53
rect 13 47 19 50
rect 2 41 14 47
rect 18 43 19 47
rect 2 30 6 41
rect 26 39 30 47
rect 18 38 30 39
rect 22 34 30 38
rect 18 33 30 34
rect 2 29 7 30
rect 2 25 3 29
rect 2 22 7 25
rect 2 18 3 22
rect 2 17 7 18
rect 13 28 17 29
rect 13 20 17 24
rect 13 12 17 16
rect -2 2 34 12
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
<< ntransistor >>
rect 9 15 11 30
<< ptransistor >>
rect 10 42 12 66
rect 20 42 22 58
<< polycontact >>
rect 18 34 22 38
<< ndcontact >>
rect 3 25 7 29
rect 3 18 7 22
rect 13 24 17 28
rect 13 16 17 20
<< pdcontact >>
rect 4 61 8 65
rect 4 53 8 57
rect 14 50 18 54
rect 14 43 18 47
rect 24 53 28 57
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
<< psubstratepdiff >>
rect 0 2 32 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 32 2
rect 0 -3 32 -2
<< nsubstratendiff >>
rect 0 82 32 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 32 82
rect 0 77 32 78
<< labels >>
rlabel metal1 4 32 4 32 6 z
rlabel metal1 12 44 12 44 6 z
rlabel metal1 16 6 16 6 6 vss
rlabel polycontact 20 36 20 36 6 a
rlabel metal1 16 74 16 74 6 vdd
rlabel metal1 28 40 28 40 6 a
<< end >>
