magic
tech scmos
timestamp 1180640142
<< checkpaint >>
rect -24 -26 94 126
<< ab >>
rect 0 0 70 100
<< pwell >>
rect -4 -6 74 49
<< nwell >>
rect -4 49 74 106
<< polysilicon >>
rect 31 94 33 98
rect 39 94 41 98
rect 47 94 49 98
rect 55 94 57 98
rect 15 75 17 80
rect 15 49 17 55
rect 31 49 33 55
rect 39 52 41 55
rect 15 48 23 49
rect 15 45 18 48
rect 11 44 18 45
rect 22 44 23 48
rect 11 43 23 44
rect 27 48 33 49
rect 27 44 28 48
rect 32 44 33 48
rect 27 43 33 44
rect 37 51 43 52
rect 37 47 38 51
rect 42 47 43 51
rect 37 46 43 47
rect 11 33 13 43
rect 27 38 29 43
rect 37 39 39 46
rect 47 43 49 55
rect 55 52 57 55
rect 55 51 63 52
rect 55 49 58 51
rect 57 47 58 49
rect 62 47 63 51
rect 57 46 63 47
rect 47 42 53 43
rect 47 40 48 42
rect 23 36 29 38
rect 35 36 39 39
rect 45 38 48 40
rect 52 38 53 42
rect 45 37 53 38
rect 23 33 25 36
rect 35 33 37 36
rect 45 33 47 37
rect 57 33 59 46
rect 11 18 13 23
rect 23 22 25 27
rect 35 23 37 27
rect 45 22 47 27
rect 57 22 59 27
<< ndiffusion >>
rect 3 32 11 33
rect 3 28 4 32
rect 8 28 11 32
rect 3 27 11 28
rect 6 23 11 27
rect 13 27 23 33
rect 25 32 35 33
rect 25 28 28 32
rect 32 28 35 32
rect 25 27 35 28
rect 37 27 45 33
rect 47 32 57 33
rect 47 28 50 32
rect 54 28 57 32
rect 47 27 57 28
rect 59 32 67 33
rect 59 28 62 32
rect 66 28 67 32
rect 59 27 67 28
rect 13 23 21 27
rect 15 12 21 23
rect 39 21 43 27
rect 37 20 43 21
rect 37 16 38 20
rect 42 16 43 20
rect 37 15 43 16
rect 15 8 16 12
rect 20 8 21 12
rect 15 7 21 8
<< pdiffusion >>
rect 19 92 31 94
rect 19 88 22 92
rect 26 88 31 92
rect 19 75 31 88
rect 10 70 15 75
rect 7 69 15 70
rect 7 65 8 69
rect 12 65 15 69
rect 7 60 15 65
rect 7 56 8 60
rect 12 56 15 60
rect 7 55 15 56
rect 17 55 31 75
rect 33 55 39 94
rect 41 55 47 94
rect 49 55 55 94
rect 57 83 62 94
rect 57 82 65 83
rect 57 78 60 82
rect 64 78 65 82
rect 57 77 65 78
rect 57 55 62 77
<< metal1 >>
rect -2 92 72 100
rect -2 88 22 92
rect 26 88 72 92
rect 18 78 60 82
rect 64 78 65 82
rect 8 69 12 73
rect 8 60 12 65
rect 3 28 4 32
rect 8 22 12 56
rect 18 48 22 78
rect 27 68 42 73
rect 47 68 62 73
rect 18 32 22 44
rect 28 48 32 63
rect 38 51 42 68
rect 38 46 42 47
rect 28 42 32 44
rect 48 42 52 63
rect 58 51 62 68
rect 58 46 62 47
rect 28 37 43 42
rect 52 38 63 42
rect 48 37 63 38
rect 62 32 66 33
rect 18 28 28 32
rect 32 28 50 32
rect 54 28 55 32
rect 8 17 23 22
rect 38 20 42 21
rect 38 12 42 16
rect 62 12 66 28
rect -2 8 16 12
rect 20 8 72 12
rect -2 0 72 8
<< ntransistor >>
rect 11 23 13 33
rect 23 27 25 33
rect 35 27 37 33
rect 45 27 47 33
rect 57 27 59 33
<< ptransistor >>
rect 15 55 17 75
rect 31 55 33 94
rect 39 55 41 94
rect 47 55 49 94
rect 55 55 57 94
<< polycontact >>
rect 18 44 22 48
rect 28 44 32 48
rect 38 47 42 51
rect 58 47 62 51
rect 48 38 52 42
<< ndcontact >>
rect 4 28 8 32
rect 28 28 32 32
rect 50 28 54 32
rect 62 28 66 32
rect 38 16 42 20
rect 16 8 20 12
<< pdcontact >>
rect 22 88 26 92
rect 8 65 12 69
rect 8 56 12 60
rect 60 78 64 82
<< psubstratepcontact >>
rect 48 4 52 8
rect 58 4 62 8
<< nsubstratencontact >>
rect 8 92 12 96
<< psubstratepdiff >>
rect 47 8 63 9
rect 47 4 48 8
rect 52 4 58 8
rect 62 4 63 8
rect 47 3 63 4
<< nsubstratendiff >>
rect 7 96 13 97
rect 7 92 8 96
rect 12 92 13 96
rect 7 91 13 92
<< labels >>
rlabel polycontact 19 46 19 46 6 zn
rlabel metal1 20 20 20 20 6 z
rlabel metal1 20 20 20 20 6 z
rlabel metal1 10 45 10 45 6 z
rlabel metal1 10 45 10 45 6 z
rlabel metal1 20 55 20 55 6 zn
rlabel metal1 35 6 35 6 6 vss
rlabel metal1 35 6 35 6 6 vss
rlabel metal1 30 50 30 50 6 a
rlabel metal1 30 50 30 50 6 a
rlabel metal1 30 70 30 70 6 b
rlabel metal1 30 70 30 70 6 b
rlabel metal1 35 94 35 94 6 vdd
rlabel metal1 35 94 35 94 6 vdd
rlabel metal1 36 30 36 30 6 zn
rlabel metal1 40 40 40 40 6 a
rlabel metal1 40 40 40 40 6 a
rlabel metal1 50 50 50 50 6 c
rlabel metal1 50 50 50 50 6 c
rlabel metal1 40 60 40 60 6 b
rlabel metal1 40 60 40 60 6 b
rlabel metal1 50 70 50 70 6 d
rlabel metal1 50 70 50 70 6 d
rlabel metal1 60 40 60 40 6 c
rlabel metal1 60 40 60 40 6 c
rlabel metal1 60 60 60 60 6 d
rlabel metal1 60 60 60 60 6 d
rlabel metal1 41 80 41 80 6 zn
<< end >>
