.subckt xor2v1x1 a b vdd vss z
*   SPICE3 file   created from xor2v1x1.ext -      technology: scmos
m00 an     a      vdd    vdd p w=22u  l=2.3636u ad=88p      pd=30u      as=110p     ps=39.3333u
m01 z      bn     an     vdd p w=22u  l=2.3636u ad=88p      pd=30u      as=88p      ps=30u
m02 ai     b      z      vdd p w=22u  l=2.3636u ad=88p      pd=30u      as=88p      ps=30u
m03 vdd    an     ai     vdd p w=22u  l=2.3636u ad=110p     pd=39.3333u as=88p      ps=30u
m04 bn     b      vdd    vdd p w=22u  l=2.3636u ad=122p     pd=58u      as=110p     ps=39.3333u
m05 an     a      vss    vss n w=11u  l=2.3636u ad=45p      pd=20u      as=99p      ps=32.6667u
m06 z      b      an     vss n w=11u  l=2.3636u ad=44p      pd=19u      as=45p      ps=20u
m07 ai     bn     z      vss n w=11u  l=2.3636u ad=44p      pd=19u      as=44p      ps=19u
m08 vss    an     ai     vss n w=11u  l=2.3636u ad=99p      pd=32.6667u as=44p      ps=19u
m09 bn     b      vss    vss n w=11u  l=2.3636u ad=67p      pd=36u      as=99p      ps=32.6667u
C0  z      an     0.285f
C1  ai     b      0.067f
C2  vss    a      0.028f
C3  ai     bn     0.103f
C4  z      a      0.026f
C5  vdd    b      0.051f
C6  vdd    bn     0.308f
C7  an     a      0.106f
C8  vss    ai     0.024f
C9  b      bn     0.310f
C10 ai     z      0.151f
C11 vss    vdd    0.005f
C12 ai     an     0.243f
C13 z      vdd    0.017f
C14 vss    b      0.037f
C15 vdd    an     0.028f
C16 ai     a      0.014f
C17 vss    bn     0.072f
C18 z      b      0.031f
C19 vdd    a      0.018f
C20 z      bn     0.126f
C21 an     b      0.188f
C22 an     bn     0.212f
C23 b      a      0.026f
C24 vss    z      0.025f
C25 a      bn     0.098f
C26 ai     vdd    0.012f
C27 vss    an     0.329f
C29 ai     vss    0.008f
C30 z      vss    0.009f
C32 an     vss    0.026f
C33 b      vss    0.056f
C34 a      vss    0.025f
C35 bn     vss    0.051f
.ends
