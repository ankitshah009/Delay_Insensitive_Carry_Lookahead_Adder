magic
tech scmos
timestamp 1179386711
<< checkpaint >>
rect -22 -25 158 105
<< ab >>
rect 0 0 136 80
<< pwell >>
rect -4 -7 140 36
<< nwell >>
rect -4 36 140 87
<< polysilicon >>
rect 9 70 11 74
rect 16 70 18 74
rect 26 70 28 74
rect 33 70 35 74
rect 43 70 45 74
rect 50 70 52 74
rect 60 70 62 74
rect 67 70 69 74
rect 77 70 79 74
rect 84 70 86 74
rect 94 70 96 74
rect 101 70 103 74
rect 111 70 113 74
rect 121 61 123 65
rect 9 33 11 42
rect 16 39 18 42
rect 26 39 28 42
rect 33 39 35 42
rect 43 39 45 42
rect 50 39 52 42
rect 60 39 62 42
rect 67 39 69 42
rect 77 39 79 42
rect 16 38 29 39
rect 16 37 24 38
rect 23 34 24 37
rect 28 34 29 38
rect 33 38 45 39
rect 33 37 40 38
rect 23 33 29 34
rect 9 32 19 33
rect 9 31 14 32
rect 13 28 14 31
rect 18 28 19 32
rect 13 27 19 28
rect 17 24 19 27
rect 27 24 29 33
rect 39 34 40 37
rect 44 34 45 38
rect 39 33 45 34
rect 49 38 63 39
rect 49 34 50 38
rect 54 34 63 38
rect 49 33 63 34
rect 67 38 79 39
rect 67 34 68 38
rect 72 37 79 38
rect 84 39 86 42
rect 94 39 96 42
rect 101 39 103 42
rect 111 39 113 42
rect 121 39 123 42
rect 84 38 96 39
rect 72 34 73 37
rect 67 33 73 34
rect 84 34 85 38
rect 89 37 96 38
rect 100 38 106 39
rect 89 34 90 37
rect 84 33 90 34
rect 100 34 101 38
rect 105 34 106 38
rect 100 33 106 34
rect 110 38 123 39
rect 110 34 115 38
rect 119 34 123 38
rect 110 33 123 34
rect 39 30 41 33
rect 49 30 51 33
rect 61 30 63 33
rect 71 30 73 33
rect 110 27 112 33
rect 120 27 122 33
rect 17 8 19 13
rect 27 8 29 13
rect 39 8 41 13
rect 49 8 51 13
rect 61 8 63 13
rect 71 8 73 13
rect 110 10 112 15
rect 120 10 122 15
<< ndiffusion >>
rect 31 24 39 30
rect 8 13 17 24
rect 19 22 27 24
rect 19 18 21 22
rect 25 18 27 22
rect 19 13 27 18
rect 29 13 39 24
rect 41 22 49 30
rect 41 18 43 22
rect 47 18 49 22
rect 41 13 49 18
rect 51 13 61 30
rect 63 22 71 30
rect 63 18 65 22
rect 69 18 71 22
rect 63 13 71 18
rect 73 18 81 30
rect 73 14 75 18
rect 79 14 81 18
rect 103 20 110 27
rect 103 16 104 20
rect 108 16 110 20
rect 103 15 110 16
rect 112 26 120 27
rect 112 22 114 26
rect 118 22 120 26
rect 112 15 120 22
rect 122 20 130 27
rect 122 16 124 20
rect 128 16 130 20
rect 122 15 130 16
rect 73 13 81 14
rect 8 12 15 13
rect 8 8 10 12
rect 14 8 15 12
rect 31 12 37 13
rect 31 8 32 12
rect 36 8 37 12
rect 53 12 59 13
rect 53 8 54 12
rect 58 8 59 12
rect 8 7 15 8
rect 31 7 37 8
rect 53 7 59 8
<< pdiffusion >>
rect 2 69 9 70
rect 2 65 3 69
rect 7 65 9 69
rect 2 62 9 65
rect 2 58 3 62
rect 7 58 9 62
rect 2 42 9 58
rect 11 42 16 70
rect 18 62 26 70
rect 18 58 20 62
rect 24 58 26 62
rect 18 54 26 58
rect 18 50 20 54
rect 24 50 26 54
rect 18 42 26 50
rect 28 42 33 70
rect 35 69 43 70
rect 35 65 37 69
rect 41 65 43 69
rect 35 62 43 65
rect 35 58 37 62
rect 41 58 43 62
rect 35 42 43 58
rect 45 42 50 70
rect 52 61 60 70
rect 52 57 54 61
rect 58 57 60 61
rect 52 54 60 57
rect 52 50 54 54
rect 58 50 60 54
rect 52 42 60 50
rect 62 42 67 70
rect 69 69 77 70
rect 69 65 71 69
rect 75 65 77 69
rect 69 62 77 65
rect 69 58 71 62
rect 75 58 77 62
rect 69 42 77 58
rect 79 42 84 70
rect 86 62 94 70
rect 86 58 88 62
rect 92 58 94 62
rect 86 54 94 58
rect 86 50 88 54
rect 92 50 94 54
rect 86 42 94 50
rect 96 42 101 70
rect 103 69 111 70
rect 103 65 105 69
rect 109 65 111 69
rect 103 62 111 65
rect 103 58 105 62
rect 109 58 111 62
rect 103 55 111 58
rect 103 51 105 55
rect 109 51 111 55
rect 103 42 111 51
rect 113 61 118 70
rect 113 54 121 61
rect 113 50 115 54
rect 119 50 121 54
rect 113 47 121 50
rect 113 43 115 47
rect 119 43 121 47
rect 113 42 121 43
rect 123 60 130 61
rect 123 56 125 60
rect 129 56 130 60
rect 123 53 130 56
rect 123 49 125 53
rect 129 49 130 53
rect 123 42 130 49
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect 118 78 122 82
rect 126 78 130 82
rect 134 78 138 82
rect -2 69 138 78
rect -2 68 3 69
rect 2 65 3 68
rect 7 68 37 69
rect 7 65 8 68
rect 2 62 8 65
rect 36 65 37 68
rect 41 68 71 69
rect 41 65 42 68
rect 2 58 3 62
rect 7 58 8 62
rect 18 62 24 63
rect 18 58 20 62
rect 36 62 42 65
rect 70 65 71 68
rect 75 68 105 69
rect 75 65 76 68
rect 70 62 76 65
rect 109 68 138 69
rect 36 58 37 62
rect 41 58 42 62
rect 54 61 58 62
rect 18 54 24 58
rect 70 58 71 62
rect 75 58 76 62
rect 88 62 94 63
rect 92 58 94 62
rect 54 54 58 57
rect 88 54 94 58
rect 2 50 20 54
rect 24 50 54 54
rect 58 50 88 54
rect 92 50 94 54
rect 105 62 109 65
rect 105 55 109 58
rect 124 60 130 68
rect 124 56 125 60
rect 129 56 130 60
rect 105 50 109 51
rect 115 54 119 55
rect 2 22 6 50
rect 115 47 119 50
rect 124 53 130 56
rect 124 49 125 53
rect 129 49 130 53
rect 25 42 87 46
rect 25 38 31 42
rect 49 38 55 42
rect 81 38 87 42
rect 101 43 115 46
rect 101 42 119 43
rect 101 38 105 42
rect 23 34 24 38
rect 28 34 31 38
rect 39 34 40 38
rect 44 34 45 38
rect 49 34 50 38
rect 54 34 55 38
rect 67 34 68 38
rect 72 34 73 38
rect 81 34 85 38
rect 89 34 95 38
rect 113 34 115 38
rect 119 34 127 38
rect 14 32 18 33
rect 39 30 45 34
rect 67 30 73 34
rect 101 30 105 34
rect 18 28 118 30
rect 14 26 118 28
rect 122 25 127 34
rect 2 18 21 22
rect 25 18 43 22
rect 47 18 65 22
rect 69 18 71 22
rect 114 21 118 22
rect 104 20 108 21
rect 75 18 79 19
rect 75 12 79 14
rect 104 12 108 16
rect 124 20 128 21
rect 124 12 128 16
rect -2 8 10 12
rect 14 8 32 12
rect 36 8 54 12
rect 58 8 138 12
rect -2 2 138 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 122 2
rect 126 -2 130 2
rect 134 -2 138 2
<< ntransistor >>
rect 17 13 19 24
rect 27 13 29 24
rect 39 13 41 30
rect 49 13 51 30
rect 61 13 63 30
rect 71 13 73 30
rect 110 15 112 27
rect 120 15 122 27
<< ptransistor >>
rect 9 42 11 70
rect 16 42 18 70
rect 26 42 28 70
rect 33 42 35 70
rect 43 42 45 70
rect 50 42 52 70
rect 60 42 62 70
rect 67 42 69 70
rect 77 42 79 70
rect 84 42 86 70
rect 94 42 96 70
rect 101 42 103 70
rect 111 42 113 70
rect 121 42 123 61
<< polycontact >>
rect 24 34 28 38
rect 14 28 18 32
rect 40 34 44 38
rect 50 34 54 38
rect 68 34 72 38
rect 85 34 89 38
rect 101 34 105 38
rect 115 34 119 38
<< ndcontact >>
rect 21 18 25 22
rect 43 18 47 22
rect 65 18 69 22
rect 75 14 79 18
rect 104 16 108 20
rect 114 22 118 26
rect 124 16 128 20
rect 10 8 14 12
rect 32 8 36 12
rect 54 8 58 12
<< pdcontact >>
rect 3 65 7 69
rect 3 58 7 62
rect 20 58 24 62
rect 20 50 24 54
rect 37 65 41 69
rect 37 58 41 62
rect 54 57 58 61
rect 54 50 58 54
rect 71 65 75 69
rect 71 58 75 62
rect 88 58 92 62
rect 88 50 92 54
rect 105 65 109 69
rect 105 58 109 62
rect 105 51 109 55
rect 115 50 119 54
rect 115 43 119 47
rect 125 56 129 60
rect 125 49 129 53
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
rect 90 -2 94 2
rect 98 -2 102 2
rect 106 -2 110 2
rect 114 -2 118 2
rect 122 -2 126 2
rect 130 -2 134 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
rect 90 78 94 82
rect 98 78 102 82
rect 106 78 110 82
rect 114 78 118 82
rect 122 78 126 82
rect 130 78 134 82
<< psubstratepdiff >>
rect 0 2 136 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 122 2
rect 126 -2 130 2
rect 134 -2 136 2
rect 0 -3 136 -2
<< nsubstratendiff >>
rect 0 82 136 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect 118 78 122 82
rect 126 78 130 82
rect 134 78 136 82
rect 0 77 136 78
<< labels >>
rlabel polycontact 16 30 16 30 6 an
rlabel polycontact 42 36 42 36 6 an
rlabel polycontact 70 36 70 36 6 an
rlabel ptransistor 102 53 102 53 6 an
rlabel metal1 12 20 12 20 6 z
rlabel metal1 20 20 20 20 6 z
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 52 12 52 6 z
rlabel metal1 20 56 20 56 6 z
rlabel metal1 28 20 28 20 6 z
rlabel metal1 36 20 36 20 6 z
rlabel ndcontact 44 20 44 20 6 z
rlabel metal1 42 32 42 32 6 an
rlabel metal1 28 40 28 40 6 b
rlabel metal1 36 44 36 44 6 b
rlabel metal1 44 44 44 44 6 b
rlabel metal1 36 52 36 52 6 z
rlabel metal1 44 52 44 52 6 z
rlabel metal1 28 52 28 52 6 z
rlabel metal1 68 6 68 6 6 vss
rlabel metal1 52 20 52 20 6 z
rlabel metal1 60 20 60 20 6 z
rlabel ndcontact 68 20 68 20 6 z
rlabel metal1 70 32 70 32 6 an
rlabel metal1 52 40 52 40 6 b
rlabel metal1 60 44 60 44 6 b
rlabel metal1 68 44 68 44 6 b
rlabel metal1 76 44 76 44 6 b
rlabel metal1 60 52 60 52 6 z
rlabel metal1 68 52 68 52 6 z
rlabel metal1 76 52 76 52 6 z
rlabel metal1 52 52 52 52 6 z
rlabel metal1 68 74 68 74 6 vdd
rlabel polycontact 103 36 103 36 6 an
rlabel metal1 84 40 84 40 6 b
rlabel metal1 92 36 92 36 6 b
rlabel metal1 84 52 84 52 6 z
rlabel metal1 92 60 92 60 6 z
rlabel metal1 66 28 66 28 6 an
rlabel ndcontact 116 25 116 25 6 an
rlabel metal1 124 32 124 32 6 a
rlabel polycontact 116 36 116 36 6 a
rlabel metal1 117 48 117 48 6 an
<< end >>
