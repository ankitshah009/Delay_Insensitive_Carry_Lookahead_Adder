magic
tech scmos
timestamp 1179386626
<< checkpaint >>
rect -22 -25 150 105
<< ab >>
rect 0 0 128 80
<< pwell >>
rect -4 -7 132 36
<< nwell >>
rect -4 36 132 87
<< polysilicon >>
rect 9 70 11 74
rect 19 70 21 74
rect 40 69 42 74
rect 50 69 52 74
rect 60 69 62 74
rect 70 69 72 74
rect 97 69 99 74
rect 107 69 109 74
rect 117 69 119 74
rect 9 39 11 43
rect 19 39 21 43
rect 40 39 42 42
rect 50 39 52 42
rect 60 39 62 42
rect 70 39 72 42
rect 97 39 99 42
rect 107 39 109 42
rect 117 39 119 42
rect 2 38 11 39
rect 2 34 3 38
rect 7 34 11 38
rect 2 33 11 34
rect 9 30 11 33
rect 16 38 23 39
rect 16 34 18 38
rect 22 35 23 38
rect 33 38 45 39
rect 22 34 28 35
rect 16 33 28 34
rect 16 30 18 33
rect 26 30 28 33
rect 33 34 34 38
rect 38 34 45 38
rect 33 33 45 34
rect 33 30 35 33
rect 43 30 45 33
rect 50 38 62 39
rect 50 34 51 38
rect 55 34 62 38
rect 50 33 62 34
rect 50 30 52 33
rect 60 30 62 33
rect 67 38 73 39
rect 67 34 68 38
rect 72 34 73 38
rect 97 38 119 39
rect 97 35 98 38
rect 67 33 73 34
rect 77 34 98 35
rect 102 34 106 38
rect 110 34 119 38
rect 77 33 119 34
rect 67 30 69 33
rect 77 30 79 33
rect 87 30 89 33
rect 97 30 99 33
rect 107 30 109 33
rect 117 30 119 33
rect 107 15 109 20
rect 117 15 119 20
rect 9 6 11 10
rect 16 6 18 10
rect 26 6 28 10
rect 33 6 35 10
rect 43 6 45 10
rect 50 6 52 10
rect 60 6 62 10
rect 67 6 69 10
rect 77 6 79 10
rect 87 6 89 10
rect 97 6 99 10
<< ndiffusion >>
rect 2 29 9 30
rect 2 25 3 29
rect 7 25 9 29
rect 2 22 9 25
rect 2 18 3 22
rect 7 18 9 22
rect 2 17 9 18
rect 4 10 9 17
rect 11 10 16 30
rect 18 15 26 30
rect 18 11 20 15
rect 24 11 26 15
rect 18 10 26 11
rect 28 10 33 30
rect 35 22 43 30
rect 35 18 37 22
rect 41 18 43 22
rect 35 10 43 18
rect 45 10 50 30
rect 52 15 60 30
rect 52 11 54 15
rect 58 11 60 15
rect 52 10 60 11
rect 62 10 67 30
rect 69 29 77 30
rect 69 25 71 29
rect 75 25 77 29
rect 69 22 77 25
rect 69 18 71 22
rect 75 18 77 22
rect 69 10 77 18
rect 79 29 87 30
rect 79 25 81 29
rect 85 25 87 29
rect 79 10 87 25
rect 89 22 97 30
rect 89 18 91 22
rect 95 18 97 22
rect 89 10 97 18
rect 99 29 107 30
rect 99 25 101 29
rect 105 25 107 29
rect 99 20 107 25
rect 109 25 117 30
rect 109 21 111 25
rect 115 21 117 25
rect 109 20 117 21
rect 119 29 126 30
rect 119 25 121 29
rect 125 25 126 29
rect 119 24 126 25
rect 119 20 124 24
rect 99 10 104 20
<< pdiffusion >>
rect 2 69 9 70
rect 2 65 3 69
rect 7 65 9 69
rect 2 62 9 65
rect 2 58 3 62
rect 7 58 9 62
rect 2 43 9 58
rect 11 62 19 70
rect 11 58 13 62
rect 17 58 19 62
rect 11 55 19 58
rect 11 51 13 55
rect 17 51 19 55
rect 11 43 19 51
rect 21 69 28 70
rect 21 65 23 69
rect 27 65 28 69
rect 21 62 28 65
rect 21 58 23 62
rect 27 58 28 62
rect 21 43 28 58
rect 33 68 40 69
rect 33 64 34 68
rect 38 64 40 68
rect 33 61 40 64
rect 33 57 34 61
rect 38 57 40 61
rect 33 42 40 57
rect 42 61 50 69
rect 42 57 44 61
rect 48 57 50 61
rect 42 54 50 57
rect 42 50 44 54
rect 48 50 50 54
rect 42 42 50 50
rect 52 68 60 69
rect 52 64 54 68
rect 58 64 60 68
rect 52 61 60 64
rect 52 57 54 61
rect 58 57 60 61
rect 52 42 60 57
rect 62 61 70 69
rect 62 57 64 61
rect 68 57 70 61
rect 62 54 70 57
rect 62 50 64 54
rect 68 50 70 54
rect 62 42 70 50
rect 72 63 77 69
rect 92 63 97 69
rect 72 62 97 63
rect 72 58 74 62
rect 78 58 82 62
rect 86 58 91 62
rect 95 58 97 62
rect 72 42 97 58
rect 99 61 107 69
rect 99 57 101 61
rect 105 57 107 61
rect 99 54 107 57
rect 99 50 101 54
rect 105 50 107 54
rect 99 42 107 50
rect 109 68 117 69
rect 109 64 111 68
rect 115 64 117 68
rect 109 61 117 64
rect 109 57 111 61
rect 115 57 117 61
rect 109 42 117 57
rect 119 55 124 69
rect 119 54 126 55
rect 119 50 121 54
rect 125 50 126 54
rect 119 47 126 50
rect 119 43 121 47
rect 125 43 126 47
rect 119 42 126 43
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect 118 78 122 82
rect 126 78 130 82
rect -2 69 130 78
rect -2 68 3 69
rect 2 65 3 68
rect 7 68 23 69
rect 7 65 8 68
rect 2 62 8 65
rect 22 65 23 68
rect 27 68 130 69
rect 27 65 28 68
rect 2 58 3 62
rect 7 58 8 62
rect 13 62 17 63
rect 22 62 28 65
rect 22 58 23 62
rect 27 58 28 62
rect 33 64 34 68
rect 38 64 39 68
rect 33 61 39 64
rect 53 64 54 68
rect 58 64 59 68
rect 13 55 17 58
rect 33 57 34 61
rect 38 57 39 61
rect 44 61 48 62
rect 53 61 59 64
rect 53 57 54 61
rect 58 57 59 61
rect 64 61 70 63
rect 68 57 70 61
rect 73 62 79 68
rect 90 62 96 68
rect 110 64 111 68
rect 115 64 116 68
rect 73 58 74 62
rect 78 58 82 62
rect 86 58 91 62
rect 95 58 96 62
rect 101 61 105 62
rect 2 46 6 55
rect 44 54 48 57
rect 64 54 70 57
rect 110 61 116 64
rect 110 57 111 61
rect 115 57 116 61
rect 101 54 105 57
rect 121 54 126 55
rect 17 51 44 54
rect 13 50 44 51
rect 48 50 64 54
rect 68 50 101 54
rect 105 50 121 54
rect 125 50 126 54
rect 2 42 64 46
rect 2 38 7 42
rect 33 38 39 42
rect 60 38 64 42
rect 2 34 3 38
rect 17 34 18 38
rect 22 34 29 38
rect 33 34 34 38
rect 38 34 39 38
rect 43 34 51 38
rect 55 34 56 38
rect 60 34 68 38
rect 72 34 73 38
rect 2 33 7 34
rect 25 30 29 34
rect 43 30 47 34
rect 82 30 86 50
rect 121 47 126 50
rect 97 38 103 46
rect 125 43 126 47
rect 97 34 98 38
rect 102 34 106 38
rect 110 34 111 38
rect 2 25 3 29
rect 7 25 8 29
rect 25 26 47 30
rect 71 29 75 30
rect 2 22 8 25
rect 80 29 106 30
rect 80 25 81 29
rect 85 25 101 29
rect 105 25 106 29
rect 121 29 126 43
rect 111 25 115 26
rect 71 22 75 25
rect 2 18 3 22
rect 7 18 37 22
rect 41 18 71 22
rect 75 18 91 22
rect 95 21 111 22
rect 95 18 115 21
rect 125 25 126 29
rect 121 17 126 25
rect 19 12 20 15
rect -2 11 20 12
rect 24 12 25 15
rect 53 12 54 15
rect 24 11 54 12
rect 58 12 59 15
rect 58 11 130 12
rect -2 2 130 11
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 122 2
rect 126 -2 130 2
<< ntransistor >>
rect 9 10 11 30
rect 16 10 18 30
rect 26 10 28 30
rect 33 10 35 30
rect 43 10 45 30
rect 50 10 52 30
rect 60 10 62 30
rect 67 10 69 30
rect 77 10 79 30
rect 87 10 89 30
rect 97 10 99 30
rect 107 20 109 30
rect 117 20 119 30
<< ptransistor >>
rect 9 43 11 70
rect 19 43 21 70
rect 40 42 42 69
rect 50 42 52 69
rect 60 42 62 69
rect 70 42 72 69
rect 97 42 99 69
rect 107 42 109 69
rect 117 42 119 69
<< polycontact >>
rect 3 34 7 38
rect 18 34 22 38
rect 34 34 38 38
rect 51 34 55 38
rect 68 34 72 38
rect 98 34 102 38
rect 106 34 110 38
<< ndcontact >>
rect 3 25 7 29
rect 3 18 7 22
rect 20 11 24 15
rect 37 18 41 22
rect 54 11 58 15
rect 71 25 75 29
rect 71 18 75 22
rect 81 25 85 29
rect 91 18 95 22
rect 101 25 105 29
rect 111 21 115 25
rect 121 25 125 29
<< pdcontact >>
rect 3 65 7 69
rect 3 58 7 62
rect 13 58 17 62
rect 13 51 17 55
rect 23 65 27 69
rect 23 58 27 62
rect 34 64 38 68
rect 34 57 38 61
rect 44 57 48 61
rect 44 50 48 54
rect 54 64 58 68
rect 54 57 58 61
rect 64 57 68 61
rect 64 50 68 54
rect 74 58 78 62
rect 82 58 86 62
rect 91 58 95 62
rect 101 57 105 61
rect 101 50 105 54
rect 111 64 115 68
rect 111 57 115 61
rect 121 50 125 54
rect 121 43 125 47
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
rect 90 -2 94 2
rect 98 -2 102 2
rect 106 -2 110 2
rect 114 -2 118 2
rect 122 -2 126 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
rect 90 78 94 82
rect 98 78 102 82
rect 106 78 110 82
rect 114 78 118 82
rect 122 78 126 82
<< psubstratepdiff >>
rect 0 2 128 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 122 2
rect 126 -2 128 2
rect 0 -3 128 -2
<< nsubstratendiff >>
rect 0 82 128 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect 118 78 122 82
rect 126 78 128 82
rect 0 77 128 78
<< labels >>
rlabel metal1 5 23 5 23 6 n2
rlabel metal1 12 44 12 44 6 b
rlabel metal1 4 44 4 44 6 b
rlabel metal1 28 28 28 28 6 a
rlabel metal1 36 28 36 28 6 a
rlabel polycontact 20 36 20 36 6 a
rlabel metal1 28 44 28 44 6 b
rlabel metal1 36 40 36 40 6 b
rlabel metal1 20 44 20 44 6 b
rlabel metal1 20 52 20 52 6 z
rlabel metal1 28 52 28 52 6 z
rlabel metal1 36 52 36 52 6 z
rlabel metal1 44 28 44 28 6 a
rlabel polycontact 52 36 52 36 6 a
rlabel metal1 52 44 52 44 6 b
rlabel metal1 60 44 60 44 6 b
rlabel metal1 44 44 44 44 6 b
rlabel metal1 44 52 44 52 6 z
rlabel metal1 52 52 52 52 6 z
rlabel metal1 60 52 60 52 6 z
rlabel metal1 64 6 64 6 6 vss
rlabel metal1 73 24 73 24 6 n2
rlabel metal1 68 36 68 36 6 b
rlabel metal1 84 40 84 40 6 z
rlabel metal1 76 52 76 52 6 z
rlabel metal1 68 56 68 56 6 z
rlabel metal1 64 74 64 74 6 vdd
rlabel metal1 92 28 92 28 6 z
rlabel metal1 100 28 100 28 6 z
rlabel metal1 100 40 100 40 6 c
rlabel metal1 92 52 92 52 6 z
rlabel metal1 100 52 100 52 6 z
rlabel metal1 58 20 58 20 6 n2
rlabel ndcontact 113 22 113 22 6 n2
rlabel polycontact 108 36 108 36 6 c
rlabel metal1 124 36 124 36 6 z
rlabel metal1 108 52 108 52 6 z
rlabel metal1 116 52 116 52 6 z
<< end >>
