magic
tech scmos
timestamp 1179385357
<< checkpaint >>
rect -22 -22 78 94
<< ab >>
rect 0 0 56 72
<< pwell >>
rect -4 -4 60 32
<< nwell >>
rect -4 32 60 76
<< polysilicon >>
rect 9 66 11 70
rect 19 66 21 70
rect 29 66 31 70
rect 39 66 41 70
rect 9 29 11 39
rect 19 36 21 39
rect 29 36 31 39
rect 19 35 25 36
rect 19 31 20 35
rect 24 31 25 35
rect 19 30 25 31
rect 29 35 35 36
rect 29 31 30 35
rect 34 31 35 35
rect 29 30 35 31
rect 39 35 41 39
rect 39 34 47 35
rect 39 30 42 34
rect 46 30 47 34
rect 9 28 15 29
rect 9 24 10 28
rect 14 24 15 28
rect 23 26 25 30
rect 31 26 33 30
rect 39 29 47 30
rect 39 26 41 29
rect 9 23 15 24
rect 13 20 15 23
rect 13 8 15 13
rect 23 5 25 10
rect 31 5 33 10
rect 39 5 41 10
<< ndiffusion >>
rect 18 20 23 26
rect 4 13 13 20
rect 15 18 23 20
rect 15 14 17 18
rect 21 14 23 18
rect 15 13 23 14
rect 4 8 11 13
rect 18 10 23 13
rect 25 10 31 26
rect 33 10 39 26
rect 41 15 48 26
rect 41 11 43 15
rect 47 11 48 15
rect 41 10 48 11
rect 4 4 6 8
rect 10 4 11 8
rect 4 3 11 4
<< pdiffusion >>
rect 4 60 9 66
rect 2 59 9 60
rect 2 55 3 59
rect 7 55 9 59
rect 2 51 9 55
rect 2 47 3 51
rect 7 47 9 51
rect 2 46 9 47
rect 4 39 9 46
rect 11 58 19 66
rect 11 54 13 58
rect 17 54 19 58
rect 11 51 19 54
rect 11 47 13 51
rect 17 47 19 51
rect 11 39 19 47
rect 21 65 29 66
rect 21 61 23 65
rect 27 61 29 65
rect 21 58 29 61
rect 21 54 23 58
rect 27 54 29 58
rect 21 39 29 54
rect 31 58 39 66
rect 31 54 33 58
rect 37 54 39 58
rect 31 51 39 54
rect 31 47 33 51
rect 37 47 39 51
rect 31 39 39 47
rect 41 65 48 66
rect 41 61 43 65
rect 47 61 48 65
rect 41 58 48 61
rect 41 54 43 58
rect 47 54 48 58
rect 41 39 48 54
<< metal1 >>
rect -2 65 58 72
rect -2 64 23 65
rect 22 61 23 64
rect 27 64 43 65
rect 27 61 28 64
rect 2 55 3 59
rect 7 55 8 59
rect 2 51 8 55
rect 2 47 3 51
rect 7 47 8 51
rect 13 58 17 59
rect 22 58 28 61
rect 42 61 43 64
rect 47 64 58 65
rect 47 61 48 64
rect 22 54 23 58
rect 27 54 28 58
rect 33 58 37 59
rect 42 58 48 61
rect 42 54 43 58
rect 47 54 48 58
rect 13 51 17 54
rect 33 51 37 54
rect 17 47 33 50
rect 2 18 6 47
rect 13 46 37 47
rect 10 37 24 43
rect 41 42 47 50
rect 17 35 24 37
rect 17 31 20 35
rect 29 38 47 42
rect 29 35 35 38
rect 29 31 30 35
rect 34 31 35 35
rect 17 30 24 31
rect 41 30 42 34
rect 46 30 47 34
rect 10 28 14 29
rect 41 27 47 30
rect 14 24 30 26
rect 10 22 30 24
rect 2 14 17 18
rect 21 14 22 18
rect 2 13 22 14
rect 26 13 30 22
rect 34 21 47 27
rect 43 15 47 16
rect 43 8 47 11
rect -2 4 6 8
rect 10 4 58 8
rect -2 0 58 4
<< ntransistor >>
rect 13 13 15 20
rect 23 10 25 26
rect 31 10 33 26
rect 39 10 41 26
<< ptransistor >>
rect 9 39 11 66
rect 19 39 21 66
rect 29 39 31 66
rect 39 39 41 66
<< polycontact >>
rect 20 31 24 35
rect 30 31 34 35
rect 42 30 46 34
rect 10 24 14 28
<< ndcontact >>
rect 17 14 21 18
rect 43 11 47 15
rect 6 4 10 8
<< pdcontact >>
rect 3 55 7 59
rect 3 47 7 51
rect 13 54 17 58
rect 13 47 17 51
rect 23 61 27 65
rect 23 54 27 58
rect 33 54 37 58
rect 33 47 37 51
rect 43 61 47 65
rect 43 54 47 58
<< labels >>
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 16 12 16 6 z
rlabel metal1 20 24 20 24 6 b
rlabel metal1 20 36 20 36 6 a3
rlabel metal1 12 40 12 40 6 a3
rlabel metal1 15 52 15 52 6 n3
rlabel metal1 28 4 28 4 6 vss
rlabel metal1 28 16 28 16 6 b
rlabel metal1 36 24 36 24 6 a1
rlabel metal1 36 40 36 40 6 a2
rlabel metal1 35 52 35 52 6 n3
rlabel metal1 28 68 28 68 6 vdd
rlabel metal1 44 28 44 28 6 a1
rlabel metal1 44 44 44 44 6 a2
<< end >>
