magic
tech scmos
timestamp 1179387097
<< checkpaint >>
rect -22 -22 94 94
<< ab >>
rect 0 0 72 72
<< pwell >>
rect -4 -4 76 32
<< nwell >>
rect -4 32 76 76
<< polysilicon >>
rect 11 63 13 68
rect 18 63 20 68
rect 28 63 30 68
rect 35 63 37 68
rect 47 62 49 67
rect 57 62 59 67
rect 11 44 13 47
rect 3 43 13 44
rect 3 39 4 43
rect 8 42 13 43
rect 8 39 9 42
rect 3 38 9 39
rect 18 37 20 47
rect 28 43 30 47
rect 35 44 37 47
rect 47 44 49 49
rect 57 46 59 49
rect 57 45 64 46
rect 35 43 53 44
rect 13 35 20 37
rect 25 42 31 43
rect 25 38 26 42
rect 30 38 31 42
rect 25 37 31 38
rect 35 42 48 43
rect 13 34 15 35
rect 9 33 15 34
rect 9 29 10 33
rect 14 29 15 33
rect 25 31 27 37
rect 35 31 37 42
rect 47 39 48 42
rect 52 39 53 43
rect 57 41 59 45
rect 63 41 64 45
rect 57 40 64 41
rect 47 38 53 39
rect 51 35 53 38
rect 9 28 15 29
rect 13 25 15 28
rect 23 28 27 31
rect 33 28 37 31
rect 41 33 47 34
rect 51 33 56 35
rect 41 29 42 33
rect 46 29 47 33
rect 41 28 47 29
rect 23 25 25 28
rect 33 25 35 28
rect 43 25 45 28
rect 54 25 56 33
rect 61 25 63 40
rect 13 13 15 18
rect 23 13 25 18
rect 33 13 35 18
rect 43 13 45 18
rect 54 9 56 14
rect 61 9 63 14
<< ndiffusion >>
rect 4 18 13 25
rect 15 23 23 25
rect 15 19 17 23
rect 21 19 23 23
rect 15 18 23 19
rect 25 24 33 25
rect 25 20 27 24
rect 31 20 33 24
rect 25 18 33 20
rect 35 23 43 25
rect 35 19 37 23
rect 41 19 43 23
rect 35 18 43 19
rect 45 19 54 25
rect 45 18 48 19
rect 4 8 11 18
rect 47 15 48 18
rect 52 15 54 19
rect 47 14 54 15
rect 56 14 61 25
rect 63 24 70 25
rect 63 20 65 24
rect 69 20 70 24
rect 63 19 70 20
rect 63 14 68 19
rect 4 4 6 8
rect 10 4 11 8
rect 4 3 11 4
<< pdiffusion >>
rect 39 68 45 69
rect 39 64 40 68
rect 44 64 45 68
rect 61 68 68 69
rect 39 63 45 64
rect 2 62 11 63
rect 2 58 3 62
rect 7 58 11 62
rect 2 55 11 58
rect 2 51 3 55
rect 7 51 11 55
rect 2 47 11 51
rect 13 47 18 63
rect 20 52 28 63
rect 20 48 22 52
rect 26 48 28 52
rect 20 47 28 48
rect 30 47 35 63
rect 37 62 45 63
rect 61 64 62 68
rect 66 64 68 68
rect 61 62 68 64
rect 37 49 47 62
rect 49 59 57 62
rect 49 55 51 59
rect 55 55 57 59
rect 49 49 57 55
rect 59 49 68 62
rect 37 47 45 49
<< metal1 >>
rect -2 68 74 72
rect -2 64 40 68
rect 44 64 62 68
rect 66 64 74 68
rect 3 62 7 64
rect 3 55 7 58
rect 3 50 7 51
rect 10 55 51 59
rect 55 55 70 59
rect 10 43 14 55
rect 3 39 4 43
rect 8 39 14 43
rect 10 33 14 35
rect 18 33 22 52
rect 26 48 27 52
rect 33 46 63 50
rect 33 43 38 46
rect 59 45 63 46
rect 26 42 38 43
rect 30 38 38 42
rect 26 37 38 38
rect 47 39 48 43
rect 52 42 53 43
rect 52 39 55 42
rect 59 40 63 41
rect 47 37 55 39
rect 51 34 55 37
rect 18 29 32 33
rect 41 29 42 33
rect 46 29 48 33
rect 51 30 63 34
rect 10 27 14 29
rect 2 21 14 27
rect 26 24 32 29
rect 44 26 48 29
rect 66 26 70 55
rect 44 24 70 26
rect 17 23 21 24
rect 2 13 6 21
rect 26 20 27 24
rect 31 20 32 24
rect 37 23 41 24
rect 17 17 21 19
rect 44 22 65 24
rect 64 20 65 22
rect 69 20 70 24
rect 37 17 41 19
rect 17 13 41 17
rect 47 15 48 19
rect 52 15 53 19
rect 47 8 53 15
rect -2 4 6 8
rect 10 4 26 8
rect 30 4 34 8
rect 38 4 74 8
rect -2 0 74 4
<< ntransistor >>
rect 13 18 15 25
rect 23 18 25 25
rect 33 18 35 25
rect 43 18 45 25
rect 54 14 56 25
rect 61 14 63 25
<< ptransistor >>
rect 11 47 13 63
rect 18 47 20 63
rect 28 47 30 63
rect 35 47 37 63
rect 47 49 49 62
rect 57 49 59 62
<< polycontact >>
rect 4 39 8 43
rect 26 38 30 42
rect 10 29 14 33
rect 48 39 52 43
rect 59 41 63 45
rect 42 29 46 33
<< ndcontact >>
rect 17 19 21 23
rect 27 20 31 24
rect 37 19 41 23
rect 48 15 52 19
rect 65 20 69 24
rect 6 4 10 8
<< pdcontact >>
rect 40 64 44 68
rect 3 58 7 62
rect 3 51 7 55
rect 22 48 26 52
rect 62 64 66 68
rect 51 55 55 59
<< psubstratepcontact >>
rect 26 4 30 8
rect 34 4 38 8
<< psubstratepdiff >>
rect 25 8 39 9
rect 25 4 26 8
rect 30 4 34 8
rect 38 4 39 8
rect 25 3 39 4
<< labels >>
rlabel polycontact 6 41 6 41 6 b
rlabel metal1 4 20 4 20 6 a3
rlabel metal1 19 18 19 18 6 n4
rlabel metal1 12 28 12 28 6 a3
rlabel metal1 20 40 20 40 6 z
rlabel metal1 8 41 8 41 6 b
rlabel metal1 36 4 36 4 6 vss
rlabel metal1 39 18 39 18 6 n4
rlabel metal1 28 24 28 24 6 z
rlabel polycontact 28 40 28 40 6 b2
rlabel metal1 36 44 36 44 6 b2
rlabel metal1 36 68 36 68 6 vdd
rlabel metal1 52 40 52 40 6 b1
rlabel metal1 44 48 44 48 6 b2
rlabel metal1 52 48 52 48 6 b2
rlabel metal1 60 32 60 32 6 b1
rlabel metal1 60 48 60 48 6 b2
rlabel metal1 40 57 40 57 6 b
rlabel metal1 68 39 68 39 6 b
<< end >>
