magic
tech scmos
timestamp 1179385359
<< checkpaint >>
rect -22 -25 78 105
<< ab >>
rect 0 0 56 80
<< pwell >>
rect -4 -7 60 36
<< nwell >>
rect -4 36 60 87
<< polysilicon >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 39 70 41 74
rect 9 33 11 43
rect 19 40 21 43
rect 29 40 31 43
rect 19 39 25 40
rect 19 35 20 39
rect 24 35 25 39
rect 19 34 25 35
rect 29 39 35 40
rect 29 35 30 39
rect 34 35 35 39
rect 29 34 35 35
rect 39 39 41 43
rect 39 38 47 39
rect 39 34 42 38
rect 46 34 47 38
rect 9 32 15 33
rect 9 28 10 32
rect 14 28 15 32
rect 23 30 25 34
rect 31 30 33 34
rect 39 33 47 34
rect 39 30 41 33
rect 9 27 15 28
rect 13 24 15 27
rect 13 12 15 17
rect 23 9 25 14
rect 31 9 33 14
rect 39 9 41 14
<< ndiffusion >>
rect 18 24 23 30
rect 4 17 13 24
rect 15 22 23 24
rect 15 18 17 22
rect 21 18 23 22
rect 15 17 23 18
rect 4 12 11 17
rect 18 14 23 17
rect 25 14 31 30
rect 33 14 39 30
rect 41 19 48 30
rect 41 15 43 19
rect 47 15 48 19
rect 41 14 48 15
rect 4 8 6 12
rect 10 8 11 12
rect 4 7 11 8
<< pdiffusion >>
rect 4 64 9 70
rect 2 63 9 64
rect 2 59 3 63
rect 7 59 9 63
rect 2 55 9 59
rect 2 51 3 55
rect 7 51 9 55
rect 2 50 9 51
rect 4 43 9 50
rect 11 62 19 70
rect 11 58 13 62
rect 17 58 19 62
rect 11 55 19 58
rect 11 51 13 55
rect 17 51 19 55
rect 11 43 19 51
rect 21 69 29 70
rect 21 65 23 69
rect 27 65 29 69
rect 21 62 29 65
rect 21 58 23 62
rect 27 58 29 62
rect 21 43 29 58
rect 31 62 39 70
rect 31 58 33 62
rect 37 58 39 62
rect 31 55 39 58
rect 31 51 33 55
rect 37 51 39 55
rect 31 43 39 51
rect 41 69 48 70
rect 41 65 43 69
rect 47 65 48 69
rect 41 62 48 65
rect 41 58 43 62
rect 47 58 48 62
rect 41 43 48 58
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect -2 69 58 78
rect -2 68 23 69
rect 22 65 23 68
rect 27 68 43 69
rect 27 65 28 68
rect 2 59 3 63
rect 7 59 8 63
rect 2 55 8 59
rect 2 51 3 55
rect 7 51 8 55
rect 13 62 17 63
rect 22 62 28 65
rect 42 65 43 68
rect 47 68 58 69
rect 47 65 48 68
rect 22 58 23 62
rect 27 58 28 62
rect 33 62 37 63
rect 42 62 48 65
rect 42 58 43 62
rect 47 58 48 62
rect 13 55 17 58
rect 33 55 37 58
rect 17 51 33 54
rect 2 22 6 51
rect 13 50 37 51
rect 10 41 24 47
rect 41 46 47 54
rect 17 39 24 41
rect 17 35 20 39
rect 29 42 47 46
rect 29 39 35 42
rect 29 35 30 39
rect 34 35 35 39
rect 17 34 24 35
rect 41 34 42 38
rect 46 34 47 38
rect 10 32 14 33
rect 41 31 47 34
rect 14 28 30 30
rect 10 26 30 28
rect 2 18 17 22
rect 21 18 22 22
rect 2 17 22 18
rect 26 17 30 26
rect 34 25 47 31
rect 43 19 47 20
rect 43 12 47 15
rect -2 8 6 12
rect 10 8 58 12
rect -2 2 58 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
<< ntransistor >>
rect 13 17 15 24
rect 23 14 25 30
rect 31 14 33 30
rect 39 14 41 30
<< ptransistor >>
rect 9 43 11 70
rect 19 43 21 70
rect 29 43 31 70
rect 39 43 41 70
<< polycontact >>
rect 20 35 24 39
rect 30 35 34 39
rect 42 34 46 38
rect 10 28 14 32
<< ndcontact >>
rect 17 18 21 22
rect 43 15 47 19
rect 6 8 10 12
<< pdcontact >>
rect 3 59 7 63
rect 3 51 7 55
rect 13 58 17 62
rect 13 51 17 55
rect 23 65 27 69
rect 23 58 27 62
rect 33 58 37 62
rect 33 51 37 55
rect 43 65 47 69
rect 43 58 47 62
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
<< psubstratepdiff >>
rect 0 2 56 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 56 2
rect 0 -3 56 -2
<< nsubstratendiff >>
rect 0 82 56 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 56 82
rect 0 77 56 78
<< labels >>
rlabel metal1 4 40 4 40 6 z
rlabel metal1 12 20 12 20 6 z
rlabel metal1 12 44 12 44 6 a3
rlabel metal1 15 56 15 56 6 n3
rlabel metal1 28 6 28 6 6 vss
rlabel metal1 20 28 20 28 6 b
rlabel metal1 28 20 28 20 6 b
rlabel metal1 20 40 20 40 6 a3
rlabel metal1 28 74 28 74 6 vdd
rlabel metal1 36 28 36 28 6 a1
rlabel metal1 44 32 44 32 6 a1
rlabel metal1 36 44 36 44 6 a2
rlabel metal1 44 48 44 48 6 a2
rlabel metal1 35 56 35 56 6 n3
<< end >>
