.subckt mx3_x2 cmd0 cmd1 i0 i1 i2 q vdd vss
*   SPICE3 file   created from mx3_x2.ext -      technology: scmos
m00 w1     i2     w2     vdd p w=19u  l=2.3636u ad=95p      pd=29.7838u as=114.339p ps=38u
m01 w3     cmd1   w1     vdd p w=18u  l=2.3636u ad=124.364p pd=41.2364u as=90p      ps=28.2162u
m02 w4     cmd1   vdd    vdd p w=14u  l=2.3636u ad=112p     pd=44u      as=97.3204p ps=30.7184u
m03 w5     w4     w3     vdd p w=19u  l=2.3636u ad=57p      pd=25u      as=131.273p ps=43.5273u
m04 w2     i1     w5     vdd p w=19u  l=2.3636u ad=114.339p pd=38u      as=57p      ps=25u
m05 vdd    w6     w2     vdd p w=18u  l=2.3636u ad=125.126p pd=39.4951u as=108.321p ps=36u
m06 w7     cmd0   vdd    vdd p w=18u  l=2.3636u ad=54p      pd=24u      as=125.126p ps=39.4951u
m07 w3     i0     w7     vdd p w=18u  l=2.3636u ad=124.364p pd=41.2364u as=54p      ps=24u
m08 w4     cmd1   vss    vss n w=8u   l=2.3636u ad=64p      pd=32u      as=65.5172p ps=24.5517u
m09 vdd    cmd0   w6     vdd p w=14u  l=2.3636u ad=97.3204p pd=30.7184u as=112p     ps=44u
m10 q      w3     vdd    vdd p w=39u  l=2.3636u ad=312p     pd=94u      as=271.107p ps=85.5728u
m11 w8     i2     w9     vss n w=12u  l=2.3636u ad=60p      pd=22u      as=82p      ps=31.3333u
m12 w3     w4     w8     vss n w=12u  l=2.3636u ad=100p     pd=37.3333u as=60p      ps=22u
m13 w10    cmd1   w3     vss n w=12u  l=2.3636u ad=36p      pd=18u      as=100p     ps=37.3333u
m14 w9     i1     w10    vss n w=12u  l=2.3636u ad=82p      pd=31.3333u as=36p      ps=18u
m15 vss    cmd0   w6     vss n w=6u   l=2.3636u ad=49.1379p pd=18.4138u as=48p      ps=28u
m16 vss    cmd0   w9     vss n w=12u  l=2.3636u ad=98.2759p pd=36.8276u as=82p      ps=31.3333u
m17 w11    w6     vss    vss n w=12u  l=2.3636u ad=36p      pd=18u      as=98.2759p ps=36.8276u
m18 w3     i0     w11    vss n w=12u  l=2.3636u ad=100p     pd=37.3333u as=36p      ps=18u
m19 q      w3     vss    vss n w=20u  l=2.3636u ad=160p     pd=56u      as=163.793p ps=61.3793u
C0  q      w3     0.275f
C1  w2     w4     0.070f
C2  i0     cmd0   0.348f
C3  vdd    w6     0.013f
C4  w3     i1     0.078f
C5  w11    vss    0.010f
C6  w8     w9     0.019f
C7  q      i0     0.027f
C8  w5     w2     0.012f
C9  w9     cmd0   0.002f
C10 i0     i1     0.029f
C11 cmd0   w6     0.316f
C12 vdd    w4     0.046f
C13 w3     cmd1   0.047f
C14 w2     i2     0.010f
C15 w8     vss    0.007f
C16 vss    cmd0   0.017f
C17 w5     vdd    0.011f
C18 q      w6     0.059f
C19 w9     i1     0.022f
C20 w6     i1     0.130f
C21 i0     cmd1   0.008f
C22 vdd    i2     0.008f
C23 cmd0   w4     0.026f
C24 q      vss    0.050f
C25 w2     vdd    0.304f
C26 vss    i1     0.015f
C27 w9     cmd1   0.005f
C28 w6     cmd1   0.045f
C29 cmd0   i2     0.012f
C30 i1     w4     0.177f
C31 w2     cmd0   0.002f
C32 w3     i0     0.186f
C33 vss    cmd1   0.055f
C34 i1     i2     0.057f
C35 w4     cmd1   0.391f
C36 w9     w3     0.108f
C37 vdd    cmd0   0.017f
C38 w3     w6     0.334f
C39 w2     i1     0.022f
C40 w10    w9     0.012f
C41 cmd1   i2     0.184f
C42 vss    w3     0.182f
C43 q      vdd    0.067f
C44 w2     cmd1   0.106f
C45 w3     w4     0.146f
C46 i0     w6     0.309f
C47 vdd    i1     0.017f
C48 w10    vss    0.004f
C49 w1     w2     0.019f
C50 q      cmd0   0.003f
C51 w7     vdd    0.011f
C52 w9     w6     0.020f
C53 vss    i0     0.022f
C54 cmd0   i1     0.078f
C55 i0     w4     0.015f
C56 vdd    cmd1   0.123f
C57 w3     i2     0.014f
C58 w9     vss    0.293f
C59 w9     w4     0.131f
C60 w2     w3     0.159f
C61 w1     vdd    0.019f
C62 vss    w6     0.075f
C63 cmd0   cmd1   0.030f
C64 w6     w4     0.038f
C65 w3     vdd    0.223f
C66 vss    w4     0.043f
C67 w9     i2     0.012f
C68 i1     cmd1   0.151f
C69 w6     i2     0.022f
C70 w3     cmd0   0.261f
C71 vdd    i0     0.023f
C72 vss    i2     0.008f
C73 w4     i2     0.165f
C74 q      vss    0.013f
C76 w3     vss    0.067f
C78 i0     vss    0.049f
C79 cmd0   vss    0.067f
C80 w6     vss    0.057f
C81 i1     vss    0.038f
C82 w4     vss    0.049f
C83 cmd1   vss    0.071f
C84 i2     vss    0.032f
.ends
