magic
tech scmos
timestamp 1179387754
<< checkpaint >>
rect -22 -25 94 105
<< ab >>
rect 0 0 72 80
<< pwell >>
rect -4 -7 76 36
<< nwell >>
rect -4 36 76 87
<< polysilicon >>
rect 20 69 22 74
rect 30 69 32 74
rect 40 69 42 74
rect 50 69 52 74
rect 2 61 8 62
rect 2 57 3 61
rect 7 58 8 61
rect 7 57 11 58
rect 2 56 11 57
rect 9 53 11 56
rect 61 55 63 60
rect 9 39 11 42
rect 20 39 22 42
rect 30 39 32 42
rect 9 37 22 39
rect 26 38 32 39
rect 9 28 11 37
rect 26 34 27 38
rect 31 34 32 38
rect 26 33 32 34
rect 40 39 42 42
rect 50 39 52 42
rect 61 39 63 44
rect 40 38 46 39
rect 40 34 41 38
rect 45 34 46 38
rect 40 33 46 34
rect 50 38 70 39
rect 50 37 65 38
rect 19 31 28 33
rect 19 28 21 31
rect 40 30 42 33
rect 50 30 52 37
rect 61 34 65 37
rect 69 34 70 38
rect 61 33 70 34
rect 61 30 63 33
rect 9 8 11 22
rect 29 23 31 27
rect 19 12 21 16
rect 61 19 63 24
rect 40 13 42 18
rect 50 13 52 18
rect 29 8 31 11
rect 9 6 31 8
<< ndiffusion >>
rect 33 29 40 30
rect 2 27 9 28
rect 2 23 3 27
rect 7 23 9 27
rect 2 22 9 23
rect 11 27 19 28
rect 11 23 13 27
rect 17 23 19 27
rect 11 22 19 23
rect 13 16 19 22
rect 21 23 26 28
rect 33 25 34 29
rect 38 25 40 29
rect 33 23 40 25
rect 21 21 29 23
rect 21 17 23 21
rect 27 17 29 21
rect 21 16 29 17
rect 24 11 29 16
rect 31 18 40 23
rect 42 23 50 30
rect 42 19 44 23
rect 48 19 50 23
rect 42 18 50 19
rect 52 24 61 30
rect 63 29 70 30
rect 63 25 65 29
rect 69 25 70 29
rect 63 24 70 25
rect 52 23 59 24
rect 52 19 54 23
rect 58 19 59 23
rect 52 18 59 19
rect 31 11 36 18
<< pdiffusion >>
rect 13 66 20 69
rect 13 62 14 66
rect 18 62 20 66
rect 13 53 20 62
rect 4 48 9 53
rect 2 47 9 48
rect 2 43 3 47
rect 7 43 9 47
rect 2 42 9 43
rect 11 42 20 53
rect 22 63 30 69
rect 22 59 24 63
rect 28 59 30 63
rect 22 42 30 59
rect 32 54 40 69
rect 32 50 34 54
rect 38 50 40 54
rect 32 47 40 50
rect 32 43 34 47
rect 38 43 40 47
rect 32 42 40 43
rect 42 63 50 69
rect 42 59 44 63
rect 48 59 50 63
rect 42 42 50 59
rect 52 62 59 69
rect 52 58 54 62
rect 58 58 59 62
rect 52 55 59 58
rect 52 44 61 55
rect 63 54 70 55
rect 63 50 65 54
rect 69 50 70 54
rect 63 49 70 50
rect 63 44 68 49
rect 52 42 59 44
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect -2 68 74 78
rect 13 66 19 68
rect 2 61 7 63
rect 13 62 14 66
rect 18 62 19 66
rect 2 57 3 61
rect 23 59 24 63
rect 28 59 44 63
rect 48 59 49 63
rect 53 62 59 68
rect 53 58 54 62
rect 58 58 59 62
rect 7 57 14 58
rect 2 54 14 57
rect 10 49 14 54
rect 26 54 38 55
rect 26 50 34 54
rect 26 49 38 50
rect 3 47 7 48
rect 3 37 7 43
rect 34 47 38 49
rect 27 38 31 39
rect 3 34 27 37
rect 3 33 31 34
rect 3 27 7 33
rect 34 29 38 43
rect 50 50 65 54
rect 69 50 70 54
rect 50 39 54 50
rect 57 42 70 46
rect 41 38 54 39
rect 45 34 54 38
rect 41 33 54 34
rect 65 38 70 42
rect 69 34 70 38
rect 65 33 70 34
rect 3 22 7 23
rect 13 27 17 28
rect 50 30 54 33
rect 50 29 70 30
rect 50 26 65 29
rect 64 25 65 26
rect 69 25 70 29
rect 34 24 38 25
rect 13 12 17 23
rect 43 21 44 23
rect 22 17 23 21
rect 27 19 44 21
rect 48 19 49 23
rect 27 17 49 19
rect 53 19 54 23
rect 58 19 59 23
rect 53 12 59 19
rect -2 2 74 12
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
<< ntransistor >>
rect 9 22 11 28
rect 19 16 21 28
rect 29 11 31 23
rect 40 18 42 30
rect 50 18 52 30
rect 61 24 63 30
<< ptransistor >>
rect 9 42 11 53
rect 20 42 22 69
rect 30 42 32 69
rect 40 42 42 69
rect 50 42 52 69
rect 61 44 63 55
<< polycontact >>
rect 3 57 7 61
rect 27 34 31 38
rect 41 34 45 38
rect 65 34 69 38
<< ndcontact >>
rect 3 23 7 27
rect 13 23 17 27
rect 34 25 38 29
rect 23 17 27 21
rect 44 19 48 23
rect 65 25 69 29
rect 54 19 58 23
<< pdcontact >>
rect 14 62 18 66
rect 3 43 7 47
rect 24 59 28 63
rect 34 50 38 54
rect 34 43 38 47
rect 44 59 48 63
rect 54 58 58 62
rect 65 50 69 54
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
<< psubstratepdiff >>
rect 0 2 72 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 72 2
rect 0 -3 72 -2
<< nsubstratendiff >>
rect 0 82 72 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 72 82
rect 0 77 72 78
<< labels >>
rlabel polycontact 29 36 29 36 6 bn
rlabel polycontact 43 36 43 36 6 an
rlabel metal1 12 52 12 52 6 b
rlabel polycontact 4 60 4 60 6 b
rlabel metal1 17 35 17 35 6 bn
rlabel metal1 28 52 28 52 6 z
rlabel metal1 36 6 36 6 6 vss
rlabel metal1 35 19 35 19 6 n2
rlabel metal1 47 36 47 36 6 an
rlabel metal1 36 40 36 40 6 z
rlabel metal1 36 61 36 61 6 n1
rlabel metal1 36 74 36 74 6 vdd
rlabel ndcontact 67 27 67 27 6 an
rlabel polycontact 68 36 68 36 6 a
rlabel metal1 60 44 60 44 6 a
rlabel metal1 60 52 60 52 6 an
<< end >>
