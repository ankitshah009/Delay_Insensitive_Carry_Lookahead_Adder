magic
tech scmos
timestamp 1179385231
<< checkpaint >>
rect -22 -22 94 94
<< ab >>
rect 0 0 72 72
<< pwell >>
rect -4 -4 76 32
<< nwell >>
rect -4 32 76 76
<< polysilicon >>
rect 9 59 11 64
rect 21 59 23 64
rect 41 59 43 64
rect 51 59 53 64
rect 61 59 63 64
rect 9 44 11 47
rect 9 43 15 44
rect 9 39 10 43
rect 14 39 15 43
rect 9 38 15 39
rect 9 18 11 38
rect 21 34 23 47
rect 41 35 43 43
rect 51 35 53 43
rect 61 40 63 43
rect 60 39 70 40
rect 60 35 65 39
rect 69 35 70 39
rect 33 34 43 35
rect 16 33 24 34
rect 16 29 17 33
rect 21 29 24 33
rect 33 30 34 34
rect 38 31 43 34
rect 49 34 55 35
rect 38 30 45 31
rect 33 29 45 30
rect 49 30 50 34
rect 54 30 55 34
rect 49 29 55 30
rect 16 28 24 29
rect 22 25 24 28
rect 43 26 45 29
rect 53 26 55 29
rect 60 34 70 35
rect 60 26 62 34
rect 22 14 24 19
rect 9 7 11 12
rect 43 15 45 20
rect 53 14 55 19
rect 60 14 62 19
<< ndiffusion >>
rect 13 19 22 25
rect 24 24 31 25
rect 24 20 26 24
rect 30 20 31 24
rect 24 19 31 20
rect 35 20 43 26
rect 45 25 53 26
rect 45 21 47 25
rect 51 21 53 25
rect 45 20 53 21
rect 13 18 20 19
rect 2 17 9 18
rect 2 13 3 17
rect 7 13 9 17
rect 2 12 9 13
rect 11 12 20 18
rect 13 8 20 12
rect 13 4 14 8
rect 18 4 20 8
rect 13 3 20 4
rect 35 8 41 20
rect 48 19 53 20
rect 55 19 60 26
rect 62 24 69 26
rect 62 20 64 24
rect 68 20 69 24
rect 62 19 69 20
rect 35 4 36 8
rect 40 4 41 8
rect 35 3 41 4
<< pdiffusion >>
rect 13 68 19 69
rect 13 64 14 68
rect 18 64 19 68
rect 13 59 19 64
rect 4 53 9 59
rect 2 52 9 53
rect 2 48 3 52
rect 7 48 9 52
rect 2 47 9 48
rect 11 47 21 59
rect 23 53 28 59
rect 23 52 30 53
rect 23 48 25 52
rect 29 48 30 52
rect 36 49 41 59
rect 23 47 30 48
rect 34 48 41 49
rect 34 44 35 48
rect 39 44 41 48
rect 34 43 41 44
rect 43 58 51 59
rect 43 54 45 58
rect 49 54 51 58
rect 43 51 51 54
rect 43 47 45 51
rect 49 47 51 51
rect 43 43 51 47
rect 53 58 61 59
rect 53 54 55 58
rect 59 54 61 58
rect 53 43 61 54
rect 63 58 70 59
rect 63 54 65 58
rect 69 54 70 58
rect 63 51 70 54
rect 63 47 65 51
rect 69 47 70 51
rect 63 46 70 47
rect 63 43 68 46
<< metal1 >>
rect -2 68 74 72
rect -2 64 14 68
rect 18 64 30 68
rect 34 64 74 68
rect 10 53 22 59
rect 54 58 60 64
rect 44 54 45 58
rect 49 54 50 58
rect 54 54 55 58
rect 59 54 60 58
rect 64 54 65 58
rect 69 54 70 58
rect 2 52 7 53
rect 2 48 3 52
rect 2 47 7 48
rect 2 17 6 47
rect 10 43 14 53
rect 25 52 29 53
rect 10 37 14 39
rect 18 33 22 43
rect 10 29 17 33
rect 21 29 22 33
rect 25 34 29 48
rect 34 48 39 52
rect 34 44 35 48
rect 44 51 50 54
rect 64 51 70 54
rect 44 47 45 51
rect 49 47 65 51
rect 69 47 70 51
rect 34 43 39 44
rect 34 39 46 43
rect 25 30 34 34
rect 38 30 39 34
rect 10 21 14 29
rect 25 24 31 30
rect 25 20 26 24
rect 30 20 31 24
rect 42 25 46 39
rect 57 39 70 43
rect 57 38 65 39
rect 69 35 70 39
rect 49 30 50 34
rect 54 30 60 34
rect 42 21 47 25
rect 51 21 52 25
rect 56 17 60 30
rect 65 29 70 35
rect 2 13 3 17
rect 7 13 60 17
rect 64 24 68 25
rect 64 8 68 20
rect -2 4 14 8
rect 18 4 25 8
rect 29 4 36 8
rect 40 4 56 8
rect 60 4 64 8
rect 68 4 74 8
rect -2 0 74 4
<< ntransistor >>
rect 22 19 24 25
rect 43 20 45 26
rect 9 12 11 18
rect 53 19 55 26
rect 60 19 62 26
<< ptransistor >>
rect 9 47 11 59
rect 21 47 23 59
rect 41 43 43 59
rect 51 43 53 59
rect 61 43 63 59
<< polycontact >>
rect 10 39 14 43
rect 65 35 69 39
rect 17 29 21 33
rect 34 30 38 34
rect 50 30 54 34
<< ndcontact >>
rect 26 20 30 24
rect 47 21 51 25
rect 3 13 7 17
rect 14 4 18 8
rect 64 20 68 24
rect 36 4 40 8
<< pdcontact >>
rect 14 64 18 68
rect 3 48 7 52
rect 25 48 29 52
rect 35 44 39 48
rect 45 54 49 58
rect 45 47 49 51
rect 55 54 59 58
rect 65 54 69 58
rect 65 47 69 51
<< psubstratepcontact >>
rect 25 4 29 8
rect 56 4 60 8
rect 64 4 68 8
<< nsubstratencontact >>
rect 30 64 34 68
<< psubstratepdiff >>
rect 24 8 30 9
rect 24 4 25 8
rect 29 4 30 8
rect 24 3 30 4
rect 55 8 69 9
rect 55 4 56 8
rect 60 4 64 8
rect 68 4 69 8
rect 55 3 69 4
<< nsubstratendiff >>
rect 29 68 35 69
rect 29 64 30 68
rect 34 64 35 68
rect 29 63 35 64
<< labels >>
rlabel polysilicon 38 32 38 32 6 bn
rlabel polycontact 52 32 52 32 6 a2n
rlabel metal1 12 24 12 24 6 b
rlabel pdcontact 4 50 4 50 6 a2n
rlabel metal1 12 48 12 48 6 a2
rlabel metal1 27 36 27 36 6 bn
rlabel metal1 20 36 20 36 6 b
rlabel metal1 20 56 20 56 6 a2
rlabel metal1 36 4 36 4 6 vss
rlabel metal1 32 32 32 32 6 bn
rlabel metal1 44 32 44 32 6 z
rlabel metal1 36 48 36 48 6 z
rlabel metal1 47 52 47 52 6 n1
rlabel metal1 36 68 36 68 6 vdd
rlabel metal1 31 15 31 15 6 a2n
rlabel metal1 54 32 54 32 6 a2n
rlabel metal1 60 40 60 40 6 a1
rlabel polycontact 68 36 68 36 6 a1
rlabel metal1 57 49 57 49 6 n1
rlabel metal1 67 52 67 52 6 n1
<< end >>
