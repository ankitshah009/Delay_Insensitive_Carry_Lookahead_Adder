.subckt iv1v0x4 a vdd vss z
*   SPICE3 file   created from iv1v0x4.ext -      technology: scmos
m00 vdd    a      z      vdd p w=28u  l=2.3636u ad=176p     pd=50u      as=196p     ps=70u
m01 z      a      vdd    vdd p w=28u  l=2.3636u ad=196p     pd=70u      as=176p     ps=50u
m02 vss    a      z      vss n w=20u  l=2.3636u ad=136p     pd=42u      as=140p     ps=54u
m03 z      a      vss    vss n w=20u  l=2.3636u ad=140p     pd=54u      as=136p     ps=42u
C0  vss    z      0.182f
C1  z      a      0.329f
C2  a      vdd    0.246f
C3  vss    a      0.019f
C4  z      vdd    0.065f
C6  z      vss    0.002f
C7  a      vss    0.094f
.ends
