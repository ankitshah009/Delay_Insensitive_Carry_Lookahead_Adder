.subckt iv1v0x6 a vdd vss z
*   SPICE3 file   created from iv1v0x6.ext -      technology: scmos
m00 vdd    a      z      vdd p w=27u  l=2.3636u ad=135p     pd=46u      as=125.667p ps=46u
m01 z      a      vdd    vdd p w=27u  l=2.3636u ad=125.667p pd=46u      as=135p     ps=46u
m02 vdd    a      z      vdd p w=27u  l=2.3636u ad=135p     pd=46u      as=125.667p ps=46u
m03 z      a      vss    vss n w=20u  l=2.3636u ad=80p      pd=28u      as=143p     ps=55u
m04 vss    a      z      vss n w=20u  l=2.3636u ad=143p     pd=55u      as=80p      ps=28u
C0  vss    z      0.230f
C1  vdd    a      0.051f
C2  vss    vdd    0.009f
C3  vdd    z      0.083f
C4  vss    a      0.088f
C5  z      a      0.143f
C8  z      vss    0.006f
C9  a      vss    0.054f
.ends
