magic
tech scmos
timestamp 1180600701
<< checkpaint >>
rect -22 -22 92 122
<< ab >>
rect 0 0 70 100
<< pwell >>
rect -4 -4 74 48
<< nwell >>
rect -4 48 74 104
<< polysilicon >>
rect 23 94 25 98
rect 33 94 35 98
rect 45 94 47 98
rect 57 94 59 98
rect 11 85 13 89
rect 11 41 13 65
rect 23 53 25 56
rect 17 52 25 53
rect 17 48 18 52
rect 22 51 25 52
rect 22 48 23 51
rect 17 47 23 48
rect 33 43 35 55
rect 45 53 47 56
rect 57 53 59 56
rect 45 52 53 53
rect 45 51 48 52
rect 47 48 48 51
rect 52 48 53 52
rect 47 47 53 48
rect 57 52 63 53
rect 57 48 58 52
rect 62 48 63 52
rect 57 47 63 48
rect 27 42 35 43
rect 27 41 28 42
rect 11 39 28 41
rect 11 25 13 39
rect 27 38 28 39
rect 32 41 35 42
rect 32 39 47 41
rect 32 38 33 39
rect 27 37 33 38
rect 17 32 23 33
rect 17 28 18 32
rect 22 29 23 32
rect 29 32 35 33
rect 22 28 25 29
rect 17 27 25 28
rect 29 28 30 32
rect 34 28 35 32
rect 29 27 35 28
rect 23 24 25 27
rect 33 24 35 27
rect 45 25 47 39
rect 57 32 63 33
rect 57 28 58 32
rect 62 28 63 32
rect 57 27 63 28
rect 11 11 13 15
rect 57 24 59 27
rect 23 2 25 6
rect 33 2 35 6
rect 45 2 47 6
rect 57 2 59 6
<< ndiffusion >>
rect 3 22 11 25
rect 3 18 4 22
rect 8 18 11 22
rect 3 15 11 18
rect 13 24 18 25
rect 40 24 45 25
rect 13 15 23 24
rect 15 12 23 15
rect 15 8 16 12
rect 20 8 23 12
rect 15 6 23 8
rect 25 6 33 24
rect 35 22 45 24
rect 35 18 38 22
rect 42 18 45 22
rect 35 6 45 18
rect 47 24 52 25
rect 47 6 57 24
rect 59 12 67 24
rect 59 8 62 12
rect 66 8 67 12
rect 59 6 67 8
<< pdiffusion >>
rect 15 92 23 94
rect 15 88 16 92
rect 20 88 23 92
rect 15 85 23 88
rect 3 82 11 85
rect 3 78 4 82
rect 8 78 11 82
rect 3 72 11 78
rect 3 68 4 72
rect 8 68 11 72
rect 3 65 11 68
rect 13 65 23 85
rect 15 56 23 65
rect 25 56 33 94
rect 28 55 33 56
rect 35 72 45 94
rect 35 68 38 72
rect 42 68 45 72
rect 35 62 45 68
rect 35 58 38 62
rect 42 58 45 62
rect 35 56 45 58
rect 47 56 57 94
rect 59 92 67 94
rect 59 88 62 92
rect 66 88 67 92
rect 59 56 67 88
rect 35 55 40 56
<< metal1 >>
rect -2 92 72 100
rect -2 88 16 92
rect 20 88 62 92
rect 66 88 72 92
rect 4 82 8 83
rect 8 78 52 82
rect 4 72 8 78
rect 4 22 8 68
rect 18 52 22 73
rect 18 32 22 48
rect 28 42 32 73
rect 28 37 32 38
rect 38 72 42 73
rect 38 62 42 68
rect 38 42 42 58
rect 48 52 52 78
rect 48 47 52 48
rect 58 52 62 83
rect 38 37 44 42
rect 40 32 44 37
rect 58 32 62 48
rect 18 27 22 28
rect 29 28 30 32
rect 34 28 35 32
rect 40 28 53 32
rect 29 22 33 28
rect 40 22 44 28
rect 8 18 33 22
rect 37 18 38 22
rect 42 18 44 22
rect 4 17 8 18
rect 58 17 62 28
rect -2 8 16 12
rect 20 8 62 12
rect 66 8 72 12
rect -2 0 72 8
<< ntransistor >>
rect 11 15 13 25
rect 23 6 25 24
rect 33 6 35 24
rect 45 6 47 25
rect 57 6 59 24
<< ptransistor >>
rect 11 65 13 85
rect 23 56 25 94
rect 33 55 35 94
rect 45 56 47 94
rect 57 56 59 94
<< polycontact >>
rect 18 48 22 52
rect 48 48 52 52
rect 58 48 62 52
rect 28 38 32 42
rect 18 28 22 32
rect 30 28 34 32
rect 58 28 62 32
<< ndcontact >>
rect 4 18 8 22
rect 16 8 20 12
rect 38 18 42 22
rect 62 8 66 12
<< pdcontact >>
rect 16 88 20 92
rect 4 78 8 82
rect 4 68 8 72
rect 38 68 42 72
rect 38 58 42 62
rect 62 88 66 92
<< labels >>
rlabel polycontact 20 50 20 50 6 i0
rlabel metal1 30 55 30 55 6 cmd
rlabel metal1 35 6 35 6 6 vss
rlabel ndcontact 40 20 40 20 6 nq
rlabel metal1 50 30 50 30 6 nq
rlabel metal1 40 55 40 55 6 nq
rlabel metal1 35 94 35 94 6 vdd
rlabel polycontact 60 50 60 50 6 i1
<< end >>
