magic
tech scmos
timestamp 1179385339
<< checkpaint >>
rect -22 -25 78 105
<< ab >>
rect 0 0 56 80
<< pwell >>
rect -4 -7 60 36
<< nwell >>
rect -4 36 60 87
<< polysilicon >>
rect 9 66 11 71
rect 19 66 21 71
rect 29 66 31 71
rect 39 66 41 71
rect 9 47 11 50
rect 9 46 15 47
rect 9 42 10 46
rect 14 42 15 46
rect 9 41 15 42
rect 19 37 21 50
rect 29 44 31 50
rect 14 35 21 37
rect 25 42 31 44
rect 39 47 41 50
rect 39 46 47 47
rect 39 42 42 46
rect 46 42 47 46
rect 14 31 16 35
rect 25 31 27 42
rect 39 41 47 42
rect 39 37 41 41
rect 9 30 16 31
rect 9 26 10 30
rect 14 26 16 30
rect 9 25 16 26
rect 14 22 16 25
rect 21 30 27 31
rect 21 26 22 30
rect 26 26 27 30
rect 21 25 27 26
rect 31 35 41 37
rect 21 22 23 25
rect 31 22 33 35
rect 38 30 47 31
rect 38 26 42 30
rect 46 26 47 30
rect 38 25 47 26
rect 38 22 40 25
rect 14 10 16 15
rect 21 10 23 15
rect 31 10 33 15
rect 38 10 40 15
<< ndiffusion >>
rect 5 15 14 22
rect 16 15 21 22
rect 23 21 31 22
rect 23 17 25 21
rect 29 17 31 21
rect 23 15 31 17
rect 33 15 38 22
rect 40 20 48 22
rect 40 16 43 20
rect 47 16 48 20
rect 40 15 48 16
rect 5 12 12 15
rect 5 8 7 12
rect 11 8 12 12
rect 5 7 12 8
<< pdiffusion >>
rect 2 65 9 66
rect 2 61 3 65
rect 7 61 9 65
rect 2 50 9 61
rect 11 63 19 66
rect 11 59 13 63
rect 17 59 19 63
rect 11 50 19 59
rect 21 55 29 66
rect 21 51 23 55
rect 27 51 29 55
rect 21 50 29 51
rect 31 63 39 66
rect 31 59 33 63
rect 37 59 39 63
rect 31 50 39 59
rect 41 65 49 66
rect 41 61 43 65
rect 47 61 49 65
rect 41 50 49 61
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect -2 68 58 78
rect 3 65 7 68
rect 43 65 47 68
rect 3 60 7 61
rect 12 59 13 63
rect 17 59 33 63
rect 37 59 38 63
rect 43 60 47 61
rect 22 54 23 55
rect 2 51 23 54
rect 27 51 28 55
rect 2 50 28 51
rect 33 50 47 54
rect 2 21 6 50
rect 10 46 14 47
rect 41 46 47 50
rect 14 42 34 46
rect 41 42 42 46
rect 46 42 47 46
rect 10 41 34 42
rect 30 38 34 41
rect 10 34 23 38
rect 30 34 46 38
rect 10 30 14 34
rect 42 30 46 34
rect 21 26 22 30
rect 26 26 38 30
rect 10 25 14 26
rect 2 17 25 21
rect 29 17 30 21
rect 34 17 38 26
rect 42 25 46 26
rect 43 20 47 21
rect 43 12 47 16
rect -2 8 7 12
rect 11 8 58 12
rect -2 2 58 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
<< ntransistor >>
rect 14 15 16 22
rect 21 15 23 22
rect 31 15 33 22
rect 38 15 40 22
<< ptransistor >>
rect 9 50 11 66
rect 19 50 21 66
rect 29 50 31 66
rect 39 50 41 66
<< polycontact >>
rect 10 42 14 46
rect 42 42 46 46
rect 10 26 14 30
rect 22 26 26 30
rect 42 26 46 30
<< ndcontact >>
rect 25 17 29 21
rect 43 16 47 20
rect 7 8 11 12
<< pdcontact >>
rect 3 61 7 65
rect 13 59 17 63
rect 23 51 27 55
rect 33 59 37 63
rect 43 61 47 65
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
<< psubstratepdiff >>
rect 0 2 56 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 56 2
rect 0 -3 56 -2
<< nsubstratendiff >>
rect 0 82 56 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 56 82
rect 0 77 56 78
<< labels >>
rlabel metal1 4 32 4 32 6 z
rlabel polycontact 12 28 12 28 6 b1
rlabel metal1 12 52 12 52 6 z
rlabel metal1 28 6 28 6 6 vss
rlabel metal1 28 28 28 28 6 b2
rlabel metal1 20 36 20 36 6 b1
rlabel metal1 20 44 20 44 6 a1
rlabel metal1 28 44 28 44 6 a1
rlabel metal1 20 52 20 52 6 z
rlabel metal1 28 74 28 74 6 vdd
rlabel metal1 36 20 36 20 6 b2
rlabel polycontact 44 28 44 28 6 a1
rlabel metal1 36 36 36 36 6 a1
rlabel metal1 44 48 44 48 6 a2
rlabel metal1 36 52 36 52 6 a2
rlabel metal1 25 61 25 61 6 n3
<< end >>
