magic
tech scmos
timestamp 1179387674
<< checkpaint >>
rect -22 -25 262 105
<< ab >>
rect 0 0 240 80
<< pwell >>
rect -4 -7 244 36
<< nwell >>
rect -4 36 244 87
<< polysilicon >>
rect 9 69 11 74
rect 19 69 21 74
rect 29 69 31 74
rect 39 69 41 74
rect 49 69 51 74
rect 59 69 61 74
rect 79 72 91 74
rect 79 69 81 72
rect 89 69 91 72
rect 119 69 121 74
rect 129 69 131 74
rect 139 69 141 74
rect 149 69 151 74
rect 159 69 161 74
rect 169 69 171 74
rect 179 69 181 74
rect 189 69 191 74
rect 199 69 201 74
rect 209 69 211 74
rect 219 69 221 74
rect 99 56 101 61
rect 109 56 111 61
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 39 39 41 42
rect 49 39 51 42
rect 59 39 61 42
rect 9 38 61 39
rect 79 38 81 42
rect 89 39 91 42
rect 99 39 101 42
rect 109 39 111 42
rect 119 39 121 42
rect 129 39 131 42
rect 139 39 141 42
rect 149 39 151 42
rect 85 38 91 39
rect 9 34 10 38
rect 14 34 61 38
rect 9 33 61 34
rect 9 30 11 33
rect 19 30 21 33
rect 29 30 31 33
rect 59 30 61 33
rect 69 30 71 35
rect 85 34 86 38
rect 90 34 91 38
rect 79 30 81 34
rect 85 33 91 34
rect 95 38 115 39
rect 95 34 96 38
rect 100 34 110 38
rect 114 34 115 38
rect 95 33 115 34
rect 119 38 131 39
rect 119 34 123 38
rect 127 34 131 38
rect 119 33 131 34
rect 135 38 151 39
rect 135 34 136 38
rect 140 37 151 38
rect 140 34 141 37
rect 135 33 141 34
rect 159 35 161 42
rect 169 39 171 42
rect 169 38 175 39
rect 169 35 170 38
rect 159 34 170 35
rect 174 34 175 38
rect 159 33 175 34
rect 89 30 91 33
rect 96 30 98 33
rect 112 30 114 33
rect 119 30 121 33
rect 129 30 131 33
rect 136 30 138 33
rect 152 32 161 33
rect 9 7 11 12
rect 19 7 21 12
rect 29 7 31 12
rect 59 9 61 12
rect 69 9 71 12
rect 79 9 81 12
rect 152 28 153 32
rect 157 28 161 32
rect 172 30 174 33
rect 179 30 181 42
rect 189 39 191 42
rect 199 39 201 42
rect 209 39 211 42
rect 219 39 221 42
rect 189 38 231 39
rect 189 34 226 38
rect 230 34 231 38
rect 189 33 231 34
rect 189 30 191 33
rect 199 30 201 33
rect 209 30 211 33
rect 152 27 161 28
rect 59 7 81 9
rect 89 6 91 10
rect 96 6 98 10
rect 112 6 114 10
rect 119 6 121 10
rect 129 7 131 12
rect 136 8 138 12
rect 172 12 174 16
rect 179 8 181 16
rect 136 6 181 8
rect 189 7 191 12
rect 199 7 201 12
rect 209 7 211 12
<< ndiffusion >>
rect 2 25 9 30
rect 2 21 3 25
rect 7 21 9 25
rect 2 17 9 21
rect 2 13 3 17
rect 7 13 9 17
rect 2 12 9 13
rect 11 29 19 30
rect 11 25 13 29
rect 17 25 19 29
rect 11 22 19 25
rect 11 18 13 22
rect 17 18 19 22
rect 11 12 19 18
rect 21 17 29 30
rect 21 13 23 17
rect 27 13 29 17
rect 21 12 29 13
rect 31 29 38 30
rect 31 25 33 29
rect 37 25 38 29
rect 31 22 38 25
rect 31 18 33 22
rect 37 18 38 22
rect 31 17 38 18
rect 52 29 59 30
rect 52 25 53 29
rect 57 25 59 29
rect 52 22 59 25
rect 52 18 53 22
rect 57 18 59 22
rect 52 17 59 18
rect 31 12 36 17
rect 54 12 59 17
rect 61 22 69 30
rect 61 18 63 22
rect 67 18 69 22
rect 61 12 69 18
rect 71 29 79 30
rect 71 25 73 29
rect 77 25 79 29
rect 71 12 79 25
rect 81 22 89 30
rect 81 18 83 22
rect 87 18 89 22
rect 81 12 89 18
rect 84 10 89 12
rect 91 10 96 30
rect 98 15 112 30
rect 98 11 103 15
rect 107 11 112 15
rect 98 10 112 11
rect 114 10 119 30
rect 121 22 129 30
rect 121 18 123 22
rect 127 18 129 22
rect 121 12 129 18
rect 131 12 136 30
rect 138 15 147 30
rect 165 29 172 30
rect 165 25 166 29
rect 170 25 172 29
rect 165 24 172 25
rect 167 16 172 24
rect 174 16 179 30
rect 181 28 189 30
rect 181 24 183 28
rect 187 24 189 28
rect 181 21 189 24
rect 181 17 183 21
rect 187 17 189 21
rect 181 16 189 17
rect 138 12 141 15
rect 121 10 126 12
rect 140 11 141 12
rect 145 11 147 15
rect 140 10 147 11
rect 184 12 189 16
rect 191 29 199 30
rect 191 25 193 29
rect 197 25 199 29
rect 191 22 199 25
rect 191 18 193 22
rect 197 18 199 22
rect 191 12 199 18
rect 201 25 209 30
rect 201 21 203 25
rect 207 21 209 25
rect 201 17 209 21
rect 201 13 203 17
rect 207 13 209 17
rect 201 12 209 13
rect 211 29 218 30
rect 211 25 213 29
rect 217 25 218 29
rect 211 22 218 25
rect 211 18 213 22
rect 217 18 218 22
rect 211 17 218 18
rect 211 12 216 17
<< pdiffusion >>
rect 2 68 9 69
rect 2 64 3 68
rect 7 64 9 68
rect 2 61 9 64
rect 2 57 3 61
rect 7 57 9 61
rect 2 42 9 57
rect 11 54 19 69
rect 11 50 13 54
rect 17 50 19 54
rect 11 47 19 50
rect 11 43 13 47
rect 17 43 19 47
rect 11 42 19 43
rect 21 68 29 69
rect 21 64 23 68
rect 27 64 29 68
rect 21 61 29 64
rect 21 57 23 61
rect 27 57 29 61
rect 21 42 29 57
rect 31 54 39 69
rect 31 50 33 54
rect 37 50 39 54
rect 31 47 39 50
rect 31 43 33 47
rect 37 43 39 47
rect 31 42 39 43
rect 41 68 49 69
rect 41 64 43 68
rect 47 64 49 68
rect 41 61 49 64
rect 41 57 43 61
rect 47 57 49 61
rect 41 42 49 57
rect 51 54 59 69
rect 51 50 53 54
rect 57 50 59 54
rect 51 47 59 50
rect 51 43 53 47
rect 57 43 59 47
rect 51 42 59 43
rect 61 68 68 69
rect 61 64 63 68
rect 67 64 68 68
rect 61 61 68 64
rect 74 62 79 69
rect 61 57 63 61
rect 67 57 68 61
rect 61 42 68 57
rect 72 61 79 62
rect 72 57 73 61
rect 77 57 79 61
rect 72 54 79 57
rect 72 50 73 54
rect 77 50 79 54
rect 72 49 79 50
rect 74 42 79 49
rect 81 54 89 69
rect 81 50 83 54
rect 87 50 89 54
rect 81 47 89 50
rect 81 43 83 47
rect 87 43 89 47
rect 81 42 89 43
rect 91 56 96 69
rect 114 56 119 69
rect 91 55 99 56
rect 91 51 93 55
rect 97 51 99 55
rect 91 42 99 51
rect 101 47 109 56
rect 101 43 103 47
rect 107 43 109 47
rect 101 42 109 43
rect 111 55 119 56
rect 111 51 113 55
rect 117 51 119 55
rect 111 42 119 51
rect 121 47 129 69
rect 121 43 123 47
rect 127 43 129 47
rect 121 42 129 43
rect 131 62 139 69
rect 131 58 133 62
rect 137 58 139 62
rect 131 42 139 58
rect 141 47 149 69
rect 141 43 143 47
rect 147 43 149 47
rect 141 42 149 43
rect 151 62 159 69
rect 151 58 153 62
rect 157 58 159 62
rect 151 42 159 58
rect 161 54 169 69
rect 161 50 163 54
rect 167 50 169 54
rect 161 42 169 50
rect 171 61 179 69
rect 171 57 173 61
rect 177 57 179 61
rect 171 54 179 57
rect 171 50 173 54
rect 177 50 179 54
rect 171 47 179 50
rect 171 43 173 47
rect 177 43 179 47
rect 171 42 179 43
rect 181 54 189 69
rect 181 50 183 54
rect 187 50 189 54
rect 181 47 189 50
rect 181 43 183 47
rect 187 43 189 47
rect 181 42 189 43
rect 191 68 199 69
rect 191 64 193 68
rect 197 64 199 68
rect 191 61 199 64
rect 191 57 193 61
rect 197 57 199 61
rect 191 42 199 57
rect 201 54 209 69
rect 201 50 203 54
rect 207 50 209 54
rect 201 47 209 50
rect 201 43 203 47
rect 207 43 209 47
rect 201 42 209 43
rect 211 68 219 69
rect 211 64 213 68
rect 217 64 219 68
rect 211 61 219 64
rect 211 57 213 61
rect 217 57 219 61
rect 211 42 219 57
rect 221 55 226 69
rect 221 54 228 55
rect 221 50 223 54
rect 227 50 228 54
rect 221 47 228 50
rect 221 43 223 47
rect 227 43 228 47
rect 221 42 228 43
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect 118 78 122 82
rect 126 78 130 82
rect 134 78 138 82
rect 142 78 146 82
rect 150 78 154 82
rect 158 78 162 82
rect 166 78 170 82
rect 174 78 178 82
rect 182 78 186 82
rect 190 78 194 82
rect 198 78 202 82
rect 206 78 210 82
rect 214 78 218 82
rect 222 78 226 82
rect 230 78 234 82
rect 238 78 242 82
rect -2 68 242 78
rect 3 61 7 64
rect 3 56 7 57
rect 23 61 27 64
rect 23 56 27 57
rect 43 61 47 64
rect 43 56 47 57
rect 63 61 67 64
rect 63 56 67 57
rect 73 61 133 62
rect 77 58 133 61
rect 137 58 153 62
rect 157 61 177 62
rect 157 58 173 61
rect 77 57 78 58
rect 13 54 17 55
rect 13 47 17 50
rect 2 38 6 47
rect 33 54 37 55
rect 33 47 37 50
rect 17 43 33 46
rect 53 54 57 55
rect 53 47 57 50
rect 73 54 78 57
rect 92 55 98 58
rect 77 50 78 54
rect 73 49 78 50
rect 83 54 87 55
rect 92 51 93 55
rect 97 51 98 55
rect 112 55 118 58
rect 112 51 113 55
rect 117 51 118 55
rect 173 54 177 57
rect 193 61 197 64
rect 193 56 197 57
rect 213 61 217 64
rect 213 56 217 57
rect 37 43 53 46
rect 83 47 87 50
rect 134 50 163 54
rect 167 50 168 54
rect 57 43 83 46
rect 103 47 107 48
rect 134 47 138 50
rect 173 47 177 50
rect 87 43 100 46
rect 13 42 100 43
rect 2 34 10 38
rect 14 34 15 38
rect 2 33 15 34
rect 33 29 37 42
rect 86 38 90 39
rect 86 30 90 34
rect 96 38 100 42
rect 96 33 100 34
rect 103 30 107 43
rect 110 43 123 47
rect 127 43 138 47
rect 142 43 143 47
rect 147 43 149 47
rect 110 38 114 43
rect 134 38 138 43
rect 110 33 114 34
rect 122 34 123 38
rect 127 34 128 38
rect 134 34 136 38
rect 140 34 141 38
rect 122 30 128 34
rect 145 32 149 43
rect 162 43 173 46
rect 162 42 177 43
rect 183 54 187 55
rect 183 47 187 50
rect 203 54 207 55
rect 203 47 207 50
rect 223 54 228 55
rect 227 50 228 54
rect 223 47 228 50
rect 187 43 203 47
rect 207 43 223 47
rect 227 43 228 47
rect 145 30 153 32
rect 3 25 7 26
rect 3 17 7 21
rect 12 25 13 29
rect 17 25 33 29
rect 12 22 17 25
rect 12 18 13 22
rect 33 22 37 25
rect 12 17 17 18
rect 23 17 27 18
rect 33 17 37 18
rect 53 29 153 30
rect 57 26 73 29
rect 72 25 73 26
rect 77 28 153 29
rect 157 28 158 32
rect 77 26 149 28
rect 77 25 78 26
rect 53 22 57 25
rect 162 22 166 42
rect 183 38 187 43
rect 169 34 170 38
rect 174 34 187 38
rect 193 29 197 43
rect 170 25 171 29
rect 183 28 187 29
rect 62 18 63 22
rect 67 18 83 22
rect 87 18 123 22
rect 127 18 166 22
rect 183 21 187 24
rect 53 17 57 18
rect 213 29 217 43
rect 226 38 238 39
rect 230 34 238 38
rect 226 33 238 34
rect 193 22 197 25
rect 193 17 197 18
rect 203 25 207 26
rect 203 17 207 21
rect 234 25 238 33
rect 213 22 217 25
rect 213 17 217 18
rect 3 12 7 13
rect 23 12 27 13
rect 102 12 103 15
rect -2 11 103 12
rect 107 12 108 15
rect 140 12 141 15
rect 107 11 141 12
rect 145 12 146 15
rect 155 12 161 15
rect 183 12 187 17
rect 203 12 207 13
rect 145 11 242 12
rect -2 2 242 11
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 122 2
rect 126 -2 130 2
rect 134 -2 138 2
rect 142 -2 146 2
rect 150 -2 154 2
rect 158 -2 162 2
rect 166 -2 170 2
rect 174 -2 178 2
rect 182 -2 186 2
rect 190 -2 194 2
rect 198 -2 202 2
rect 206 -2 210 2
rect 214 -2 218 2
rect 222 -2 226 2
rect 230 -2 234 2
rect 238 -2 242 2
<< ntransistor >>
rect 9 12 11 30
rect 19 12 21 30
rect 29 12 31 30
rect 59 12 61 30
rect 69 12 71 30
rect 79 12 81 30
rect 89 10 91 30
rect 96 10 98 30
rect 112 10 114 30
rect 119 10 121 30
rect 129 12 131 30
rect 136 12 138 30
rect 172 16 174 30
rect 179 16 181 30
rect 189 12 191 30
rect 199 12 201 30
rect 209 12 211 30
<< ptransistor >>
rect 9 42 11 69
rect 19 42 21 69
rect 29 42 31 69
rect 39 42 41 69
rect 49 42 51 69
rect 59 42 61 69
rect 79 42 81 69
rect 89 42 91 69
rect 99 42 101 56
rect 109 42 111 56
rect 119 42 121 69
rect 129 42 131 69
rect 139 42 141 69
rect 149 42 151 69
rect 159 42 161 69
rect 169 42 171 69
rect 179 42 181 69
rect 189 42 191 69
rect 199 42 201 69
rect 209 42 211 69
rect 219 42 221 69
<< polycontact >>
rect 10 34 14 38
rect 86 34 90 38
rect 96 34 100 38
rect 110 34 114 38
rect 123 34 127 38
rect 136 34 140 38
rect 170 34 174 38
rect 153 28 157 32
rect 226 34 230 38
<< ndcontact >>
rect 3 21 7 25
rect 3 13 7 17
rect 13 25 17 29
rect 13 18 17 22
rect 23 13 27 17
rect 33 25 37 29
rect 33 18 37 22
rect 53 25 57 29
rect 53 18 57 22
rect 63 18 67 22
rect 73 25 77 29
rect 83 18 87 22
rect 103 11 107 15
rect 123 18 127 22
rect 166 25 170 29
rect 183 24 187 28
rect 183 17 187 21
rect 141 11 145 15
rect 193 25 197 29
rect 193 18 197 22
rect 203 21 207 25
rect 203 13 207 17
rect 213 25 217 29
rect 213 18 217 22
<< pdcontact >>
rect 3 64 7 68
rect 3 57 7 61
rect 13 50 17 54
rect 13 43 17 47
rect 23 64 27 68
rect 23 57 27 61
rect 33 50 37 54
rect 33 43 37 47
rect 43 64 47 68
rect 43 57 47 61
rect 53 50 57 54
rect 53 43 57 47
rect 63 64 67 68
rect 63 57 67 61
rect 73 57 77 61
rect 73 50 77 54
rect 83 50 87 54
rect 83 43 87 47
rect 93 51 97 55
rect 103 43 107 47
rect 113 51 117 55
rect 123 43 127 47
rect 133 58 137 62
rect 143 43 147 47
rect 153 58 157 62
rect 163 50 167 54
rect 173 57 177 61
rect 173 50 177 54
rect 173 43 177 47
rect 183 50 187 54
rect 183 43 187 47
rect 193 64 197 68
rect 193 57 197 61
rect 203 50 207 54
rect 203 43 207 47
rect 213 64 217 68
rect 213 57 217 61
rect 223 50 227 54
rect 223 43 227 47
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
rect 90 -2 94 2
rect 98 -2 102 2
rect 106 -2 110 2
rect 114 -2 118 2
rect 122 -2 126 2
rect 130 -2 134 2
rect 138 -2 142 2
rect 146 -2 150 2
rect 154 -2 158 2
rect 162 -2 166 2
rect 170 -2 174 2
rect 178 -2 182 2
rect 186 -2 190 2
rect 194 -2 198 2
rect 202 -2 206 2
rect 210 -2 214 2
rect 218 -2 222 2
rect 226 -2 230 2
rect 234 -2 238 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
rect 90 78 94 82
rect 98 78 102 82
rect 106 78 110 82
rect 114 78 118 82
rect 122 78 126 82
rect 130 78 134 82
rect 138 78 142 82
rect 146 78 150 82
rect 154 78 158 82
rect 162 78 166 82
rect 170 78 174 82
rect 178 78 182 82
rect 186 78 190 82
rect 194 78 198 82
rect 202 78 206 82
rect 210 78 214 82
rect 218 78 222 82
rect 226 78 230 82
rect 234 78 238 82
<< psubstratepdiff >>
rect 0 2 240 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 122 2
rect 126 -2 130 2
rect 134 -2 138 2
rect 142 -2 146 2
rect 150 -2 154 2
rect 158 -2 162 2
rect 166 -2 170 2
rect 174 -2 178 2
rect 182 -2 186 2
rect 190 -2 194 2
rect 198 -2 202 2
rect 206 -2 210 2
rect 214 -2 218 2
rect 222 -2 226 2
rect 230 -2 234 2
rect 238 -2 240 2
rect 0 -3 240 -2
<< nsubstratendiff >>
rect 0 82 240 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect 118 78 122 82
rect 126 78 130 82
rect 134 78 138 82
rect 142 78 146 82
rect 150 78 154 82
rect 158 78 162 82
rect 166 78 170 82
rect 174 78 178 82
rect 182 78 186 82
rect 190 78 194 82
rect 198 78 202 82
rect 206 78 210 82
rect 214 78 218 82
rect 222 78 226 82
rect 230 78 234 82
rect 238 78 240 82
rect 0 77 240 78
<< labels >>
rlabel polycontact 88 36 88 36 6 an
rlabel polysilicon 105 36 105 36 6 bn
rlabel polycontact 125 36 125 36 6 an
rlabel polycontact 138 36 138 36 6 bn
rlabel polycontact 156 30 156 30 6 an
rlabel polycontact 172 36 172 36 6 an
rlabel metal1 14 23 14 23 6 bn
rlabel polycontact 12 36 12 36 6 b
rlabel metal1 4 40 4 40 6 b
rlabel metal1 35 36 35 36 6 bn
rlabel metal1 15 48 15 48 6 bn
rlabel metal1 76 20 76 20 6 z
rlabel metal1 68 20 68 20 6 z
rlabel metal1 55 23 55 23 6 an
rlabel metal1 76 56 76 56 6 z
rlabel metal1 55 48 55 48 6 bn
rlabel metal1 100 20 100 20 6 z
rlabel metal1 108 20 108 20 6 z
rlabel metal1 116 20 116 20 6 z
rlabel metal1 92 20 92 20 6 z
rlabel ndcontact 84 20 84 20 6 z
rlabel metal1 88 32 88 32 6 an
rlabel metal1 98 39 98 39 6 bn
rlabel metal1 112 40 112 40 6 bn
rlabel metal1 105 37 105 37 6 an
rlabel metal1 85 48 85 48 6 bn
rlabel metal1 116 60 116 60 6 z
rlabel metal1 108 60 108 60 6 z
rlabel metal1 100 60 100 60 6 z
rlabel metal1 92 60 92 60 6 z
rlabel metal1 84 60 84 60 6 z
rlabel metal1 120 6 120 6 6 vss
rlabel ndcontact 124 20 124 20 6 z
rlabel metal1 156 20 156 20 6 z
rlabel metal1 148 20 148 20 6 z
rlabel metal1 132 20 132 20 6 z
rlabel metal1 140 20 140 20 6 z
rlabel metal1 151 30 151 30 6 an
rlabel metal1 125 32 125 32 6 an
rlabel metal1 101 28 101 28 6 an
rlabel metal1 136 44 136 44 6 bn
rlabel pdcontact 124 45 124 45 6 bn
rlabel pdcontact 145 45 145 45 6 an
rlabel metal1 124 60 124 60 6 z
rlabel pdcontact 156 60 156 60 6 z
rlabel metal1 148 60 148 60 6 z
rlabel metal1 140 60 140 60 6 z
rlabel metal1 132 60 132 60 6 z
rlabel metal1 120 74 120 74 6 vdd
rlabel metal1 164 32 164 32 6 z
rlabel metal1 178 36 178 36 6 an
rlabel metal1 172 44 172 44 6 z
rlabel metal1 195 32 195 32 6 an
rlabel metal1 151 52 151 52 6 bn
rlabel metal1 164 60 164 60 6 z
rlabel metal1 172 60 172 60 6 z
rlabel polycontact 228 36 228 36 6 a
rlabel metal1 236 32 236 32 6 a
rlabel metal1 215 32 215 32 6 an
rlabel pdcontact 205 45 205 45 6 an
rlabel metal1 225 49 225 49 6 an
rlabel metal1 205 49 205 49 6 an
<< end >>
