magic
tech scmos
timestamp 1179386383
<< checkpaint >>
rect -22 -25 110 105
<< ab >>
rect 0 0 88 80
<< pwell >>
rect -4 -7 92 36
<< nwell >>
rect -4 36 92 87
<< polysilicon >>
rect 9 66 11 71
rect 19 66 21 71
rect 29 66 31 71
rect 39 66 41 71
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 9 38 15 39
rect 9 34 10 38
rect 14 34 15 38
rect 9 33 15 34
rect 19 38 31 39
rect 19 34 26 38
rect 30 34 31 38
rect 39 39 41 42
rect 39 38 47 39
rect 39 35 42 38
rect 19 33 31 34
rect 12 30 14 33
rect 19 30 21 33
rect 29 30 31 33
rect 36 34 42 35
rect 46 35 47 38
rect 57 38 63 39
rect 57 35 58 38
rect 46 34 50 35
rect 36 33 50 34
rect 36 30 38 33
rect 48 30 50 33
rect 55 34 58 35
rect 62 35 63 38
rect 72 38 79 39
rect 62 34 67 35
rect 55 33 67 34
rect 55 30 57 33
rect 65 30 67 33
rect 72 34 74 38
rect 78 34 79 38
rect 72 33 79 34
rect 72 30 74 33
rect 12 6 14 10
rect 19 6 21 10
rect 29 6 31 10
rect 36 6 38 10
rect 48 6 50 10
rect 55 6 57 10
rect 65 6 67 10
rect 72 6 74 10
<< ndiffusion >>
rect 3 15 12 30
rect 3 11 5 15
rect 9 11 12 15
rect 3 10 12 11
rect 14 10 19 30
rect 21 22 29 30
rect 21 18 23 22
rect 27 18 29 22
rect 21 10 29 18
rect 31 10 36 30
rect 38 15 48 30
rect 38 11 41 15
rect 45 11 48 15
rect 38 10 48 11
rect 50 10 55 30
rect 57 22 65 30
rect 57 18 59 22
rect 63 18 65 22
rect 57 10 65 18
rect 67 10 72 30
rect 74 22 82 30
rect 74 18 76 22
rect 80 18 82 22
rect 74 15 82 18
rect 74 11 76 15
rect 80 11 82 15
rect 74 10 82 11
<< pdiffusion >>
rect 2 65 9 66
rect 2 61 3 65
rect 7 61 9 65
rect 2 42 9 61
rect 11 61 19 66
rect 11 57 13 61
rect 17 57 19 61
rect 11 54 19 57
rect 11 50 13 54
rect 17 50 19 54
rect 11 42 19 50
rect 21 65 29 66
rect 21 61 23 65
rect 27 61 29 65
rect 21 42 29 61
rect 31 62 39 66
rect 31 58 33 62
rect 37 58 39 62
rect 31 54 39 58
rect 31 50 33 54
rect 37 50 39 54
rect 31 42 39 50
rect 41 65 49 66
rect 41 61 43 65
rect 47 61 49 65
rect 41 57 49 61
rect 41 53 43 57
rect 47 53 49 57
rect 41 42 49 53
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect -2 68 90 78
rect 3 65 7 68
rect 23 65 27 68
rect 3 60 7 61
rect 13 61 17 62
rect 43 65 47 68
rect 23 60 27 61
rect 33 62 38 63
rect 13 54 17 57
rect 37 58 38 62
rect 33 54 38 58
rect 2 50 13 54
rect 17 50 33 54
rect 37 50 38 54
rect 43 57 47 61
rect 43 52 47 53
rect 2 22 6 50
rect 25 42 63 46
rect 10 38 14 39
rect 25 38 31 42
rect 57 38 63 42
rect 25 34 26 38
rect 30 34 31 38
rect 41 34 42 38
rect 46 34 47 38
rect 57 34 58 38
rect 62 34 63 38
rect 73 34 74 38
rect 78 34 79 38
rect 10 30 14 34
rect 41 30 47 34
rect 73 30 79 34
rect 10 26 79 30
rect 2 18 23 22
rect 27 18 59 22
rect 63 18 64 22
rect 75 18 76 22
rect 80 18 81 22
rect 75 15 81 18
rect 4 12 5 15
rect -2 11 5 12
rect 9 12 10 15
rect 40 12 41 15
rect 9 11 41 12
rect 45 12 46 15
rect 75 12 76 15
rect 45 11 76 12
rect 80 12 81 15
rect 80 11 90 12
rect -2 2 90 11
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
<< ntransistor >>
rect 12 10 14 30
rect 19 10 21 30
rect 29 10 31 30
rect 36 10 38 30
rect 48 10 50 30
rect 55 10 57 30
rect 65 10 67 30
rect 72 10 74 30
<< ptransistor >>
rect 9 42 11 66
rect 19 42 21 66
rect 29 42 31 66
rect 39 42 41 66
<< polycontact >>
rect 10 34 14 38
rect 26 34 30 38
rect 42 34 46 38
rect 58 34 62 38
rect 74 34 78 38
<< ndcontact >>
rect 5 11 9 15
rect 23 18 27 22
rect 41 11 45 15
rect 59 18 63 22
rect 76 18 80 22
rect 76 11 80 15
<< pdcontact >>
rect 3 61 7 65
rect 13 57 17 61
rect 13 50 17 54
rect 23 61 27 65
rect 33 58 37 62
rect 33 50 37 54
rect 43 61 47 65
rect 43 53 47 57
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
<< psubstratepdiff >>
rect 0 2 88 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 88 2
rect 0 -3 88 -2
<< nsubstratendiff >>
rect 0 82 88 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 88 82
rect 0 77 88 78
<< labels >>
rlabel metal1 12 20 12 20 6 z
rlabel polycontact 12 36 12 36 6 a
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 52 12 52 6 z
rlabel metal1 20 20 20 20 6 z
rlabel metal1 20 28 20 28 6 a
rlabel metal1 28 20 28 20 6 z
rlabel metal1 28 28 28 28 6 a
rlabel polycontact 28 36 28 36 6 b
rlabel metal1 28 40 28 40 6 b
rlabel metal1 20 52 20 52 6 z
rlabel metal1 28 52 28 52 6 z
rlabel metal1 44 6 44 6 6 vss
rlabel metal1 36 20 36 20 6 z
rlabel metal1 36 28 36 28 6 a
rlabel metal1 44 20 44 20 6 z
rlabel metal1 44 32 44 32 6 a
rlabel metal1 36 44 36 44 6 b
rlabel metal1 44 44 44 44 6 b
rlabel pdcontact 36 60 36 60 6 z
rlabel metal1 44 74 44 74 6 vdd
rlabel metal1 52 20 52 20 6 z
rlabel metal1 52 28 52 28 6 a
rlabel ndcontact 60 20 60 20 6 z
rlabel metal1 60 28 60 28 6 a
rlabel metal1 68 28 68 28 6 a
rlabel metal1 52 44 52 44 6 b
rlabel polycontact 60 36 60 36 6 b
rlabel metal1 60 40 60 40 6 b
rlabel metal1 76 32 76 32 6 a
<< end >>
