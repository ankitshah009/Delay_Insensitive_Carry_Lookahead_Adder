magic
tech scmos
timestamp 1180639944
<< checkpaint >>
rect -24 -26 94 126
<< ab >>
rect 0 0 70 100
<< pwell >>
rect -4 -6 74 49
<< nwell >>
rect -4 49 74 106
<< polysilicon >>
rect 11 83 13 88
rect 23 83 25 88
rect 35 83 37 88
rect 47 83 49 88
rect 59 83 61 87
rect 23 63 25 67
rect 11 45 13 63
rect 23 62 31 63
rect 23 58 26 62
rect 30 58 31 62
rect 23 57 31 58
rect 11 44 23 45
rect 11 43 18 44
rect 15 40 18 43
rect 22 40 23 44
rect 15 39 23 40
rect 15 36 17 39
rect 29 36 31 57
rect 35 52 37 67
rect 47 63 49 67
rect 47 62 53 63
rect 47 58 48 62
rect 52 58 53 62
rect 47 57 53 58
rect 35 51 43 52
rect 35 47 38 51
rect 42 47 43 51
rect 35 46 43 47
rect 37 36 39 46
rect 47 42 49 57
rect 59 53 61 67
rect 45 39 49 42
rect 57 52 63 53
rect 57 48 58 52
rect 62 48 63 52
rect 57 47 63 48
rect 57 41 59 47
rect 53 39 59 41
rect 45 36 47 39
rect 53 36 55 39
rect 15 21 17 26
rect 29 12 31 17
rect 37 12 39 17
rect 45 12 47 17
rect 53 12 55 17
<< ndiffusion >>
rect 7 35 15 36
rect 7 31 8 35
rect 12 31 15 35
rect 7 30 15 31
rect 10 26 15 30
rect 17 26 29 36
rect 19 22 29 26
rect 19 18 21 22
rect 25 18 29 22
rect 19 17 29 18
rect 31 17 37 36
rect 39 17 45 36
rect 47 17 53 36
rect 55 31 60 36
rect 55 30 63 31
rect 55 26 58 30
rect 62 26 63 30
rect 55 22 63 26
rect 55 18 58 22
rect 62 18 63 22
rect 55 17 63 18
<< pdiffusion >>
rect 15 92 21 93
rect 15 88 16 92
rect 20 88 21 92
rect 61 94 67 95
rect 39 92 45 93
rect 39 88 40 92
rect 44 88 45 92
rect 61 90 62 94
rect 66 90 67 94
rect 61 89 67 90
rect 15 83 21 88
rect 39 83 45 88
rect 63 83 67 89
rect 6 77 11 83
rect 3 76 11 77
rect 3 72 4 76
rect 8 72 11 76
rect 3 68 11 72
rect 3 64 4 68
rect 8 64 11 68
rect 3 63 11 64
rect 13 67 23 83
rect 25 82 35 83
rect 25 78 28 82
rect 32 78 35 82
rect 25 67 35 78
rect 37 67 47 83
rect 49 82 59 83
rect 49 78 52 82
rect 56 78 59 82
rect 49 67 59 78
rect 61 67 67 83
rect 13 63 21 67
<< metal1 >>
rect -2 94 72 100
rect -2 92 62 94
rect -2 88 16 92
rect 20 88 40 92
rect 44 90 62 92
rect 66 90 72 94
rect 44 88 72 90
rect 3 72 4 76
rect 3 64 4 68
rect 8 35 12 83
rect 18 78 28 82
rect 32 78 52 82
rect 56 78 57 82
rect 18 44 22 78
rect 28 68 43 73
rect 47 68 62 73
rect 28 63 32 68
rect 26 62 32 63
rect 30 58 32 62
rect 37 62 52 63
rect 37 58 48 62
rect 26 57 32 58
rect 28 47 32 57
rect 38 51 42 54
rect 22 40 33 43
rect 18 39 33 40
rect 12 31 22 33
rect 8 27 22 31
rect 21 22 25 23
rect 29 22 33 39
rect 38 32 42 47
rect 48 37 52 58
rect 58 52 62 68
rect 58 47 62 48
rect 38 27 53 32
rect 57 26 58 30
rect 62 26 63 30
rect 57 22 63 26
rect 29 18 58 22
rect 62 18 63 22
rect 21 12 25 18
rect -2 0 72 12
<< ntransistor >>
rect 15 26 17 36
rect 29 17 31 36
rect 37 17 39 36
rect 45 17 47 36
rect 53 17 55 36
<< ptransistor >>
rect 11 63 13 83
rect 23 67 25 83
rect 35 67 37 83
rect 47 67 49 83
rect 59 67 61 83
<< polycontact >>
rect 26 58 30 62
rect 18 40 22 44
rect 48 58 52 62
rect 38 47 42 51
rect 58 48 62 52
<< ndcontact >>
rect 8 31 12 35
rect 21 18 25 22
rect 58 26 62 30
rect 58 18 62 22
<< pdcontact >>
rect 16 88 20 92
rect 40 88 44 92
rect 62 90 66 94
rect 4 72 8 76
rect 4 64 8 68
rect 28 78 32 82
rect 52 78 56 82
<< psubstratepcontact >>
rect 8 4 12 8
rect 18 4 22 8
<< nsubstratencontact >>
rect 28 92 32 96
<< psubstratepdiff >>
rect 7 8 23 9
rect 7 4 8 8
rect 12 4 18 8
rect 22 4 23 8
rect 7 3 23 4
<< nsubstratendiff >>
rect 27 96 33 97
rect 27 92 28 96
rect 32 92 33 96
rect 27 91 33 92
<< labels >>
rlabel polycontact 19 42 19 42 6 zn
rlabel metal1 20 30 20 30 6 z
rlabel metal1 20 30 20 30 6 z
rlabel metal1 10 55 10 55 6 z
rlabel metal1 10 55 10 55 6 z
rlabel metal1 20 60 20 60 6 zn
rlabel metal1 35 6 35 6 6 vss
rlabel metal1 35 6 35 6 6 vss
rlabel metal1 30 60 30 60 6 a
rlabel metal1 30 60 30 60 6 a
rlabel metal1 35 94 35 94 6 vdd
rlabel metal1 35 94 35 94 6 vdd
rlabel metal1 50 30 50 30 6 b
rlabel metal1 50 30 50 30 6 b
rlabel metal1 40 40 40 40 6 b
rlabel metal1 40 40 40 40 6 b
rlabel metal1 50 50 50 50 6 c
rlabel metal1 50 50 50 50 6 c
rlabel metal1 40 60 40 60 6 c
rlabel metal1 40 60 40 60 6 c
rlabel metal1 40 70 40 70 6 a
rlabel metal1 40 70 40 70 6 a
rlabel metal1 50 70 50 70 6 d
rlabel metal1 50 70 50 70 6 d
rlabel metal1 60 24 60 24 6 zn
rlabel metal1 46 20 46 20 6 zn
rlabel metal1 60 60 60 60 6 d
rlabel metal1 60 60 60 60 6 d
rlabel metal1 37 80 37 80 6 zn
<< end >>
