magic
tech scmos
timestamp 1179385125
<< checkpaint >>
rect -22 -25 86 105
<< ab >>
rect 0 0 64 80
<< pwell >>
rect -4 -7 68 36
<< nwell >>
rect -4 36 68 87
<< polysilicon >>
rect 20 66 22 71
rect 30 66 32 71
rect 42 66 44 71
rect 52 66 54 71
rect 9 60 11 65
rect 9 39 11 48
rect 20 39 22 56
rect 30 53 32 56
rect 30 52 38 53
rect 30 48 33 52
rect 37 48 38 52
rect 30 47 38 48
rect 42 47 44 56
rect 9 38 16 39
rect 9 34 11 38
rect 15 34 16 38
rect 9 33 16 34
rect 20 38 28 39
rect 20 34 23 38
rect 27 34 28 38
rect 20 33 28 34
rect 9 28 11 33
rect 25 30 27 33
rect 32 30 34 47
rect 42 46 48 47
rect 42 43 43 46
rect 39 42 43 43
rect 47 42 48 46
rect 39 41 48 42
rect 39 30 41 41
rect 52 39 54 56
rect 52 38 58 39
rect 52 35 53 38
rect 46 34 53 35
rect 57 34 58 38
rect 46 33 58 34
rect 46 30 48 33
rect 9 17 11 22
rect 25 13 27 18
rect 32 13 34 18
rect 39 13 41 18
rect 46 13 48 18
<< ndiffusion >>
rect 13 28 25 30
rect 2 27 9 28
rect 2 23 3 27
rect 7 23 9 27
rect 2 22 9 23
rect 11 22 25 28
rect 13 18 25 22
rect 27 18 32 30
rect 34 18 39 30
rect 41 18 46 30
rect 48 24 53 30
rect 48 23 55 24
rect 48 19 50 23
rect 54 19 55 23
rect 48 18 55 19
rect 13 12 23 18
rect 13 8 16 12
rect 20 8 23 12
rect 13 7 23 8
<< pdiffusion >>
rect 34 72 40 73
rect 34 68 35 72
rect 39 68 40 72
rect 34 66 40 68
rect 13 63 20 66
rect 13 60 14 63
rect 4 54 9 60
rect 2 53 9 54
rect 2 49 3 53
rect 7 49 9 53
rect 2 48 9 49
rect 11 59 14 60
rect 18 59 20 63
rect 11 56 20 59
rect 22 63 30 66
rect 22 59 24 63
rect 28 59 30 63
rect 22 56 30 59
rect 32 56 42 66
rect 44 63 52 66
rect 44 59 46 63
rect 50 59 52 63
rect 44 56 52 59
rect 54 65 61 66
rect 54 61 56 65
rect 60 61 61 65
rect 54 56 61 61
rect 11 48 18 56
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect -2 72 66 78
rect -2 68 35 72
rect 39 68 66 72
rect 14 63 18 68
rect 56 65 60 68
rect 2 53 7 63
rect 14 58 18 59
rect 23 59 24 63
rect 28 59 46 63
rect 50 59 51 63
rect 56 60 60 61
rect 23 54 27 59
rect 2 49 3 53
rect 2 48 7 49
rect 14 50 27 54
rect 33 52 47 54
rect 2 28 6 48
rect 14 38 18 50
rect 37 50 47 52
rect 33 46 37 48
rect 58 46 62 55
rect 25 42 37 46
rect 41 42 43 46
rect 47 42 62 46
rect 10 34 11 38
rect 15 34 18 38
rect 22 34 23 38
rect 27 34 31 38
rect 41 34 53 38
rect 57 34 62 38
rect 14 31 18 34
rect 2 27 7 28
rect 14 27 22 31
rect 2 23 3 27
rect 2 17 14 23
rect 18 21 22 27
rect 26 30 31 34
rect 26 26 39 30
rect 50 23 54 24
rect 18 19 50 21
rect 18 17 54 19
rect 58 17 62 34
rect -2 8 16 12
rect 20 8 66 12
rect -2 2 66 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
<< ntransistor >>
rect 9 22 11 28
rect 25 18 27 30
rect 32 18 34 30
rect 39 18 41 30
rect 46 18 48 30
<< ptransistor >>
rect 9 48 11 60
rect 20 56 22 66
rect 30 56 32 66
rect 42 56 44 66
rect 52 56 54 66
<< polycontact >>
rect 33 48 37 52
rect 11 34 15 38
rect 23 34 27 38
rect 43 42 47 46
rect 53 34 57 38
<< ndcontact >>
rect 3 23 7 27
rect 50 19 54 23
rect 16 8 20 12
<< pdcontact >>
rect 35 68 39 72
rect 3 49 7 53
rect 14 59 18 63
rect 24 59 28 63
rect 46 59 50 63
rect 56 61 60 65
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
<< psubstratepdiff >>
rect 0 2 64 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 64 2
rect 0 -3 64 -2
<< nsubstratendiff >>
rect 0 82 64 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 64 82
rect 0 77 64 78
<< labels >>
rlabel polycontact 12 36 12 36 6 zn
rlabel metal1 4 40 4 40 6 z
rlabel metal1 12 20 12 20 6 z
rlabel metal1 16 40 16 40 6 zn
rlabel metal1 32 6 32 6 6 vss
rlabel metal1 36 28 36 28 6 a
rlabel metal1 28 36 28 36 6 a
rlabel metal1 28 44 28 44 6 b
rlabel metal1 36 52 36 52 6 b
rlabel metal1 32 74 32 74 6 vdd
rlabel polycontact 44 44 44 44 6 c
rlabel metal1 44 36 44 36 6 d
rlabel metal1 44 52 44 52 6 b
rlabel metal1 37 61 37 61 6 zn
rlabel metal1 36 19 36 19 6 zn
rlabel metal1 60 24 60 24 6 d
rlabel metal1 52 36 52 36 6 d
rlabel metal1 52 44 52 44 6 c
rlabel metal1 60 52 60 52 6 c
<< end >>
