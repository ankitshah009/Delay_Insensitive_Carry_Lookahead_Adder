magic
tech scmos
timestamp 1179385450
<< checkpaint >>
rect -22 -25 54 105
<< ab >>
rect 0 0 32 80
<< pwell >>
rect -4 -7 36 36
<< nwell >>
rect -4 36 36 87
<< polysilicon >>
rect 9 57 11 62
rect 21 63 27 64
rect 21 59 22 63
rect 26 59 27 63
rect 21 58 27 59
rect 21 55 23 58
rect 9 39 11 45
rect 9 38 16 39
rect 9 34 11 38
rect 15 34 16 38
rect 9 33 16 34
rect 9 30 11 33
rect 21 30 23 45
rect 9 19 11 24
rect 21 18 23 23
<< ndiffusion >>
rect 2 29 9 30
rect 2 25 3 29
rect 7 25 9 29
rect 2 24 9 25
rect 11 28 21 30
rect 11 24 14 28
rect 18 24 21 28
rect 13 23 21 24
rect 23 29 30 30
rect 23 25 25 29
rect 29 25 30 29
rect 23 23 30 25
<< pdiffusion >>
rect 13 72 19 73
rect 13 68 14 72
rect 18 68 19 72
rect 13 57 19 68
rect 4 51 9 57
rect 2 50 9 51
rect 2 46 3 50
rect 7 46 9 50
rect 2 45 9 46
rect 11 55 19 57
rect 11 45 21 55
rect 23 51 28 55
rect 23 50 30 51
rect 23 46 25 50
rect 29 46 30 50
rect 23 45 30 46
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect -2 72 34 78
rect -2 68 14 72
rect 18 68 34 72
rect 18 59 22 63
rect 26 59 30 63
rect 18 57 30 59
rect 2 50 14 55
rect 2 46 3 50
rect 7 49 14 50
rect 18 49 22 57
rect 25 50 29 51
rect 2 45 7 46
rect 2 29 6 45
rect 25 38 29 46
rect 10 34 11 38
rect 15 34 30 38
rect 24 29 30 34
rect 2 25 3 29
rect 7 25 8 29
rect 14 28 18 29
rect 24 25 25 29
rect 29 25 30 29
rect 14 12 18 24
rect -2 2 34 12
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
<< ntransistor >>
rect 9 24 11 30
rect 21 23 23 30
<< ptransistor >>
rect 9 45 11 57
rect 21 45 23 55
<< polycontact >>
rect 22 59 26 63
rect 11 34 15 38
<< ndcontact >>
rect 3 25 7 29
rect 14 24 18 28
rect 25 25 29 29
<< pdcontact >>
rect 14 68 18 72
rect 3 46 7 50
rect 25 46 29 50
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
<< psubstratepdiff >>
rect 0 2 32 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 32 2
rect 0 -3 32 -2
<< nsubstratendiff >>
rect 0 82 32 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 32 82
rect 0 77 32 78
<< labels >>
rlabel polycontact 12 36 12 36 6 an
rlabel metal1 4 40 4 40 6 z
rlabel metal1 12 52 12 52 6 z
rlabel metal1 16 6 16 6 6 vss
rlabel metal1 20 56 20 56 6 a
rlabel metal1 16 74 16 74 6 vdd
rlabel metal1 20 36 20 36 6 an
rlabel metal1 27 38 27 38 6 an
rlabel metal1 28 60 28 60 6 a
<< end >>
