magic
tech scmos
timestamp 1179386702
<< checkpaint >>
rect -22 -25 126 105
<< ab >>
rect 0 0 104 80
<< pwell >>
rect -4 -7 108 36
<< nwell >>
rect -4 36 108 87
<< polysilicon >>
rect 9 70 11 74
rect 16 70 18 74
rect 26 70 28 74
rect 33 70 35 74
rect 43 70 45 74
rect 50 70 52 74
rect 60 70 62 74
rect 67 70 69 74
rect 78 61 80 66
rect 88 61 90 65
rect 9 33 11 42
rect 16 39 18 42
rect 26 39 28 42
rect 33 39 35 42
rect 43 39 45 42
rect 50 39 52 42
rect 60 39 62 42
rect 16 38 28 39
rect 16 37 23 38
rect 22 34 23 37
rect 27 34 28 38
rect 22 33 28 34
rect 32 38 46 39
rect 32 34 41 38
rect 45 34 46 38
rect 32 33 46 34
rect 9 32 15 33
rect 9 28 10 32
rect 14 28 15 32
rect 22 30 24 33
rect 32 30 34 33
rect 9 27 15 28
rect 44 22 46 33
rect 50 37 62 39
rect 67 39 69 42
rect 78 39 80 42
rect 88 39 90 42
rect 67 38 73 39
rect 50 30 56 37
rect 67 34 68 38
rect 72 34 73 38
rect 67 33 73 34
rect 78 38 90 39
rect 78 34 84 38
rect 88 34 90 38
rect 78 33 90 34
rect 78 30 80 33
rect 50 26 51 30
rect 55 26 56 30
rect 50 25 56 26
rect 54 22 56 25
rect 22 6 24 11
rect 32 6 34 11
rect 44 6 46 11
rect 54 6 56 11
rect 78 6 80 11
<< ndiffusion >>
rect 17 24 22 30
rect 13 15 22 24
rect 13 11 15 15
rect 19 11 22 15
rect 24 22 32 30
rect 24 18 26 22
rect 30 18 32 22
rect 24 11 32 18
rect 34 22 42 30
rect 71 29 78 30
rect 71 25 72 29
rect 76 25 78 29
rect 71 22 78 25
rect 34 15 44 22
rect 34 11 37 15
rect 41 11 44 15
rect 46 21 54 22
rect 46 17 48 21
rect 52 17 54 21
rect 46 11 54 17
rect 56 16 66 22
rect 71 18 72 22
rect 76 18 78 22
rect 71 17 78 18
rect 56 12 60 16
rect 64 12 66 16
rect 56 11 66 12
rect 73 11 78 17
rect 80 24 87 30
rect 80 20 82 24
rect 86 20 87 24
rect 80 16 87 20
rect 80 12 82 16
rect 86 12 87 16
rect 80 11 87 12
rect 13 9 20 11
rect 36 9 42 11
<< pdiffusion >>
rect 2 69 9 70
rect 2 65 3 69
rect 7 65 9 69
rect 2 62 9 65
rect 2 58 3 62
rect 7 58 9 62
rect 2 42 9 58
rect 11 42 16 70
rect 18 62 26 70
rect 18 58 20 62
rect 24 58 26 62
rect 18 54 26 58
rect 18 50 20 54
rect 24 50 26 54
rect 18 42 26 50
rect 28 42 33 70
rect 35 69 43 70
rect 35 65 37 69
rect 41 65 43 69
rect 35 62 43 65
rect 35 58 37 62
rect 41 58 43 62
rect 35 42 43 58
rect 45 42 50 70
rect 52 54 60 70
rect 52 50 54 54
rect 58 50 60 54
rect 52 47 60 50
rect 52 43 54 47
rect 58 43 60 47
rect 52 42 60 43
rect 62 42 67 70
rect 69 69 76 70
rect 69 65 71 69
rect 75 65 76 69
rect 69 62 76 65
rect 69 58 71 62
rect 75 61 76 62
rect 75 58 78 61
rect 69 55 78 58
rect 69 51 71 55
rect 75 51 78 55
rect 69 42 78 51
rect 80 54 88 61
rect 80 50 82 54
rect 86 50 88 54
rect 80 47 88 50
rect 80 43 82 47
rect 86 43 88 47
rect 80 42 88 43
rect 90 60 97 61
rect 90 56 92 60
rect 96 56 97 60
rect 90 42 97 56
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect -2 69 106 78
rect -2 68 3 69
rect 2 65 3 68
rect 7 68 37 69
rect 7 65 8 68
rect 2 62 8 65
rect 36 65 37 68
rect 41 68 71 69
rect 41 65 42 68
rect 2 58 3 62
rect 7 58 8 62
rect 18 62 24 63
rect 18 58 20 62
rect 36 62 42 65
rect 36 58 37 62
rect 41 58 42 62
rect 75 68 106 69
rect 71 62 75 65
rect 18 54 24 58
rect 71 55 75 58
rect 92 60 96 68
rect 92 55 96 56
rect 2 50 20 54
rect 24 50 54 54
rect 58 50 63 54
rect 71 50 75 51
rect 82 54 86 55
rect 2 22 6 50
rect 54 47 58 50
rect 14 42 40 46
rect 82 47 86 50
rect 54 42 58 43
rect 72 43 82 46
rect 72 42 86 43
rect 14 33 18 42
rect 36 38 40 42
rect 22 34 23 38
rect 27 34 31 38
rect 36 34 41 38
rect 45 34 68 38
rect 10 32 18 33
rect 14 28 18 32
rect 10 27 18 28
rect 25 30 31 34
rect 25 26 51 30
rect 55 26 63 30
rect 72 29 76 42
rect 90 38 94 47
rect 81 34 84 38
rect 88 34 94 38
rect 90 25 94 34
rect 72 22 76 25
rect 2 18 26 22
rect 30 21 55 22
rect 30 18 48 21
rect 47 17 48 18
rect 52 18 55 21
rect 52 17 53 18
rect 72 17 76 18
rect 82 24 86 25
rect 60 16 64 17
rect 14 12 15 15
rect -2 11 15 12
rect 19 12 20 15
rect 36 12 37 15
rect 19 11 37 12
rect 41 12 42 15
rect 82 16 86 20
rect 41 11 106 12
rect -2 2 106 11
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
<< ntransistor >>
rect 22 11 24 30
rect 32 11 34 30
rect 44 11 46 22
rect 54 11 56 22
rect 78 11 80 30
<< ptransistor >>
rect 9 42 11 70
rect 16 42 18 70
rect 26 42 28 70
rect 33 42 35 70
rect 43 42 45 70
rect 50 42 52 70
rect 60 42 62 70
rect 67 42 69 70
rect 78 42 80 61
rect 88 42 90 61
<< polycontact >>
rect 23 34 27 38
rect 41 34 45 38
rect 10 28 14 32
rect 68 34 72 38
rect 84 34 88 38
rect 51 26 55 30
<< ndcontact >>
rect 15 11 19 15
rect 26 18 30 22
rect 72 25 76 29
rect 37 11 41 15
rect 48 17 52 21
rect 72 18 76 22
rect 60 12 64 16
rect 82 20 86 24
rect 82 12 86 16
<< pdcontact >>
rect 3 65 7 69
rect 3 58 7 62
rect 20 58 24 62
rect 20 50 24 54
rect 37 65 41 69
rect 37 58 41 62
rect 54 50 58 54
rect 54 43 58 47
rect 71 65 75 69
rect 71 58 75 62
rect 71 51 75 55
rect 82 50 86 54
rect 82 43 86 47
rect 92 56 96 60
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
rect 90 -2 94 2
rect 98 -2 102 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
rect 90 78 94 82
rect 98 78 102 82
<< psubstratepdiff >>
rect 0 2 104 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 104 2
rect 0 -3 104 -2
<< nsubstratendiff >>
rect 0 82 104 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 104 82
rect 0 77 104 78
<< labels >>
rlabel polycontact 12 30 12 30 6 an
rlabel polysilicon 39 36 39 36 6 an
rlabel polycontact 70 36 70 36 6 an
rlabel metal1 12 20 12 20 6 z
rlabel metal1 14 30 14 30 6 an
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 52 12 52 6 z
rlabel metal1 20 20 20 20 6 z
rlabel ndcontact 28 20 28 20 6 z
rlabel metal1 36 20 36 20 6 z
rlabel metal1 36 28 36 28 6 b
rlabel metal1 28 32 28 32 6 b
rlabel metal1 28 52 28 52 6 z
rlabel metal1 36 52 36 52 6 z
rlabel metal1 20 56 20 56 6 z
rlabel metal1 52 6 52 6 6 vss
rlabel metal1 44 20 44 20 6 z
rlabel metal1 44 28 44 28 6 b
rlabel metal1 52 20 52 20 6 z
rlabel polycontact 52 28 52 28 6 b
rlabel metal1 60 28 60 28 6 b
rlabel metal1 52 52 52 52 6 z
rlabel metal1 60 52 60 52 6 z
rlabel metal1 44 52 44 52 6 z
rlabel metal1 52 74 52 74 6 vdd
rlabel metal1 74 31 74 31 6 an
rlabel metal1 56 36 56 36 6 an
rlabel metal1 84 36 84 36 6 a
rlabel metal1 92 36 92 36 6 a
rlabel metal1 84 48 84 48 6 an
<< end >>
