magic
tech scmos
timestamp 1185039112
<< checkpaint >>
rect -22 -24 122 124
<< ab >>
rect 0 0 100 100
<< pwell >>
rect -2 -4 102 49
<< nwell >>
rect -2 49 102 104
<< polysilicon >>
rect 73 95 75 98
rect 85 95 87 98
rect 11 85 13 88
rect 23 85 25 88
rect 35 85 37 88
rect 47 85 49 88
rect 11 43 13 65
rect 23 43 25 65
rect 7 42 13 43
rect 7 38 8 42
rect 12 38 13 42
rect 7 37 13 38
rect 17 42 25 43
rect 17 38 18 42
rect 22 38 25 42
rect 17 37 25 38
rect 11 25 13 37
rect 23 25 25 37
rect 35 43 37 65
rect 47 43 49 65
rect 73 43 75 55
rect 35 42 43 43
rect 35 38 38 42
rect 42 38 43 42
rect 35 37 43 38
rect 47 42 53 43
rect 47 38 48 42
rect 52 38 53 42
rect 47 37 53 38
rect 67 42 75 43
rect 67 38 68 42
rect 72 41 75 42
rect 85 41 87 55
rect 72 39 87 41
rect 72 38 75 39
rect 67 37 75 38
rect 35 25 37 37
rect 47 25 49 37
rect 73 25 75 37
rect 85 25 87 39
rect 11 12 13 15
rect 23 12 25 15
rect 35 12 37 15
rect 47 12 49 15
rect 73 2 75 5
rect 85 2 87 5
<< ndiffusion >>
rect 3 15 11 25
rect 13 15 23 25
rect 25 22 35 25
rect 25 18 28 22
rect 32 18 35 22
rect 25 15 35 18
rect 37 15 47 25
rect 49 15 57 25
rect 3 12 9 15
rect 51 12 57 15
rect 3 8 4 12
rect 8 8 9 12
rect 3 7 9 8
rect 51 8 52 12
rect 56 8 57 12
rect 51 7 57 8
rect 65 22 73 25
rect 65 18 66 22
rect 70 18 73 22
rect 65 12 73 18
rect 65 8 66 12
rect 70 8 73 12
rect 65 5 73 8
rect 75 22 85 25
rect 75 18 78 22
rect 82 18 85 22
rect 75 5 85 18
rect 87 22 95 25
rect 87 18 90 22
rect 94 18 95 22
rect 87 12 95 18
rect 87 8 90 12
rect 94 8 95 12
rect 87 5 95 8
<< pdiffusion >>
rect 39 92 45 93
rect 39 88 40 92
rect 44 88 45 92
rect 65 92 73 95
rect 65 88 66 92
rect 70 88 73 92
rect 39 85 45 88
rect 3 82 11 85
rect 3 78 4 82
rect 8 78 11 82
rect 3 65 11 78
rect 13 72 23 85
rect 13 68 16 72
rect 20 68 23 72
rect 13 65 23 68
rect 25 82 35 85
rect 25 78 28 82
rect 32 78 35 82
rect 25 65 35 78
rect 37 65 47 85
rect 49 82 57 85
rect 49 78 52 82
rect 56 78 57 82
rect 49 65 57 78
rect 65 82 73 88
rect 65 78 66 82
rect 70 78 73 82
rect 65 55 73 78
rect 75 82 85 95
rect 75 78 78 82
rect 82 78 85 82
rect 75 72 85 78
rect 75 68 78 72
rect 82 68 85 72
rect 75 62 85 68
rect 75 58 78 62
rect 82 58 85 62
rect 75 55 85 58
rect 87 92 95 95
rect 87 88 90 92
rect 94 88 95 92
rect 87 82 95 88
rect 87 78 90 82
rect 94 78 95 82
rect 87 72 95 78
rect 87 68 90 72
rect 94 68 95 72
rect 87 62 95 68
rect 87 58 90 62
rect 94 58 95 62
rect 87 55 95 58
<< metal1 >>
rect -2 96 102 101
rect -2 92 4 96
rect 8 92 16 96
rect 20 92 28 96
rect 32 92 102 96
rect -2 88 40 92
rect 44 88 66 92
rect 70 88 90 92
rect 94 88 102 92
rect -2 87 102 88
rect 3 82 9 83
rect 27 82 33 83
rect 51 82 57 83
rect 3 78 4 82
rect 8 78 28 82
rect 32 78 52 82
rect 56 78 57 82
rect 3 77 9 78
rect 27 77 33 78
rect 51 77 57 78
rect 65 82 71 87
rect 65 78 66 82
rect 70 78 71 82
rect 65 77 71 78
rect 77 82 83 83
rect 77 78 78 82
rect 82 78 83 82
rect 15 72 21 73
rect 77 72 83 78
rect 15 68 16 72
rect 20 68 72 72
rect 15 67 21 68
rect 7 42 13 62
rect 7 38 8 42
rect 12 38 13 42
rect 7 18 13 38
rect 17 42 23 62
rect 17 38 18 42
rect 22 38 23 42
rect 17 18 23 38
rect 28 23 32 68
rect 37 42 43 62
rect 37 38 38 42
rect 42 38 43 42
rect 27 22 33 23
rect 27 18 28 22
rect 32 18 33 22
rect 37 18 43 38
rect 47 42 53 62
rect 68 43 72 68
rect 77 68 78 72
rect 82 68 83 72
rect 77 62 83 68
rect 77 58 78 62
rect 82 58 83 62
rect 47 38 48 42
rect 52 38 53 42
rect 47 18 53 38
rect 67 42 73 43
rect 67 38 68 42
rect 72 38 73 42
rect 67 37 73 38
rect 65 22 71 23
rect 65 18 66 22
rect 70 18 71 22
rect 27 17 33 18
rect 65 13 71 18
rect 77 22 83 58
rect 89 82 95 87
rect 89 78 90 82
rect 94 78 95 82
rect 89 72 95 78
rect 89 68 90 72
rect 94 68 95 72
rect 89 62 95 68
rect 89 58 90 62
rect 94 58 95 62
rect 89 57 95 58
rect 77 18 78 22
rect 82 18 83 22
rect 77 17 83 18
rect 89 22 95 23
rect 89 18 90 22
rect 94 18 95 22
rect 89 13 95 18
rect -2 12 102 13
rect -2 8 4 12
rect 8 8 52 12
rect 56 8 66 12
rect 70 8 90 12
rect 94 8 102 12
rect -2 4 16 8
rect 20 4 28 8
rect 32 4 40 8
rect 44 4 102 8
rect -2 -1 102 4
<< ntransistor >>
rect 11 15 13 25
rect 23 15 25 25
rect 35 15 37 25
rect 47 15 49 25
rect 73 5 75 25
rect 85 5 87 25
<< ptransistor >>
rect 11 65 13 85
rect 23 65 25 85
rect 35 65 37 85
rect 47 65 49 85
rect 73 55 75 95
rect 85 55 87 95
<< polycontact >>
rect 8 38 12 42
rect 18 38 22 42
rect 38 38 42 42
rect 48 38 52 42
rect 68 38 72 42
<< ndcontact >>
rect 28 18 32 22
rect 4 8 8 12
rect 52 8 56 12
rect 66 18 70 22
rect 66 8 70 12
rect 78 18 82 22
rect 90 18 94 22
rect 90 8 94 12
<< pdcontact >>
rect 40 88 44 92
rect 66 88 70 92
rect 4 78 8 82
rect 16 68 20 72
rect 28 78 32 82
rect 52 78 56 82
rect 66 78 70 82
rect 78 78 82 82
rect 78 68 82 72
rect 78 58 82 62
rect 90 88 94 92
rect 90 78 94 82
rect 90 68 94 72
rect 90 58 94 62
<< psubstratepcontact >>
rect 16 4 20 8
rect 28 4 32 8
rect 40 4 44 8
<< nsubstratencontact >>
rect 4 92 8 96
rect 16 92 20 96
rect 28 92 32 96
<< psubstratepdiff >>
rect 15 8 45 9
rect 15 4 16 8
rect 20 4 28 8
rect 32 4 40 8
rect 44 4 45 8
rect 15 3 45 4
<< nsubstratendiff >>
rect 3 96 33 97
rect 3 92 4 96
rect 8 92 16 96
rect 20 92 28 96
rect 32 92 33 96
rect 3 91 33 92
<< labels >>
rlabel polycontact 10 40 10 40 6 i0
rlabel polycontact 20 40 20 40 6 i1
rlabel polycontact 20 40 20 40 6 i1
rlabel polycontact 10 40 10 40 6 i0
rlabel polycontact 40 40 40 40 6 i2
rlabel polycontact 40 40 40 40 6 i2
rlabel metal1 50 6 50 6 6 vss
rlabel metal1 50 6 50 6 6 vss
rlabel polycontact 50 40 50 40 6 i3
rlabel polycontact 50 40 50 40 6 i3
rlabel metal1 50 94 50 94 6 vdd
rlabel metal1 50 94 50 94 6 vdd
rlabel metal1 80 50 80 50 6 q
rlabel metal1 80 50 80 50 6 q
<< end >>
