.subckt nd2v6x4 a b vdd vss z
*   SPICE3 file   created from nd2v6x4.ext -      technology: scmos
m00 z      a      vdd    vdd p w=26u  l=2.3636u ad=130p     pd=36u      as=182p     ps=66u
m01 vdd    a      z      vdd p w=26u  l=2.3636u ad=182p     pd=66u      as=130p     ps=36u
m02 z      b      vdd    vdd p w=26u  l=2.3636u ad=130p     pd=36u      as=182p     ps=66u
m03 vdd    b      z      vdd p w=26u  l=2.3636u ad=182p     pd=66u      as=130p     ps=36u
m04 w1     a      vss    vss n w=18u  l=2.3636u ad=108p     pd=39u      as=126p     ps=50u
m05 vss    a      w1     vss n w=18u  l=2.3636u ad=126p     pd=50u      as=108p     ps=39u
m06 z      b      w1     vss n w=18u  l=2.3636u ad=90p      pd=28u      as=108p     ps=39u
m07 w1     b      z      vss n w=18u  l=2.3636u ad=108p     pd=39u      as=90p      ps=28u
C0  a      vdd    0.034f
C1  w1     z      0.169f
C2  vss    b      0.013f
C3  w1     a      0.023f
C4  z      a      0.279f
C5  vss    vdd    0.006f
C6  b      vdd    0.050f
C7  w1     vss    0.208f
C8  vss    z      0.041f
C9  w1     b      0.040f
C10 vss    a      0.098f
C11 z      b      0.299f
C12 z      vdd    0.186f
C13 b      a      0.211f
C14 w1     vss    0.002f
C16 z      vss    0.016f
C17 b      vss    0.126f
C18 a      vss    0.126f
.ends
