.subckt cgi2bv0x1 a b c vdd vss z
*   SPICE3 file   created from cgi2bv0x1.ext -      technology: scmos
m00 vdd    a      n1     vdd p w=27u  l=2.3636u ad=108p     pd=35u      as=125.667p ps=46u
m01 w1     a      vdd    vdd p w=27u  l=2.3636u ad=67.5p    pd=32u      as=108p     ps=35u
m02 z      bn     w1     vdd p w=27u  l=2.3636u ad=108p     pd=35u      as=67.5p    ps=32u
m03 n1     c      z      vdd p w=27u  l=2.3636u ad=125.667p pd=46u      as=108p     ps=35u
m04 vdd    bn     n1     vdd p w=27u  l=2.3636u ad=108p     pd=35u      as=125.667p ps=46u
m05 bn     b      vdd    vdd p w=27u  l=2.3636u ad=161p     pd=68u      as=108p     ps=35u
m06 vss    a      n3     vss n w=12u  l=2.3636u ad=73.5p    pd=27u      as=56p      ps=26u
m07 w2     a      vss    vss n w=12u  l=2.3636u ad=30p      pd=17u      as=73.5p    ps=27u
m08 z      bn     w2     vss n w=12u  l=2.3636u ad=48p      pd=20u      as=30p      ps=17u
m09 n3     c      z      vss n w=12u  l=2.3636u ad=56p      pd=26u      as=48p      ps=20u
m10 vss    bn     n3     vss n w=12u  l=2.3636u ad=73.5p    pd=27u      as=56p      ps=26u
m11 bn     b      vss    vss n w=12u  l=2.3636u ad=72p      pd=38u      as=73.5p    ps=27u
C0  z      a      0.098f
C1  vdd    c      0.018f
C2  n3     z      0.177f
C3  n1     bn     0.017f
C4  vdd    a      0.022f
C5  b      c      0.035f
C6  n3     vdd    0.005f
C7  b      a      0.015f
C8  c      bn     0.239f
C9  z      vdd    0.062f
C10 vss    n1     0.018f
C11 bn     a      0.119f
C12 n3     bn     0.005f
C13 vss    c      0.024f
C14 w1     n1     0.023f
C15 z      b      0.014f
C16 w2     n3     0.006f
C17 vdd    b      0.024f
C18 z      bn     0.065f
C19 vss    a      0.020f
C20 n3     vss    0.337f
C21 w2     z      0.008f
C22 vdd    bn     0.152f
C23 n1     c      0.025f
C24 vss    z      0.068f
C25 n1     a      0.042f
C26 b      bn     0.403f
C27 vss    vdd    0.004f
C28 n3     n1     0.038f
C29 z      w1     0.007f
C30 c      a      0.043f
C31 n3     c      0.097f
C32 w1     vdd    0.004f
C33 z      n1     0.191f
C34 vss    b      0.019f
C35 vdd    n1     0.403f
C36 z      c      0.116f
C37 vss    bn     0.125f
C38 n3     a      0.041f
C39 n3     vss    0.003f
C41 z      vss    0.003f
C43 b      vss    0.021f
C44 c      vss    0.021f
C45 bn     vss    0.041f
C46 a      vss    0.042f
.ends
