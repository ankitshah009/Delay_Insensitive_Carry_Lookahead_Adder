magic
tech scmos
timestamp 1185039105
<< checkpaint >>
rect -22 -24 82 124
<< ab >>
rect 0 0 60 100
<< pwell >>
rect -2 -4 62 49
<< nwell >>
rect -2 49 62 104
<< polysilicon >>
rect 47 95 49 98
rect 11 85 13 88
rect 23 85 25 88
rect 35 85 37 88
rect 11 43 13 65
rect 23 63 25 65
rect 17 62 25 63
rect 17 58 18 62
rect 22 58 25 62
rect 17 57 25 58
rect 35 53 37 65
rect 35 52 43 53
rect 35 48 38 52
rect 42 48 43 52
rect 35 47 43 48
rect 7 42 13 43
rect 7 38 8 42
rect 12 38 13 42
rect 7 37 13 38
rect 27 42 33 43
rect 27 38 28 42
rect 32 41 33 42
rect 47 41 49 55
rect 32 39 49 41
rect 32 38 33 39
rect 27 37 33 38
rect 11 25 13 37
rect 17 32 25 33
rect 17 28 18 32
rect 22 28 25 32
rect 17 27 25 28
rect 23 25 25 27
rect 35 32 43 33
rect 35 28 38 32
rect 42 28 43 32
rect 35 27 43 28
rect 35 25 37 27
rect 47 25 49 39
rect 11 12 13 15
rect 23 12 25 15
rect 35 12 37 15
rect 47 2 49 5
<< ndiffusion >>
rect 3 15 11 25
rect 13 15 23 25
rect 25 22 35 25
rect 25 18 28 22
rect 32 18 35 22
rect 25 15 35 18
rect 37 15 47 25
rect 3 12 9 15
rect 39 12 47 15
rect 3 8 4 12
rect 8 8 9 12
rect 3 7 9 8
rect 39 8 40 12
rect 44 8 47 12
rect 39 5 47 8
rect 49 22 57 25
rect 49 18 52 22
rect 56 18 57 22
rect 49 5 57 18
<< pdiffusion >>
rect 39 92 47 95
rect 39 88 40 92
rect 44 88 47 92
rect 39 85 47 88
rect 3 82 11 85
rect 3 78 4 82
rect 8 78 11 82
rect 3 72 11 78
rect 3 68 4 72
rect 8 68 11 72
rect 3 65 11 68
rect 13 72 23 85
rect 13 68 16 72
rect 20 68 23 72
rect 13 65 23 68
rect 25 82 35 85
rect 25 78 28 82
rect 32 78 35 82
rect 25 65 35 78
rect 37 65 47 85
rect 39 55 47 65
rect 49 82 57 95
rect 49 78 52 82
rect 56 78 57 82
rect 49 72 57 78
rect 49 68 52 72
rect 56 68 57 72
rect 49 62 57 68
rect 49 58 52 62
rect 56 58 57 62
rect 49 55 57 58
<< metal1 >>
rect -2 96 62 101
rect -2 92 4 96
rect 8 92 16 96
rect 20 92 28 96
rect 32 92 62 96
rect -2 88 40 92
rect 44 88 62 92
rect -2 87 62 88
rect 3 82 9 83
rect 27 82 33 83
rect 47 82 57 83
rect 3 78 4 82
rect 8 78 28 82
rect 32 78 33 82
rect 3 77 9 78
rect 27 77 33 78
rect 4 73 8 77
rect 3 72 9 73
rect 3 68 4 72
rect 8 68 9 72
rect 3 67 9 68
rect 15 72 21 73
rect 15 68 16 72
rect 20 68 32 72
rect 15 67 21 68
rect 17 62 23 63
rect 7 42 13 62
rect 7 38 8 42
rect 12 38 13 42
rect 7 18 13 38
rect 17 58 18 62
rect 22 58 23 62
rect 17 32 23 58
rect 28 43 32 68
rect 37 52 43 82
rect 37 48 38 52
rect 42 48 43 52
rect 27 42 33 43
rect 27 38 28 42
rect 32 38 33 42
rect 27 37 33 38
rect 17 28 18 32
rect 22 28 23 32
rect 17 18 23 28
rect 28 23 32 37
rect 37 32 43 48
rect 37 28 38 32
rect 42 28 43 32
rect 27 22 33 23
rect 27 18 28 22
rect 32 18 33 22
rect 37 18 43 28
rect 47 78 52 82
rect 56 78 57 82
rect 47 77 57 78
rect 47 73 53 77
rect 47 72 57 73
rect 47 68 52 72
rect 56 68 57 72
rect 47 67 57 68
rect 47 63 53 67
rect 47 62 57 63
rect 47 58 52 62
rect 56 58 57 62
rect 47 57 57 58
rect 47 23 53 57
rect 47 22 57 23
rect 47 18 52 22
rect 56 18 57 22
rect 27 17 33 18
rect 47 17 57 18
rect -2 12 62 13
rect -2 8 4 12
rect 8 8 40 12
rect 44 8 62 12
rect -2 4 16 8
rect 20 4 28 8
rect 32 4 62 8
rect -2 -1 62 4
<< ntransistor >>
rect 11 15 13 25
rect 23 15 25 25
rect 35 15 37 25
rect 47 5 49 25
<< ptransistor >>
rect 11 65 13 85
rect 23 65 25 85
rect 35 65 37 85
rect 47 55 49 95
<< polycontact >>
rect 18 58 22 62
rect 38 48 42 52
rect 8 38 12 42
rect 28 38 32 42
rect 18 28 22 32
rect 38 28 42 32
<< ndcontact >>
rect 28 18 32 22
rect 4 8 8 12
rect 40 8 44 12
rect 52 18 56 22
<< pdcontact >>
rect 40 88 44 92
rect 4 78 8 82
rect 4 68 8 72
rect 16 68 20 72
rect 28 78 32 82
rect 52 78 56 82
rect 52 68 56 72
rect 52 58 56 62
<< psubstratepcontact >>
rect 16 4 20 8
rect 28 4 32 8
<< nsubstratencontact >>
rect 4 92 8 96
rect 16 92 20 96
rect 28 92 32 96
<< psubstratepdiff >>
rect 15 8 33 9
rect 15 4 16 8
rect 20 4 28 8
rect 32 4 33 8
rect 15 3 33 4
<< nsubstratendiff >>
rect 3 96 33 97
rect 3 92 4 96
rect 8 92 16 96
rect 20 92 28 96
rect 32 92 33 96
rect 3 91 33 92
<< labels >>
rlabel polycontact 10 40 10 40 6 i0
rlabel polycontact 10 40 10 40 6 i0
rlabel metal1 20 40 20 40 6 i1
rlabel metal1 20 40 20 40 6 i1
rlabel psubstratepcontact 30 6 30 6 6 vss
rlabel psubstratepcontact 30 6 30 6 6 vss
rlabel polycontact 40 50 40 50 6 i2
rlabel polycontact 40 50 40 50 6 i2
rlabel nsubstratencontact 30 94 30 94 6 vdd
rlabel nsubstratencontact 30 94 30 94 6 vdd
rlabel metal1 50 50 50 50 6 q
rlabel metal1 50 50 50 50 6 q
<< end >>
