magic
tech scmos
timestamp 1179385959
<< checkpaint >>
rect -22 -22 62 94
<< ab >>
rect 0 0 40 72
<< pwell >>
rect -4 -4 44 32
<< nwell >>
rect -4 32 44 76
<< polysilicon >>
rect 19 64 21 69
rect 29 64 31 69
rect 9 54 11 59
rect 9 35 11 38
rect 19 35 21 38
rect 29 35 31 38
rect 9 34 31 35
rect 9 30 16 34
rect 20 33 31 34
rect 20 30 21 33
rect 9 29 21 30
rect 9 26 11 29
rect 9 4 11 9
<< ndiffusion >>
rect 2 25 9 26
rect 2 21 3 25
rect 7 21 9 25
rect 2 18 9 21
rect 2 14 3 18
rect 7 14 9 18
rect 2 13 9 14
rect 4 9 9 13
rect 11 22 19 26
rect 11 18 13 22
rect 17 18 19 22
rect 11 14 19 18
rect 11 10 13 14
rect 17 10 19 14
rect 11 9 19 10
<< pdiffusion >>
rect 13 54 19 64
rect 4 51 9 54
rect 2 50 9 51
rect 2 46 3 50
rect 7 46 9 50
rect 2 43 9 46
rect 2 39 3 43
rect 7 39 9 43
rect 2 38 9 39
rect 11 53 19 54
rect 11 49 13 53
rect 17 49 19 53
rect 11 38 19 49
rect 21 50 29 64
rect 21 46 23 50
rect 27 46 29 50
rect 21 43 29 46
rect 21 39 23 43
rect 27 39 29 43
rect 21 38 29 39
rect 31 63 38 64
rect 31 59 33 63
rect 37 59 38 63
rect 31 55 38 59
rect 31 51 33 55
rect 37 51 38 55
rect 31 38 38 51
<< metal1 >>
rect -2 68 42 72
rect -2 64 4 68
rect 8 64 42 68
rect 13 53 17 64
rect 2 50 7 51
rect 2 46 3 50
rect 33 63 37 64
rect 33 55 37 59
rect 13 48 17 49
rect 23 50 27 51
rect 33 50 37 51
rect 2 43 7 46
rect 2 39 3 43
rect 23 43 27 46
rect 7 39 23 42
rect 27 39 31 42
rect 2 38 31 39
rect 2 26 6 38
rect 15 30 16 34
rect 20 30 31 34
rect 2 25 7 26
rect 2 21 3 25
rect 2 18 7 21
rect 2 14 3 18
rect 2 13 7 14
rect 13 22 17 23
rect 25 22 31 30
rect 13 14 17 18
rect 13 8 17 10
rect -2 4 24 8
rect 28 4 32 8
rect 36 4 42 8
rect -2 0 42 4
<< ntransistor >>
rect 9 9 11 26
<< ptransistor >>
rect 9 38 11 54
rect 19 38 21 64
rect 29 38 31 64
<< polycontact >>
rect 16 30 20 34
<< ndcontact >>
rect 3 21 7 25
rect 3 14 7 18
rect 13 18 17 22
rect 13 10 17 14
<< pdcontact >>
rect 3 46 7 50
rect 3 39 7 43
rect 13 49 17 53
rect 23 46 27 50
rect 23 39 27 43
rect 33 59 37 63
rect 33 51 37 55
<< psubstratepcontact >>
rect 24 4 28 8
rect 32 4 36 8
<< nsubstratencontact >>
rect 4 64 8 68
<< psubstratepdiff >>
rect 23 8 37 24
rect 23 4 24 8
rect 28 4 32 8
rect 36 4 37 8
rect 23 3 37 4
<< nsubstratendiff >>
rect 3 68 9 69
rect 3 64 4 68
rect 8 64 9 68
rect 3 62 9 64
<< labels >>
rlabel metal1 4 32 4 32 6 z
rlabel metal1 12 40 12 40 6 z
rlabel metal1 20 4 20 4 6 vss
rlabel metal1 20 32 20 32 6 a
rlabel metal1 28 28 28 28 6 a
rlabel metal1 28 40 28 40 6 z
rlabel metal1 20 40 20 40 6 z
rlabel metal1 20 68 20 68 6 vdd
<< end >>
