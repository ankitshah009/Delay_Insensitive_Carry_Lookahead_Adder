magic
tech scmos
timestamp 1185094696
<< checkpaint >>
rect -22 -22 172 122
<< ab >>
rect 0 0 150 100
<< pwell >>
rect -4 -4 154 48
<< nwell >>
rect -4 48 154 104
<< polysilicon >>
rect 11 83 13 88
rect 23 83 25 88
rect 35 83 37 88
rect 47 83 49 88
rect 59 83 61 88
rect 67 83 69 88
rect 79 83 81 88
rect 87 83 89 88
rect 99 83 101 88
rect 111 83 113 88
rect 123 83 125 88
rect 135 83 137 88
rect 11 53 13 57
rect 7 52 13 53
rect 7 48 8 52
rect 12 48 13 52
rect 7 47 13 48
rect 11 39 13 47
rect 23 53 25 57
rect 35 53 37 57
rect 23 52 37 53
rect 47 54 49 57
rect 59 54 61 57
rect 47 52 63 54
rect 23 48 28 52
rect 32 48 37 52
rect 57 48 58 52
rect 62 48 63 52
rect 23 47 37 48
rect 23 30 25 47
rect 35 30 37 47
rect 47 47 53 48
rect 57 47 63 48
rect 47 43 48 47
rect 52 43 53 47
rect 47 42 53 43
rect 47 39 49 42
rect 59 30 61 47
rect 67 43 69 57
rect 79 43 81 57
rect 67 42 81 43
rect 67 38 72 42
rect 76 38 81 42
rect 67 37 81 38
rect 67 30 69 37
rect 79 30 81 37
rect 87 53 89 57
rect 99 53 101 57
rect 111 53 113 57
rect 87 52 93 53
rect 87 48 88 52
rect 92 48 93 52
rect 87 47 93 48
rect 97 52 113 53
rect 97 48 98 52
rect 102 51 113 52
rect 102 48 103 51
rect 97 47 103 48
rect 123 47 125 55
rect 135 47 137 55
rect 87 30 89 47
rect 118 46 137 47
rect 118 42 119 46
rect 123 45 137 46
rect 123 42 125 45
rect 118 41 125 42
rect 123 37 125 41
rect 135 37 137 45
rect 11 13 13 18
rect 23 13 25 18
rect 35 13 37 18
rect 47 13 49 18
rect 59 13 61 18
rect 67 13 69 18
rect 79 13 81 18
rect 87 13 89 18
rect 123 17 125 22
rect 135 17 137 22
<< ndiffusion >>
rect 3 32 11 39
rect 3 28 4 32
rect 8 28 11 32
rect 3 24 11 28
rect 3 20 4 24
rect 8 20 11 24
rect 3 18 11 20
rect 13 30 18 39
rect 42 30 47 39
rect 13 23 23 30
rect 13 19 16 23
rect 20 19 23 23
rect 13 18 23 19
rect 25 29 35 30
rect 25 25 28 29
rect 32 25 35 29
rect 25 18 35 25
rect 37 23 47 30
rect 37 19 40 23
rect 44 19 47 23
rect 37 18 47 19
rect 49 30 57 39
rect 114 36 123 37
rect 114 32 116 36
rect 120 32 123 36
rect 49 23 59 30
rect 49 19 52 23
rect 56 19 59 23
rect 49 18 59 19
rect 61 18 67 30
rect 69 28 79 30
rect 69 24 72 28
rect 76 24 79 28
rect 69 18 79 24
rect 81 18 87 30
rect 89 23 98 30
rect 89 19 92 23
rect 96 19 98 23
rect 114 28 123 32
rect 114 24 116 28
rect 120 24 123 28
rect 114 22 123 24
rect 125 36 135 37
rect 125 32 128 36
rect 132 32 135 36
rect 125 28 135 32
rect 125 24 128 28
rect 132 24 135 28
rect 125 22 135 24
rect 137 36 146 37
rect 137 32 140 36
rect 144 32 146 36
rect 137 28 146 32
rect 137 24 140 28
rect 144 24 146 28
rect 137 22 146 24
rect 89 18 98 19
<< pdiffusion >>
rect 51 92 57 93
rect 51 88 52 92
rect 56 88 57 92
rect 91 92 97 93
rect 91 88 92 92
rect 96 88 97 92
rect 51 83 57 88
rect 91 83 97 88
rect 3 82 11 83
rect 3 78 4 82
rect 8 78 11 82
rect 3 57 11 78
rect 13 82 23 83
rect 13 78 16 82
rect 20 78 23 82
rect 13 57 23 78
rect 25 62 35 83
rect 25 58 28 62
rect 32 58 35 62
rect 25 57 35 58
rect 37 82 47 83
rect 37 78 40 82
rect 44 78 47 82
rect 37 57 47 78
rect 49 57 59 83
rect 61 57 67 83
rect 69 62 79 83
rect 69 58 72 62
rect 76 58 79 62
rect 69 57 79 58
rect 81 57 87 83
rect 89 57 99 83
rect 101 80 111 83
rect 101 76 104 80
rect 108 76 111 80
rect 101 72 111 76
rect 101 68 104 72
rect 108 68 111 72
rect 101 57 111 68
rect 113 82 123 83
rect 113 78 116 82
rect 120 78 123 82
rect 113 72 123 78
rect 113 68 116 72
rect 120 68 123 72
rect 113 57 123 68
rect 115 55 123 57
rect 125 72 135 83
rect 125 68 128 72
rect 132 68 135 72
rect 125 62 135 68
rect 125 58 128 62
rect 132 58 135 62
rect 125 55 135 58
rect 137 82 146 83
rect 137 78 140 82
rect 144 78 146 82
rect 137 72 146 78
rect 137 68 140 72
rect 144 68 146 72
rect 137 55 146 68
<< metal1 >>
rect -2 96 152 100
rect -2 92 8 96
rect 12 92 18 96
rect 22 92 152 96
rect -2 88 52 92
rect 56 88 92 92
rect 96 88 152 92
rect 4 82 8 88
rect 116 82 120 88
rect 15 78 16 82
rect 20 78 40 82
rect 44 80 108 82
rect 44 78 104 80
rect 4 77 8 78
rect 104 72 108 76
rect 8 68 93 72
rect 8 52 12 68
rect 8 47 12 48
rect 18 52 22 63
rect 27 58 28 62
rect 32 58 72 62
rect 76 58 77 62
rect 18 48 28 52
rect 32 48 33 52
rect 18 37 22 48
rect 4 32 8 33
rect 38 32 42 58
rect 87 52 93 68
rect 104 67 108 68
rect 116 72 120 78
rect 140 82 144 88
rect 116 67 120 68
rect 128 72 132 73
rect 128 62 132 68
rect 140 72 144 78
rect 140 67 144 68
rect 57 48 58 52
rect 62 48 88 52
rect 92 48 93 52
rect 97 52 103 62
rect 97 48 98 52
rect 102 48 103 52
rect 47 47 53 48
rect 47 43 48 47
rect 52 43 53 47
rect 47 42 53 43
rect 97 42 103 48
rect 128 52 132 58
rect 128 48 143 52
rect 47 38 72 42
rect 76 38 103 42
rect 108 42 119 46
rect 123 42 124 46
rect 108 32 112 42
rect 4 24 8 28
rect 27 29 112 32
rect 27 25 28 29
rect 32 28 112 29
rect 116 36 120 37
rect 116 28 120 32
rect 32 25 33 28
rect 52 23 56 24
rect 72 23 76 24
rect 92 23 96 24
rect 4 12 8 20
rect 15 19 16 23
rect 20 21 21 23
rect 39 21 40 23
rect 20 19 40 21
rect 44 19 45 23
rect 15 17 45 19
rect 52 12 56 19
rect 92 12 96 19
rect 116 12 120 24
rect 128 36 132 48
rect 128 28 132 32
rect 128 23 132 24
rect 140 36 144 37
rect 140 28 144 32
rect 140 12 144 24
rect -2 8 152 12
rect -2 4 8 8
rect 12 4 18 8
rect 22 4 152 8
rect -2 0 152 4
<< ntransistor >>
rect 11 18 13 39
rect 23 18 25 30
rect 35 18 37 30
rect 47 18 49 39
rect 59 18 61 30
rect 67 18 69 30
rect 79 18 81 30
rect 87 18 89 30
rect 123 22 125 37
rect 135 22 137 37
<< ptransistor >>
rect 11 57 13 83
rect 23 57 25 83
rect 35 57 37 83
rect 47 57 49 83
rect 59 57 61 83
rect 67 57 69 83
rect 79 57 81 83
rect 87 57 89 83
rect 99 57 101 83
rect 111 57 113 83
rect 123 55 125 83
rect 135 55 137 83
<< polycontact >>
rect 8 48 12 52
rect 28 48 32 52
rect 58 48 62 52
rect 48 43 52 47
rect 72 38 76 42
rect 88 48 92 52
rect 98 48 102 52
rect 119 42 123 46
<< ndcontact >>
rect 4 28 8 32
rect 4 20 8 24
rect 16 19 20 23
rect 28 25 32 29
rect 40 19 44 23
rect 116 32 120 36
rect 52 19 56 23
rect 72 24 76 28
rect 92 19 96 23
rect 116 24 120 28
rect 128 32 132 36
rect 128 24 132 28
rect 140 32 144 36
rect 140 24 144 28
<< pdcontact >>
rect 52 88 56 92
rect 92 88 96 92
rect 4 78 8 82
rect 16 78 20 82
rect 28 58 32 62
rect 40 78 44 82
rect 72 58 76 62
rect 104 76 108 80
rect 104 68 108 72
rect 116 78 120 82
rect 116 68 120 72
rect 128 68 132 72
rect 128 58 132 62
rect 140 78 144 82
rect 140 68 144 72
<< psubstratepcontact >>
rect 8 4 12 8
rect 18 4 22 8
<< nsubstratencontact >>
rect 8 92 12 96
rect 18 92 22 96
<< psubstratepdiff >>
rect 7 8 23 9
rect 7 4 8 8
rect 12 4 18 8
rect 22 4 23 8
rect 7 3 23 4
<< nsubstratendiff >>
rect 7 96 23 97
rect 7 92 8 96
rect 12 92 18 96
rect 22 92 23 96
rect 7 91 23 92
<< labels >>
rlabel polycontact 121 44 121 44 6 zn
rlabel ndcontact 18 20 18 20 6 n4
rlabel metal1 20 50 20 50 6 c
rlabel metal1 10 60 10 60 6 a
rlabel metal1 20 70 20 70 6 a
rlabel ndcontact 42 20 42 20 6 n4
rlabel ndcontact 30 28 30 28 6 zn
rlabel metal1 50 40 50 40 6 b
rlabel polycontact 30 50 30 50 6 c
rlabel metal1 30 70 30 70 6 a
rlabel metal1 50 70 50 70 6 a
rlabel metal1 40 70 40 70 6 a
rlabel metal1 75 6 75 6 6 vss
rlabel ndcontact 74 27 74 27 6 zn
rlabel metal1 80 40 80 40 6 b
rlabel metal1 70 40 70 40 6 b
rlabel metal1 60 40 60 40 6 b
rlabel polycontact 60 50 60 50 6 a
rlabel metal1 80 50 80 50 6 a
rlabel metal1 70 50 70 50 6 a
rlabel metal1 52 60 52 60 6 zn
rlabel metal1 60 70 60 70 6 a
rlabel metal1 80 70 80 70 6 a
rlabel metal1 70 70 70 70 6 a
rlabel metal1 75 94 75 94 6 vdd
rlabel metal1 90 40 90 40 6 b
rlabel polycontact 100 50 100 50 6 b
rlabel metal1 90 60 90 60 6 a
rlabel metal1 106 74 106 74 6 n2
rlabel metal1 61 80 61 80 6 n2
rlabel metal1 116 44 116 44 6 zn
rlabel metal1 130 50 130 50 6 z
rlabel metal1 140 50 140 50 6 z
<< end >>
