.subckt o3_x2 i0 i1 i2 q vdd vss
*   SPICE3 file   created from o3_x2.ext -      technology: scmos
m00 w1     i2     w2     vdd p w=30u  l=2.3636u ad=90p      pd=36u      as=240p     ps=76u
m01 w3     i1     w1     vdd p w=30u  l=2.3636u ad=90p      pd=36u      as=90p      ps=36u
m02 vdd    i0     w3     vdd p w=30u  l=2.3636u ad=300p     pd=49.7143u as=90p      ps=36u
m03 q      w2     vdd    vdd p w=40u  l=2.3636u ad=320p     pd=96u      as=400p     ps=66.2857u
m04 vss    i2     w2     vss n w=10u  l=2.3636u ad=65.6p    pd=23.2u    as=60p      ps=25.3333u
m05 w2     i1     vss    vss n w=10u  l=2.3636u ad=60p      pd=25.3333u as=65.6p    ps=23.2u
m06 vss    i0     w2     vss n w=10u  l=2.3636u ad=65.6p    pd=23.2u    as=60p      ps=25.3333u
m07 q      w2     vss    vss n w=20u  l=2.3636u ad=160p     pd=56u      as=131.2p   ps=46.4u
C0  i0     i2     0.131f
C1  w1     w2     0.012f
C2  vss    q      0.099f
C3  i1     w2     0.187f
C4  i0     vdd    0.041f
C5  i2     vdd    0.015f
C6  vss    i1     0.015f
C7  q      i0     0.095f
C8  vss    w2     0.297f
C9  q      i2     0.040f
C10 w3     i1     0.018f
C11 q      vdd    0.123f
C12 i0     i1     0.410f
C13 w1     i2     0.009f
C14 w3     w2     0.012f
C15 i0     w2     0.413f
C16 i1     i2     0.436f
C17 i1     vdd    0.017f
C18 i2     w2     0.181f
C19 vss    i0     0.015f
C20 w2     vdd    0.330f
C21 q      i1     0.056f
C22 vss    i2     0.015f
C23 w3     i0     0.009f
C24 w1     i1     0.018f
C25 q      w2     0.429f
C27 q      vss    0.015f
C28 i0     vss    0.032f
C29 i1     vss    0.032f
C30 i2     vss    0.031f
C31 w2     vss    0.036f
.ends
