.subckt xaon21_x05 a1 a2 b vdd vss z
*   SPICE3 file   created from xaon21_x05.ext -      technology: scmos
m00 vdd    a1     an     vdd p w=20u  l=2.3636u ad=140p     pd=40.6667u as=106p     ps=38.6667u
m01 an     a2     vdd    vdd p w=20u  l=2.3636u ad=106p     pd=38.6667u as=140p     ps=40.6667u
m02 z      bn     an     vdd p w=20u  l=2.3636u ad=100p     pd=30u      as=106p     ps=38.6667u
m03 bn     an     z      vdd p w=20u  l=2.3636u ad=103p     pd=32u      as=100p     ps=30u
m04 vdd    b      bn     vdd p w=20u  l=2.3636u ad=140p     pd=40.6667u as=103p     ps=32u
m05 w1     a1     vss    vss n w=12u  l=2.3636u ad=36p      pd=18u      as=176.8p   ps=58.4u
m06 an     a2     w1     vss n w=12u  l=2.3636u ad=64.5p    pd=25u      as=36p      ps=18u
m07 z      b      an     vss n w=12u  l=2.3636u ad=60p      pd=25.1429u as=64.5p    ps=25u
m08 w2     bn     z      vss n w=9u   l=2.3636u ad=27p      pd=15u      as=45p      ps=18.8571u
m09 vss    an     w2     vss n w=9u   l=2.3636u ad=132.6p   pd=43.8u    as=27p      ps=15u
m10 bn     b      vss    vss n w=9u   l=2.3636u ad=63p      pd=34u      as=132.6p   ps=43.8u
C0  z      bn     0.070f
C1  vss    a2     0.007f
C2  b      an     0.243f
C3  w1     a1     0.006f
C4  an     bn     0.386f
C5  b      a2     0.037f
C6  z      a1     0.042f
C7  an     a1     0.062f
C8  bn     a2     0.070f
C9  a2     a1     0.113f
C10 bn     vdd    0.192f
C11 vss    b      0.147f
C12 a1     vdd    0.001f
C13 vss    bn     0.014f
C14 z      an     0.411f
C15 b      bn     0.175f
C16 z      a2     0.162f
C17 vss    a1     0.064f
C18 z      vdd    0.018f
C19 an     a2     0.184f
C20 b      a1     0.014f
C21 bn     a1     0.020f
C22 an     vdd    0.192f
C23 vss    z      0.028f
C24 w2     an     0.007f
C25 a2     vdd    0.041f
C26 z      b      0.036f
C27 vss    an     0.168f
C29 z      vss    0.015f
C30 b      vss    0.063f
C31 an     vss    0.038f
C32 bn     vss    0.042f
C33 a2     vss    0.035f
C34 a1     vss    0.031f
.ends
