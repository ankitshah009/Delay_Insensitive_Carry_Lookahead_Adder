.subckt oan21v0x05 a1 a2 b vdd vss z
*   SPICE3 file   created from oan21v0x05.ext -      technology: scmos
m00 vdd    zn     z      vdd p w=12u  l=2.3636u ad=160.457p pd=43.2u    as=72p      ps=38u
m01 zn     b      vdd    vdd p w=8u   l=2.3636u ad=34.4348p pd=16u      as=106.971p ps=28.8u
m02 w1     a2     zn     vdd p w=15u  l=2.3636u ad=37.5p    pd=20u      as=64.5652p ps=30u
m03 vdd    a1     w1     vdd p w=15u  l=2.3636u ad=200.571p pd=54u      as=37.5p    ps=20u
m04 vss    zn     z      vss n w=6u   l=2.3636u ad=62.4p    pd=27.6u    as=42p      ps=26u
m05 n1     b      zn     vss n w=7u   l=2.3636u ad=35p      pd=19.3333u as=49p      ps=28u
m06 vss    a2     n1     vss n w=7u   l=2.3636u ad=72.8p    pd=32.2u    as=35p      ps=19.3333u
m07 n1     a1     vss    vss n w=7u   l=2.3636u ad=35p      pd=19.3333u as=72.8p    ps=32.2u
C0  w1     vdd    0.004f
C1  z      a2     0.012f
C2  zn     a1     0.022f
C3  n1     vss    0.202f
C4  zn     vdd    0.210f
C5  b      a2     0.095f
C6  n1     z      0.014f
C7  a1     vdd    0.029f
C8  vss    zn     0.082f
C9  n1     b      0.021f
C10 w1     b      0.003f
C11 z      zn     0.093f
C12 vss    a1     0.017f
C13 n1     a2     0.118f
C14 zn     b      0.137f
C15 vss    vdd    0.008f
C16 z      a1     0.004f
C17 zn     a2     0.039f
C18 z      vdd    0.041f
C19 b      a1     0.054f
C20 b      vdd    0.034f
C21 a1     a2     0.123f
C22 vss    z      0.097f
C23 n1     zn     0.030f
C24 a2     vdd    0.016f
C25 n1     a1     0.022f
C26 vss    b      0.016f
C27 z      b      0.011f
C28 vss    a2     0.048f
C29 n1     vdd    0.007f
C30 n1     vss    0.005f
C32 z      vss    0.009f
C33 zn     vss    0.026f
C34 b      vss    0.028f
C35 a1     vss    0.032f
C36 a2     vss    0.026f
.ends
