magic
tech scmos
timestamp 1179386983
<< checkpaint >>
rect -22 -22 86 94
<< ab >>
rect 0 0 64 72
<< pwell >>
rect -4 -4 68 32
<< nwell >>
rect -4 32 68 76
<< polysilicon >>
rect 19 62 21 67
rect 26 62 28 67
rect 9 54 11 59
rect 40 58 42 63
rect 9 34 11 46
rect 9 33 15 34
rect 9 29 10 33
rect 14 29 15 33
rect 9 28 15 29
rect 19 28 21 46
rect 26 43 28 46
rect 40 43 42 46
rect 26 42 33 43
rect 26 38 27 42
rect 31 38 33 42
rect 40 42 55 43
rect 40 41 50 42
rect 26 37 33 38
rect 49 38 50 41
rect 54 38 55 42
rect 49 37 55 38
rect 9 19 11 28
rect 19 27 25 28
rect 19 23 20 27
rect 24 23 25 27
rect 19 22 25 23
rect 19 19 21 22
rect 31 19 33 37
rect 51 26 53 37
rect 51 15 53 20
rect 9 7 11 12
rect 19 7 21 12
rect 31 7 33 12
<< ndiffusion >>
rect 44 25 51 26
rect 44 21 45 25
rect 49 21 51 25
rect 44 20 51 21
rect 53 25 60 26
rect 53 21 55 25
rect 59 21 60 25
rect 53 20 60 21
rect 2 18 9 19
rect 2 14 3 18
rect 7 14 9 18
rect 2 12 9 14
rect 11 17 19 19
rect 11 13 13 17
rect 17 13 19 17
rect 11 12 19 13
rect 21 12 31 19
rect 33 17 40 19
rect 33 13 35 17
rect 39 13 40 17
rect 33 12 40 13
rect 23 8 29 12
rect 23 4 24 8
rect 28 4 29 8
rect 23 3 29 4
<< pdiffusion >>
rect 14 54 19 62
rect 2 53 9 54
rect 2 49 3 53
rect 7 49 9 53
rect 2 46 9 49
rect 11 51 19 54
rect 11 47 13 51
rect 17 47 19 51
rect 11 46 19 47
rect 21 46 26 62
rect 28 58 37 62
rect 28 57 40 58
rect 28 53 34 57
rect 38 53 40 57
rect 28 46 40 53
rect 42 52 47 58
rect 42 51 49 52
rect 42 47 44 51
rect 48 47 49 51
rect 42 46 49 47
<< metal1 >>
rect -2 68 66 72
rect -2 64 4 68
rect 8 64 56 68
rect 60 64 66 68
rect 3 53 7 64
rect 34 57 38 64
rect 34 52 38 53
rect 3 48 7 49
rect 10 47 13 51
rect 17 47 22 51
rect 10 45 22 47
rect 10 43 14 45
rect 2 39 14 43
rect 26 42 30 51
rect 42 47 44 51
rect 48 47 49 51
rect 2 19 6 39
rect 26 38 27 42
rect 31 38 39 42
rect 10 33 23 34
rect 14 30 23 33
rect 10 21 14 29
rect 42 27 46 47
rect 50 42 62 43
rect 54 38 62 42
rect 50 37 62 38
rect 58 29 62 37
rect 19 23 20 27
rect 24 25 46 27
rect 24 23 45 25
rect 42 21 45 23
rect 49 21 50 25
rect 54 21 55 25
rect 59 21 60 25
rect 2 18 7 19
rect 2 14 3 18
rect 2 13 7 14
rect 12 13 13 17
rect 17 13 35 17
rect 39 13 40 17
rect 54 8 60 21
rect -2 4 24 8
rect 28 4 48 8
rect 52 4 56 8
rect 60 4 66 8
rect -2 0 66 4
<< ntransistor >>
rect 51 20 53 26
rect 9 12 11 19
rect 19 12 21 19
rect 31 12 33 19
<< ptransistor >>
rect 9 46 11 54
rect 19 46 21 62
rect 26 46 28 62
rect 40 46 42 58
<< polycontact >>
rect 10 29 14 33
rect 27 38 31 42
rect 50 38 54 42
rect 20 23 24 27
<< ndcontact >>
rect 45 21 49 25
rect 55 21 59 25
rect 3 14 7 18
rect 13 13 17 17
rect 35 13 39 17
rect 24 4 28 8
<< pdcontact >>
rect 3 49 7 53
rect 13 47 17 51
rect 34 53 38 57
rect 44 47 48 51
<< psubstratepcontact >>
rect 48 4 52 8
rect 56 4 60 8
<< nsubstratencontact >>
rect 4 64 8 68
rect 56 64 60 68
<< psubstratepdiff >>
rect 47 8 61 9
rect 47 4 48 8
rect 52 4 56 8
rect 60 4 61 8
rect 47 3 61 4
<< nsubstratendiff >>
rect 3 68 9 69
rect 3 64 4 68
rect 8 64 9 68
rect 55 68 61 69
rect 3 63 9 64
rect 55 64 56 68
rect 60 64 61 68
rect 55 46 61 64
<< labels >>
rlabel polycontact 22 25 22 25 6 a2n
rlabel metal1 4 28 4 28 6 z
rlabel metal1 12 24 12 24 6 b
rlabel metal1 12 48 12 48 6 z
rlabel metal1 20 32 20 32 6 b
rlabel metal1 28 48 28 48 6 a1
rlabel metal1 20 48 20 48 6 z
rlabel metal1 32 4 32 4 6 vss
rlabel metal1 26 15 26 15 6 n1
rlabel metal1 32 25 32 25 6 a2n
rlabel metal1 44 36 44 36 6 a2n
rlabel metal1 36 40 36 40 6 a1
rlabel pdcontact 45 49 45 49 6 a2n
rlabel metal1 32 68 32 68 6 vdd
rlabel metal1 60 36 60 36 6 a2
rlabel polycontact 52 40 52 40 6 a2
<< end >>
