magic
tech scmos
timestamp 1179386902
<< checkpaint >>
rect -22 -25 134 105
<< ab >>
rect 0 0 112 80
<< pwell >>
rect -4 -7 116 36
<< nwell >>
rect -4 36 116 87
<< polysilicon >>
rect 13 70 15 74
rect 21 70 23 74
rect 29 70 31 74
rect 39 70 41 74
rect 46 70 48 74
rect 53 70 55 74
rect 63 70 65 74
rect 70 70 72 74
rect 77 70 79 74
rect 87 61 89 66
rect 94 61 96 65
rect 101 61 103 65
rect 13 39 15 42
rect 21 39 23 42
rect 29 39 31 42
rect 39 39 41 42
rect 9 38 15 39
rect 9 34 10 38
rect 14 34 15 38
rect 9 33 15 34
rect 19 38 25 39
rect 19 34 20 38
rect 24 34 25 38
rect 19 33 25 34
rect 29 38 41 39
rect 29 34 36 38
rect 40 34 41 38
rect 29 33 41 34
rect 9 30 11 33
rect 21 30 23 33
rect 31 30 33 33
rect 9 6 11 11
rect 46 23 48 42
rect 53 39 55 42
rect 63 39 65 42
rect 53 38 65 39
rect 53 37 60 38
rect 59 34 60 37
rect 64 34 65 38
rect 59 33 65 34
rect 70 23 72 42
rect 77 39 79 42
rect 87 39 89 42
rect 77 37 89 39
rect 77 30 83 37
rect 77 26 78 30
rect 82 26 83 30
rect 77 25 83 26
rect 94 23 96 42
rect 101 39 103 42
rect 101 38 107 39
rect 101 34 102 38
rect 106 34 107 38
rect 101 33 107 34
rect 46 22 52 23
rect 46 18 47 22
rect 51 18 52 22
rect 46 17 52 18
rect 66 22 72 23
rect 66 18 67 22
rect 71 18 72 22
rect 66 17 72 18
rect 89 22 96 23
rect 89 18 90 22
rect 94 18 96 22
rect 89 17 96 18
rect 21 6 23 11
rect 31 6 33 11
<< ndiffusion >>
rect 2 29 9 30
rect 2 25 3 29
rect 7 25 9 29
rect 2 22 9 25
rect 2 18 3 22
rect 7 18 9 22
rect 2 17 9 18
rect 4 11 9 17
rect 11 12 21 30
rect 11 11 14 12
rect 13 8 14 11
rect 18 11 21 12
rect 23 22 31 30
rect 23 18 25 22
rect 29 18 31 22
rect 23 11 31 18
rect 33 23 41 30
rect 33 19 35 23
rect 39 19 41 23
rect 33 16 41 19
rect 33 12 35 16
rect 39 12 41 16
rect 33 11 41 12
rect 18 8 19 11
rect 13 7 19 8
<< pdiffusion >>
rect 5 69 13 70
rect 5 65 7 69
rect 11 65 13 69
rect 5 62 13 65
rect 5 58 7 62
rect 11 58 13 62
rect 5 42 13 58
rect 15 42 21 70
rect 23 42 29 70
rect 31 62 39 70
rect 31 58 33 62
rect 37 58 39 62
rect 31 54 39 58
rect 31 50 33 54
rect 37 50 39 54
rect 31 42 39 50
rect 41 42 46 70
rect 48 42 53 70
rect 55 69 63 70
rect 55 65 57 69
rect 61 65 63 69
rect 55 62 63 65
rect 55 58 57 62
rect 61 58 63 62
rect 55 42 63 58
rect 65 42 70 70
rect 72 42 77 70
rect 79 61 84 70
rect 79 54 87 61
rect 79 50 81 54
rect 85 50 87 54
rect 79 47 87 50
rect 79 43 81 47
rect 85 43 87 47
rect 79 42 87 43
rect 89 42 94 61
rect 96 42 101 61
rect 103 60 110 61
rect 103 56 105 60
rect 109 56 110 60
rect 103 53 110 56
rect 103 49 105 53
rect 109 49 110 53
rect 103 42 110 49
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect -2 69 114 78
rect -2 68 7 69
rect 6 65 7 68
rect 11 68 57 69
rect 11 65 12 68
rect 6 62 12 65
rect 56 65 57 68
rect 61 68 114 69
rect 61 65 62 68
rect 6 58 7 62
rect 11 58 12 62
rect 33 62 38 63
rect 37 58 38 62
rect 56 62 62 65
rect 56 58 57 62
rect 61 58 62 62
rect 104 60 110 68
rect 33 54 38 58
rect 104 56 105 60
rect 109 56 110 60
rect 2 50 33 54
rect 37 50 81 54
rect 85 50 87 54
rect 2 29 6 50
rect 81 47 87 50
rect 104 53 110 56
rect 104 49 105 53
rect 109 49 110 53
rect 10 42 63 46
rect 85 46 87 47
rect 85 43 95 46
rect 81 42 95 43
rect 10 38 14 42
rect 59 38 63 42
rect 19 34 20 38
rect 24 34 31 38
rect 35 34 36 38
rect 40 34 55 38
rect 59 34 60 38
rect 64 34 102 38
rect 106 34 107 38
rect 10 33 14 34
rect 25 30 31 34
rect 51 30 55 34
rect 2 25 3 29
rect 7 25 8 29
rect 25 26 47 30
rect 51 26 78 30
rect 82 26 87 30
rect 2 22 8 25
rect 2 18 3 22
rect 7 18 25 22
rect 29 18 31 22
rect 34 19 35 23
rect 39 19 40 23
rect 34 16 40 19
rect 43 18 47 26
rect 51 18 67 22
rect 71 18 90 22
rect 94 18 95 22
rect 34 12 35 16
rect 39 12 40 16
rect -2 8 14 12
rect 18 8 114 12
rect -2 2 114 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
<< ntransistor >>
rect 9 11 11 30
rect 21 11 23 30
rect 31 11 33 30
<< ptransistor >>
rect 13 42 15 70
rect 21 42 23 70
rect 29 42 31 70
rect 39 42 41 70
rect 46 42 48 70
rect 53 42 55 70
rect 63 42 65 70
rect 70 42 72 70
rect 77 42 79 70
rect 87 42 89 61
rect 94 42 96 61
rect 101 42 103 61
<< polycontact >>
rect 10 34 14 38
rect 20 34 24 38
rect 36 34 40 38
rect 60 34 64 38
rect 78 26 82 30
rect 102 34 106 38
rect 47 18 51 22
rect 67 18 71 22
rect 90 18 94 22
<< ndcontact >>
rect 3 25 7 29
rect 3 18 7 22
rect 14 8 18 12
rect 25 18 29 22
rect 35 19 39 23
rect 35 12 39 16
<< pdcontact >>
rect 7 65 11 69
rect 7 58 11 62
rect 33 58 37 62
rect 33 50 37 54
rect 57 65 61 69
rect 57 58 61 62
rect 81 50 85 54
rect 81 43 85 47
rect 105 56 109 60
rect 105 49 109 53
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
rect 90 -2 94 2
rect 98 -2 102 2
rect 106 -2 110 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
rect 90 78 94 82
rect 98 78 102 82
rect 106 78 110 82
<< psubstratepdiff >>
rect 0 2 112 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 112 2
rect 0 -3 112 -2
<< nsubstratendiff >>
rect 0 82 112 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 112 82
rect 0 77 112 78
<< labels >>
rlabel metal1 12 20 12 20 6 z
rlabel polycontact 12 36 12 36 6 a
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 52 12 52 6 z
rlabel metal1 20 20 20 20 6 z
rlabel ndcontact 28 20 28 20 6 z
rlabel metal1 28 32 28 32 6 b
rlabel metal1 28 44 28 44 6 a
rlabel metal1 20 44 20 44 6 a
rlabel metal1 20 52 20 52 6 z
rlabel metal1 28 52 28 52 6 z
rlabel metal1 52 20 52 20 6 b
rlabel metal1 44 28 44 28 6 b
rlabel metal1 36 28 36 28 6 b
rlabel metal1 52 36 52 36 6 c
rlabel metal1 44 36 44 36 6 c
rlabel metal1 44 44 44 44 6 a
rlabel metal1 52 44 52 44 6 a
rlabel metal1 36 44 36 44 6 a
rlabel metal1 44 52 44 52 6 z
rlabel metal1 52 52 52 52 6 z
rlabel metal1 36 56 36 56 6 z
rlabel metal1 56 6 56 6 6 vss
rlabel polycontact 68 20 68 20 6 b
rlabel metal1 60 20 60 20 6 b
rlabel metal1 60 28 60 28 6 c
rlabel metal1 68 28 68 28 6 c
rlabel metal1 68 36 68 36 6 a
rlabel metal1 60 44 60 44 6 a
rlabel metal1 68 52 68 52 6 z
rlabel metal1 60 52 60 52 6 z
rlabel metal1 56 74 56 74 6 vdd
rlabel metal1 76 20 76 20 6 b
rlabel polycontact 92 20 92 20 6 b
rlabel metal1 84 20 84 20 6 b
rlabel metal1 84 28 84 28 6 c
rlabel metal1 76 28 76 28 6 c
rlabel metal1 76 36 76 36 6 a
rlabel metal1 92 36 92 36 6 a
rlabel metal1 84 36 84 36 6 a
rlabel metal1 92 44 92 44 6 z
rlabel metal1 76 52 76 52 6 z
rlabel metal1 84 48 84 48 6 z
rlabel metal1 100 36 100 36 6 a
<< end >>
