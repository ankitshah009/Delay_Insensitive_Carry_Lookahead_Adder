.subckt a2_x2 i0 i1 q vdd vss
*   SPICE3 file   created from a2_x2.ext -      technology: scmos
m00 w1     i0     vdd    vdd p w=20u  l=2.3636u ad=101.5p   pd=31u      as=140.253p ps=42.5316u
m01 vdd    i1     w1     vdd p w=20u  l=2.3636u ad=140.253p pd=42.5316u as=101.5p   ps=31u
m02 q      w1     vdd    vdd p w=39u  l=2.3636u ad=312p     pd=94u      as=273.494p ps=82.9367u
m03 w2     i0     w1     vss n w=20u  l=2.3636u ad=128.421p pd=40u      as=160p     ps=56u
m04 vss    i1     w2     vss n w=18u  l=2.3636u ad=90p      pd=28.2162u as=115.579p ps=36u
m05 q      w1     vss    vss n w=19u  l=2.3636u ad=152p     pd=54u      as=95p      ps=29.7838u
C0  q      i1     0.334f
C1  q      vdd    0.070f
C2  i1     i0     0.109f
C3  w2     w1     0.034f
C4  i0     vdd    0.021f
C5  i1     w1     0.424f
C6  vdd    w1     0.056f
C7  vss    q      0.055f
C8  vss    i0     0.011f
C9  vss    w1     0.098f
C10 q      i0     0.054f
C11 i1     vdd    0.095f
C12 q      w1     0.115f
C13 i0     w1     0.349f
C14 vss    w2     0.015f
C15 vss    i1     0.054f
C17 q      vss    0.015f
C18 i1     vss    0.039f
C19 i0     vss    0.030f
C21 w1     vss    0.041f
.ends
