magic
tech scmos
timestamp 1179385749
<< checkpaint >>
rect -22 -22 190 94
<< ab >>
rect 0 0 168 72
<< pwell >>
rect -4 -4 172 32
<< nwell >>
rect -4 32 172 76
<< polysilicon >>
rect 9 66 11 70
rect 19 66 21 70
rect 29 66 31 70
rect 39 66 41 70
rect 49 66 51 70
rect 59 66 61 70
rect 69 66 71 70
rect 76 66 78 70
rect 89 66 91 70
rect 96 66 98 70
rect 106 66 108 70
rect 113 66 115 70
rect 125 66 127 70
rect 135 66 137 70
rect 145 66 147 70
rect 9 33 11 38
rect 19 33 21 38
rect 29 33 31 38
rect 9 31 31 33
rect 9 26 11 31
rect 19 26 21 31
rect 29 26 31 31
rect 39 35 41 38
rect 49 35 51 38
rect 59 35 61 38
rect 69 35 71 38
rect 76 35 78 38
rect 89 35 91 38
rect 39 34 61 35
rect 39 33 56 34
rect 39 26 41 33
rect 49 30 56 33
rect 60 30 61 34
rect 49 29 61 30
rect 66 34 72 35
rect 66 30 67 34
rect 71 30 72 34
rect 66 29 72 30
rect 76 34 91 35
rect 76 30 82 34
rect 86 30 91 34
rect 76 29 91 30
rect 49 26 51 29
rect 59 26 61 29
rect 69 26 71 29
rect 76 26 78 29
rect 89 26 91 29
rect 96 35 98 38
rect 106 35 108 38
rect 96 34 108 35
rect 96 30 97 34
rect 101 30 108 34
rect 96 29 108 30
rect 96 26 98 29
rect 106 26 108 29
rect 113 35 115 38
rect 125 35 127 38
rect 135 35 137 38
rect 145 35 147 38
rect 113 34 147 35
rect 113 30 114 34
rect 118 33 147 34
rect 118 30 128 33
rect 113 29 128 30
rect 113 26 115 29
rect 126 26 128 29
rect 136 26 138 33
rect 9 7 11 12
rect 19 7 21 12
rect 29 4 31 12
rect 39 8 41 12
rect 49 8 51 12
rect 59 8 61 12
rect 69 4 71 12
rect 76 7 78 12
rect 29 2 71 4
rect 89 7 91 12
rect 96 7 98 12
rect 106 7 108 12
rect 113 7 115 12
rect 126 2 128 6
rect 136 2 138 6
<< ndiffusion >>
rect 2 24 9 26
rect 2 20 3 24
rect 7 20 9 24
rect 2 17 9 20
rect 2 13 3 17
rect 7 13 9 17
rect 2 12 9 13
rect 11 25 19 26
rect 11 21 13 25
rect 17 21 19 25
rect 11 18 19 21
rect 11 14 13 18
rect 17 14 19 18
rect 11 12 19 14
rect 21 17 29 26
rect 21 13 23 17
rect 27 13 29 17
rect 21 12 29 13
rect 31 25 39 26
rect 31 21 33 25
rect 37 21 39 25
rect 31 18 39 21
rect 31 14 33 18
rect 37 14 39 18
rect 31 12 39 14
rect 41 25 49 26
rect 41 21 43 25
rect 47 21 49 25
rect 41 12 49 21
rect 51 18 59 26
rect 51 14 53 18
rect 57 14 59 18
rect 51 12 59 14
rect 61 25 69 26
rect 61 21 63 25
rect 67 21 69 25
rect 61 12 69 21
rect 71 12 76 26
rect 78 12 89 26
rect 91 12 96 26
rect 98 25 106 26
rect 98 21 100 25
rect 104 21 106 25
rect 98 12 106 21
rect 108 12 113 26
rect 115 12 126 26
rect 80 8 87 12
rect 80 4 81 8
rect 85 4 87 8
rect 117 11 126 12
rect 117 7 118 11
rect 122 7 126 11
rect 117 6 126 7
rect 128 25 136 26
rect 128 21 130 25
rect 134 21 136 25
rect 128 18 136 21
rect 128 14 130 18
rect 134 14 136 18
rect 128 6 136 14
rect 138 19 146 26
rect 138 15 140 19
rect 144 15 146 19
rect 138 11 146 15
rect 138 7 140 11
rect 144 7 146 11
rect 138 6 146 7
rect 80 3 87 4
<< pdiffusion >>
rect 2 65 9 66
rect 2 61 3 65
rect 7 61 9 65
rect 2 58 9 61
rect 2 54 3 58
rect 7 54 9 58
rect 2 51 9 54
rect 2 47 3 51
rect 7 47 9 51
rect 2 38 9 47
rect 11 58 19 66
rect 11 54 13 58
rect 17 54 19 58
rect 11 51 19 54
rect 11 47 13 51
rect 17 47 19 51
rect 11 38 19 47
rect 21 65 29 66
rect 21 61 23 65
rect 27 61 29 65
rect 21 58 29 61
rect 21 54 23 58
rect 27 54 29 58
rect 21 38 29 54
rect 31 58 39 66
rect 31 54 33 58
rect 37 54 39 58
rect 31 51 39 54
rect 31 47 33 51
rect 37 47 39 51
rect 31 38 39 47
rect 41 50 49 66
rect 41 46 43 50
rect 47 46 49 50
rect 41 38 49 46
rect 51 58 59 66
rect 51 54 53 58
rect 57 54 59 58
rect 51 38 59 54
rect 61 50 69 66
rect 61 46 63 50
rect 67 46 69 50
rect 61 38 69 46
rect 71 38 76 66
rect 78 65 89 66
rect 78 61 81 65
rect 85 61 89 65
rect 78 38 89 61
rect 91 38 96 66
rect 98 50 106 66
rect 98 46 100 50
rect 104 46 106 50
rect 98 38 106 46
rect 108 38 113 66
rect 115 65 125 66
rect 115 61 118 65
rect 122 61 125 65
rect 115 38 125 61
rect 127 58 135 66
rect 127 54 129 58
rect 133 54 135 58
rect 127 51 135 54
rect 127 47 129 51
rect 133 47 135 51
rect 127 38 135 47
rect 137 65 145 66
rect 137 61 139 65
rect 143 61 145 65
rect 137 58 145 61
rect 137 54 139 58
rect 143 54 145 58
rect 137 38 145 54
rect 147 51 152 66
rect 147 50 154 51
rect 147 46 149 50
rect 153 46 154 50
rect 147 43 154 46
rect 147 39 149 43
rect 153 39 154 43
rect 147 38 154 39
<< metal1 >>
rect -2 68 170 72
rect -2 65 157 68
rect -2 64 3 65
rect 7 64 23 65
rect 3 58 7 61
rect 22 61 23 64
rect 27 64 81 65
rect 27 61 28 64
rect 80 61 81 64
rect 85 64 118 65
rect 85 61 86 64
rect 117 61 118 64
rect 122 64 139 65
rect 122 61 123 64
rect 138 61 139 64
rect 143 64 157 65
rect 161 64 170 68
rect 143 61 144 64
rect 3 51 7 54
rect 3 46 7 47
rect 13 58 17 59
rect 22 58 28 61
rect 138 58 144 61
rect 22 54 23 58
rect 27 54 28 58
rect 32 54 33 58
rect 37 54 53 58
rect 57 54 129 58
rect 133 54 134 58
rect 138 54 139 58
rect 143 54 144 58
rect 157 60 161 64
rect 157 55 161 56
rect 13 51 17 54
rect 32 51 37 54
rect 32 50 33 51
rect 17 47 33 50
rect 129 51 134 54
rect 13 46 37 47
rect 42 46 43 50
rect 47 46 63 50
rect 67 46 100 50
rect 104 46 126 50
rect 133 50 134 51
rect 133 47 149 50
rect 129 46 149 47
rect 153 46 154 50
rect 13 25 37 26
rect 3 24 7 25
rect 3 17 7 20
rect 17 22 33 25
rect 13 18 17 21
rect 32 21 33 22
rect 42 25 46 46
rect 57 35 63 42
rect 81 38 118 42
rect 50 34 63 35
rect 50 30 56 34
rect 60 30 63 34
rect 50 29 63 30
rect 67 34 77 35
rect 71 30 77 34
rect 81 34 87 38
rect 114 34 118 38
rect 81 30 82 34
rect 86 30 87 34
rect 91 30 97 34
rect 101 30 103 34
rect 67 29 77 30
rect 73 26 77 29
rect 91 26 95 30
rect 114 29 118 30
rect 42 21 43 25
rect 47 21 63 25
rect 67 21 68 25
rect 73 22 95 26
rect 122 25 126 46
rect 148 43 154 46
rect 148 39 149 43
rect 153 39 154 43
rect 99 21 100 25
rect 104 21 126 25
rect 130 25 135 26
rect 134 21 135 25
rect 32 18 37 21
rect 130 18 135 21
rect 13 13 17 14
rect 23 17 27 18
rect 32 14 33 18
rect 37 14 53 18
rect 57 14 130 18
rect 134 14 135 18
rect 140 19 144 20
rect 3 8 7 13
rect 23 8 27 13
rect 140 11 144 15
rect 117 8 118 11
rect -2 4 81 8
rect 85 7 118 8
rect 122 8 123 11
rect 122 7 140 8
rect 154 16 158 17
rect 154 8 158 12
rect 144 7 154 8
rect 85 4 154 7
rect 158 4 170 8
rect -2 0 170 4
<< ntransistor >>
rect 9 12 11 26
rect 19 12 21 26
rect 29 12 31 26
rect 39 12 41 26
rect 49 12 51 26
rect 59 12 61 26
rect 69 12 71 26
rect 76 12 78 26
rect 89 12 91 26
rect 96 12 98 26
rect 106 12 108 26
rect 113 12 115 26
rect 126 6 128 26
rect 136 6 138 26
<< ptransistor >>
rect 9 38 11 66
rect 19 38 21 66
rect 29 38 31 66
rect 39 38 41 66
rect 49 38 51 66
rect 59 38 61 66
rect 69 38 71 66
rect 76 38 78 66
rect 89 38 91 66
rect 96 38 98 66
rect 106 38 108 66
rect 113 38 115 66
rect 125 38 127 66
rect 135 38 137 66
rect 145 38 147 66
<< polycontact >>
rect 56 30 60 34
rect 67 30 71 34
rect 82 30 86 34
rect 97 30 101 34
rect 114 30 118 34
<< ndcontact >>
rect 3 20 7 24
rect 3 13 7 17
rect 13 21 17 25
rect 13 14 17 18
rect 23 13 27 17
rect 33 21 37 25
rect 33 14 37 18
rect 43 21 47 25
rect 53 14 57 18
rect 63 21 67 25
rect 100 21 104 25
rect 81 4 85 8
rect 118 7 122 11
rect 130 21 134 25
rect 130 14 134 18
rect 140 15 144 19
rect 140 7 144 11
<< pdcontact >>
rect 3 61 7 65
rect 3 54 7 58
rect 3 47 7 51
rect 13 54 17 58
rect 13 47 17 51
rect 23 61 27 65
rect 23 54 27 58
rect 33 54 37 58
rect 33 47 37 51
rect 43 46 47 50
rect 53 54 57 58
rect 63 46 67 50
rect 81 61 85 65
rect 100 46 104 50
rect 118 61 122 65
rect 129 54 133 58
rect 129 47 133 51
rect 139 61 143 65
rect 139 54 143 58
rect 149 46 153 50
rect 149 39 153 43
<< psubstratepcontact >>
rect 154 12 158 16
rect 154 4 158 8
<< nsubstratencontact >>
rect 157 64 161 68
rect 157 56 161 60
<< psubstratepdiff >>
rect 153 16 159 24
rect 153 12 154 16
rect 158 12 159 16
rect 153 8 159 12
rect 153 4 154 8
rect 158 4 159 8
rect 153 3 159 4
<< nsubstratendiff >>
rect 156 68 162 69
rect 156 64 157 68
rect 161 64 162 68
rect 156 60 162 64
rect 156 56 157 60
rect 161 56 162 60
rect 156 55 162 56
<< labels >>
rlabel metal1 15 19 15 19 6 n3
rlabel metal1 15 52 15 52 6 n1
rlabel metal1 34 20 34 20 6 n3
rlabel metal1 44 32 44 32 6 z
rlabel metal1 52 32 52 32 6 c
rlabel metal1 60 36 60 36 6 c
rlabel metal1 52 48 52 48 6 z
rlabel metal1 60 48 60 48 6 z
rlabel metal1 34 52 34 52 6 n1
rlabel metal1 84 4 84 4 6 vss
rlabel metal1 76 24 76 24 6 b
rlabel metal1 84 24 84 24 6 b
rlabel metal1 92 24 92 24 6 b
rlabel metal1 92 40 92 40 6 a
rlabel metal1 84 36 84 36 6 a
rlabel metal1 68 48 68 48 6 z
rlabel metal1 76 48 76 48 6 z
rlabel metal1 84 48 84 48 6 z
rlabel metal1 92 48 92 48 6 z
rlabel metal1 84 68 84 68 6 vdd
rlabel polycontact 116 32 116 32 6 a
rlabel metal1 124 32 124 32 6 z
rlabel polycontact 100 32 100 32 6 b
rlabel metal1 100 40 100 40 6 a
rlabel metal1 108 40 108 40 6 a
rlabel metal1 100 48 100 48 6 z
rlabel metal1 108 48 108 48 6 z
rlabel metal1 116 48 116 48 6 z
rlabel metal1 131 52 131 52 6 n1
rlabel metal1 83 56 83 56 6 n1
rlabel metal1 132 20 132 20 6 n3
rlabel metal1 83 16 83 16 6 n3
rlabel metal1 151 44 151 44 6 n1
<< end >>
