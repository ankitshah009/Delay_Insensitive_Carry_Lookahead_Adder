.subckt cgi2cv0x1 a b c vdd vss z
*   SPICE3 file   created from cgi2cv0x1.ext -      technology: scmos
m00 vdd    a      n1     vdd p w=27u  l=2.3636u ad=121.5p   pd=36u      as=125.667p ps=46u
m01 w1     a      vdd    vdd p w=27u  l=2.3636u ad=67.5p    pd=32u      as=121.5p   ps=36u
m02 z      b      w1     vdd p w=27u  l=2.3636u ad=108p     pd=35u      as=67.5p    ps=32u
m03 n1     w2     z      vdd p w=27u  l=2.3636u ad=125.667p pd=46u      as=108p     ps=35u
m04 vdd    b      n1     vdd p w=27u  l=2.3636u ad=121.5p   pd=36u      as=125.667p ps=46u
m05 w2     c      vdd    vdd p w=27u  l=2.3636u ad=161p     pd=68u      as=121.5p   ps=36u
m06 vss    a      n3     vss n w=12u  l=2.3636u ad=73.5p    pd=27u      as=56p      ps=26u
m07 w3     a      vss    vss n w=12u  l=2.3636u ad=30p      pd=17u      as=73.5p    ps=27u
m08 z      b      w3     vss n w=12u  l=2.3636u ad=48p      pd=20u      as=30p      ps=17u
m09 n3     w2     z      vss n w=12u  l=2.3636u ad=56p      pd=26u      as=48p      ps=20u
m10 vss    b      n3     vss n w=12u  l=2.3636u ad=73.5p    pd=27u      as=56p      ps=26u
m11 w2     c      vss    vss n w=12u  l=2.3636u ad=72p      pd=38u      as=73.5p    ps=27u
C0  a      vdd    0.022f
C1  z      w2     0.068f
C2  vss    b      0.032f
C3  n3     a      0.041f
C4  w3     n3     0.006f
C5  n1     w2     0.024f
C6  vss    vdd    0.002f
C7  z      a      0.098f
C8  n3     vss    0.337f
C9  w3     z      0.008f
C10 w1     vdd    0.004f
C11 c      b      0.252f
C12 n1     a      0.042f
C13 vss    z      0.068f
C14 w2     a      0.041f
C15 c      vdd    0.068f
C16 z      w1     0.007f
C17 vss    n1     0.018f
C18 b      vdd    0.032f
C19 w1     n1     0.023f
C20 vss    w2     0.131f
C21 n3     b      0.014f
C22 z      c      0.033f
C23 z      b      0.120f
C24 n3     vdd    0.005f
C25 n1     c      0.008f
C26 vss    a      0.020f
C27 z      vdd    0.062f
C28 c      w2     0.291f
C29 n1     b      0.081f
C30 n3     z      0.177f
C31 c      a      0.010f
C32 w2     b      0.322f
C33 n1     vdd    0.370f
C34 n3     n1     0.038f
C35 b      a      0.126f
C36 w2     vdd    0.044f
C37 n3     w2     0.087f
C38 z      n1     0.191f
C39 vss    c      0.014f
C40 n3     vss    0.003f
C42 z      vss    0.003f
C43 c      vss    0.015f
C44 w2     vss    0.024f
C45 b      vss    0.040f
C46 a      vss    0.042f
.ends
