magic
tech scmos
timestamp 1179385983
<< checkpaint >>
rect -22 -22 94 94
<< ab >>
rect 0 0 72 72
<< pwell >>
rect -4 -4 76 32
<< nwell >>
rect -4 32 76 76
<< polysilicon >>
rect 9 66 11 70
rect 19 66 21 70
rect 29 66 31 70
rect 39 66 41 70
rect 49 66 51 70
rect 59 57 61 61
rect 9 35 11 38
rect 19 35 21 38
rect 29 35 31 38
rect 39 35 41 38
rect 49 35 51 38
rect 59 35 61 38
rect 9 34 42 35
rect 9 33 36 34
rect 20 26 22 33
rect 29 30 36 33
rect 40 30 42 34
rect 29 29 42 30
rect 49 34 61 35
rect 49 30 50 34
rect 54 33 61 34
rect 54 30 55 33
rect 49 29 55 30
rect 30 26 32 29
rect 40 26 42 29
rect 50 26 52 29
rect 20 6 22 11
rect 30 6 32 11
rect 40 5 42 10
rect 50 5 52 10
<< ndiffusion >>
rect 13 24 20 26
rect 13 20 14 24
rect 18 20 20 24
rect 13 16 20 20
rect 13 12 14 16
rect 18 12 20 16
rect 13 11 20 12
rect 22 25 30 26
rect 22 21 24 25
rect 28 21 30 25
rect 22 18 30 21
rect 22 14 24 18
rect 28 14 30 18
rect 22 11 30 14
rect 32 16 40 26
rect 32 12 34 16
rect 38 12 40 16
rect 32 11 40 12
rect 34 10 40 11
rect 42 25 50 26
rect 42 21 44 25
rect 48 21 50 25
rect 42 18 50 21
rect 42 14 44 18
rect 48 14 50 18
rect 42 10 50 14
rect 52 15 59 26
rect 52 11 54 15
rect 58 11 59 15
rect 52 10 59 11
<< pdiffusion >>
rect 2 65 9 66
rect 2 61 3 65
rect 7 61 9 65
rect 2 58 9 61
rect 2 54 3 58
rect 7 54 9 58
rect 2 51 9 54
rect 2 47 3 51
rect 7 47 9 51
rect 2 38 9 47
rect 11 50 19 66
rect 11 46 13 50
rect 17 46 19 50
rect 11 43 19 46
rect 11 39 13 43
rect 17 39 19 43
rect 11 38 19 39
rect 21 65 29 66
rect 21 61 23 65
rect 27 61 29 65
rect 21 57 29 61
rect 21 53 23 57
rect 27 53 29 57
rect 21 38 29 53
rect 31 50 39 66
rect 31 46 33 50
rect 37 46 39 50
rect 31 43 39 46
rect 31 39 33 43
rect 37 39 39 43
rect 31 38 39 39
rect 41 65 49 66
rect 41 61 43 65
rect 47 61 49 65
rect 41 57 49 61
rect 41 53 43 57
rect 47 53 49 57
rect 41 38 49 53
rect 51 57 56 66
rect 51 50 59 57
rect 51 46 53 50
rect 57 46 59 50
rect 51 43 59 46
rect 51 39 53 43
rect 57 39 59 43
rect 51 38 59 39
rect 61 56 68 57
rect 61 52 63 56
rect 67 52 68 56
rect 61 49 68 52
rect 61 45 63 49
rect 67 45 68 49
rect 61 38 68 45
<< metal1 >>
rect -2 68 74 72
rect -2 65 62 68
rect -2 64 3 65
rect 7 64 23 65
rect 3 58 7 61
rect 3 51 7 54
rect 27 64 43 65
rect 23 57 27 61
rect 23 52 27 53
rect 47 64 62 65
rect 66 64 74 68
rect 43 57 47 61
rect 43 52 47 53
rect 62 56 68 64
rect 62 52 63 56
rect 67 52 68 56
rect 3 46 7 47
rect 13 50 17 51
rect 13 43 17 46
rect 9 39 13 42
rect 33 50 38 51
rect 37 46 38 50
rect 33 43 38 46
rect 17 39 33 42
rect 37 42 38 43
rect 53 50 57 51
rect 53 43 57 46
rect 62 49 68 52
rect 62 45 63 49
rect 67 45 68 49
rect 37 39 53 42
rect 57 39 63 42
rect 9 38 63 39
rect 26 26 30 38
rect 35 30 36 34
rect 40 30 50 34
rect 54 30 63 34
rect 23 25 48 26
rect 14 24 18 25
rect 14 16 18 20
rect 23 21 24 25
rect 28 22 44 25
rect 23 18 28 21
rect 23 14 24 18
rect 42 21 44 22
rect 58 21 63 30
rect 42 18 48 21
rect 23 13 28 14
rect 34 16 38 17
rect 14 8 18 12
rect 42 14 44 18
rect 42 13 48 14
rect 54 15 58 16
rect 34 8 38 12
rect 54 8 58 11
rect -2 4 4 8
rect 8 4 64 8
rect 68 4 74 8
rect -2 0 74 4
<< ntransistor >>
rect 20 11 22 26
rect 30 11 32 26
rect 40 10 42 26
rect 50 10 52 26
<< ptransistor >>
rect 9 38 11 66
rect 19 38 21 66
rect 29 38 31 66
rect 39 38 41 66
rect 49 38 51 66
rect 59 38 61 57
<< polycontact >>
rect 36 30 40 34
rect 50 30 54 34
<< ndcontact >>
rect 14 20 18 24
rect 14 12 18 16
rect 24 21 28 25
rect 24 14 28 18
rect 34 12 38 16
rect 44 21 48 25
rect 44 14 48 18
rect 54 11 58 15
<< pdcontact >>
rect 3 61 7 65
rect 3 54 7 58
rect 3 47 7 51
rect 13 46 17 50
rect 13 39 17 43
rect 23 61 27 65
rect 23 53 27 57
rect 33 46 37 50
rect 33 39 37 43
rect 43 61 47 65
rect 43 53 47 57
rect 53 46 57 50
rect 53 39 57 43
rect 63 52 67 56
rect 63 45 67 49
<< psubstratepcontact >>
rect 4 4 8 8
rect 64 4 68 8
<< nsubstratencontact >>
rect 62 64 66 68
<< psubstratepdiff >>
rect 3 8 9 24
rect 3 4 4 8
rect 8 4 9 8
rect 63 8 69 24
rect 3 3 9 4
rect 63 4 64 8
rect 68 4 69 8
rect 63 3 69 4
<< nsubstratendiff >>
rect 61 68 67 69
rect 61 64 62 68
rect 66 64 67 68
rect 61 63 67 64
<< labels >>
rlabel metal1 12 40 12 40 6 z
rlabel metal1 28 32 28 32 6 z
rlabel metal1 20 40 20 40 6 z
rlabel metal1 36 4 36 4 6 vss
rlabel metal1 44 20 44 20 6 z
rlabel metal1 36 24 36 24 6 z
rlabel metal1 44 32 44 32 6 a
rlabel polycontact 52 32 52 32 6 a
rlabel metal1 44 40 44 40 6 z
rlabel metal1 52 40 52 40 6 z
rlabel metal1 36 44 36 44 6 z
rlabel metal1 36 68 36 68 6 vdd
rlabel metal1 60 28 60 28 6 a
rlabel metal1 60 40 60 40 6 z
<< end >>
