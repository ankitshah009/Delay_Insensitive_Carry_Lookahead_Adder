.subckt mxi2v0x2 a0 a1 s vdd vss z
*   SPICE3 file   created from mxi2v0x2.ext -      technology: scmos
m00 w1     a0     vdd    vdd p w=25u  l=2.3636u ad=62.5p    pd=30u      as=149.153p ps=44.9153u
m01 z      s      w1     vdd p w=25u  l=2.3636u ad=100p     pd=33u      as=62.5p    ps=30u
m02 w2     s      z      vdd p w=25u  l=2.3636u ad=62.5p    pd=30u      as=100p     ps=33u
m03 vdd    a0     w2     vdd p w=25u  l=2.3636u ad=149.153p pd=44.9153u as=62.5p    ps=30u
m04 w3     a1     vdd    vdd p w=25u  l=2.3636u ad=62.5p    pd=30u      as=149.153p ps=44.9153u
m05 z      sn     w3     vdd p w=25u  l=2.3636u ad=100p     pd=33u      as=62.5p    ps=30u
m06 w4     sn     z      vdd p w=25u  l=2.3636u ad=62.5p    pd=30u      as=100p     ps=33u
m07 vdd    a1     w4     vdd p w=25u  l=2.3636u ad=149.153p pd=44.9153u as=62.5p    ps=30u
m08 sn     s      vdd    vdd p w=18u  l=2.3636u ad=116p     pd=50u      as=107.39p  ps=32.339u
m09 w5     a0     vss    vss n w=11u  l=2.3636u ad=27.5p    pd=16u      as=78.4528p ps=30.717u
m10 z      sn     w5     vss n w=11u  l=2.3636u ad=44p      pd=19u      as=27.5p    ps=16u
m11 w6     sn     z      vss n w=11u  l=2.3636u ad=27.5p    pd=16u      as=44p      ps=19u
m12 vss    a0     w6     vss n w=11u  l=2.3636u ad=78.4528p pd=30.717u  as=27.5p    ps=16u
m13 w7     a1     vss    vss n w=11u  l=2.3636u ad=27.5p    pd=16u      as=78.4528p ps=30.717u
m14 z      s      w7     vss n w=11u  l=2.3636u ad=44p      pd=19u      as=27.5p    ps=16u
m15 w8     s      z      vss n w=11u  l=2.3636u ad=27.5p    pd=16u      as=44p      ps=19u
m16 vss    a1     w8     vss n w=11u  l=2.3636u ad=78.4528p pd=30.717u  as=27.5p    ps=16u
m17 sn     s      vss    vss n w=9u   l=2.3636u ad=57p      pd=32u      as=64.1887p ps=25.1321u
C0  sn     a0     0.193f
C1  a1     s      0.390f
C2  z      a0     0.288f
C3  w2     vdd    0.005f
C4  w7     a1     0.006f
C5  w6     z      0.010f
C6  a1     vdd    0.042f
C7  s      a0     0.156f
C8  w1     vdd    0.005f
C9  vss    sn     0.107f
C10 vss    z      0.396f
C11 a0     vdd    0.130f
C12 vss    s      0.055f
C13 w3     sn     0.010f
C14 w3     z      0.010f
C15 w3     s      0.004f
C16 z      sn     0.612f
C17 vss    vdd    0.007f
C18 sn     s      0.510f
C19 z      s      0.192f
C20 w3     vdd    0.005f
C21 w8     a1     0.006f
C22 w7     z      0.010f
C23 sn     vdd    0.248f
C24 a1     a0     0.091f
C25 z      vdd    0.340f
C26 w1     a0     0.002f
C27 w5     z      0.013f
C28 s      vdd    0.057f
C29 w4     sn     0.008f
C30 vss    a1     0.135f
C31 w2     sn     0.010f
C32 vss    a0     0.027f
C33 w2     z      0.010f
C34 sn     a1     0.321f
C35 z      a1     0.279f
C36 w1     sn     0.002f
C37 w2     s      0.003f
C38 w4     vdd    0.005f
C39 z      w1     0.018f
C41 z      vss    0.004f
C42 sn     vss    0.047f
C43 a1     vss    0.044f
C44 s      vss    0.072f
C45 a0     vss    0.058f
.ends
