magic
tech scmos
timestamp 1180600794
<< checkpaint >>
rect -22 -22 142 122
<< ab >>
rect 0 0 120 100
<< pwell >>
rect -4 -4 124 48
<< nwell >>
rect -4 48 124 104
<< polysilicon >>
rect 11 94 13 98
rect 23 94 25 98
rect 35 94 37 98
rect 47 94 49 98
rect 79 94 81 98
rect 91 94 93 98
rect 103 94 105 98
rect 11 53 13 56
rect 23 53 25 56
rect 35 53 37 56
rect 47 53 49 56
rect 79 53 81 56
rect 91 53 93 56
rect 11 51 19 53
rect 23 51 29 53
rect 35 52 43 53
rect 35 51 38 52
rect 17 43 19 51
rect 27 43 29 51
rect 37 48 38 51
rect 42 48 43 52
rect 37 47 43 48
rect 47 52 53 53
rect 47 48 48 52
rect 52 48 53 52
rect 47 47 53 48
rect 77 52 83 53
rect 77 48 78 52
rect 82 48 83 52
rect 77 47 83 48
rect 87 52 93 53
rect 87 48 88 52
rect 92 48 93 52
rect 87 47 93 48
rect 17 42 23 43
rect 17 38 18 42
rect 22 38 23 42
rect 17 37 23 38
rect 27 42 33 43
rect 27 38 28 42
rect 32 38 33 42
rect 27 37 33 38
rect 17 29 19 37
rect 27 29 29 37
rect 37 29 39 47
rect 47 29 49 47
rect 15 27 19 29
rect 23 27 29 29
rect 35 27 39 29
rect 43 27 49 29
rect 79 29 81 47
rect 79 27 85 29
rect 15 24 17 27
rect 23 24 25 27
rect 35 24 37 27
rect 43 24 45 27
rect 83 24 85 27
rect 91 24 93 47
rect 103 43 105 55
rect 97 42 105 43
rect 97 38 98 42
rect 102 38 105 42
rect 97 37 105 38
rect 103 25 105 37
rect 15 2 17 6
rect 23 2 25 6
rect 35 2 37 6
rect 43 2 45 6
rect 83 2 85 6
rect 91 2 93 6
rect 103 2 105 6
<< ndiffusion >>
rect 98 24 103 25
rect 7 12 15 24
rect 7 8 8 12
rect 12 8 15 12
rect 7 6 15 8
rect 17 6 23 24
rect 25 22 35 24
rect 25 18 28 22
rect 32 18 35 22
rect 25 6 35 18
rect 37 6 43 24
rect 45 12 53 24
rect 75 22 83 24
rect 75 18 76 22
rect 80 18 83 22
rect 45 8 48 12
rect 52 8 53 12
rect 45 6 53 8
rect 75 6 83 18
rect 85 6 91 24
rect 93 12 103 24
rect 93 8 96 12
rect 100 8 103 12
rect 93 6 103 8
rect 105 22 113 25
rect 105 18 108 22
rect 112 18 113 22
rect 105 6 113 18
<< pdiffusion >>
rect 3 82 11 94
rect 3 78 4 82
rect 8 78 11 82
rect 3 56 11 78
rect 13 72 23 94
rect 13 68 16 72
rect 20 68 23 72
rect 13 56 23 68
rect 25 82 35 94
rect 25 78 28 82
rect 32 78 35 82
rect 25 56 35 78
rect 37 72 47 94
rect 37 68 40 72
rect 44 68 47 72
rect 37 56 47 68
rect 49 82 57 94
rect 49 78 52 82
rect 56 78 57 82
rect 49 56 57 78
rect 71 92 79 94
rect 71 88 72 92
rect 76 88 79 92
rect 71 82 79 88
rect 71 78 72 82
rect 76 78 79 82
rect 71 56 79 78
rect 81 82 91 94
rect 81 78 84 82
rect 88 78 91 82
rect 81 56 91 78
rect 93 92 103 94
rect 93 88 96 92
rect 100 88 103 92
rect 93 82 103 88
rect 93 78 96 82
rect 100 78 103 82
rect 93 72 103 78
rect 93 68 96 72
rect 100 68 103 72
rect 93 56 103 68
rect 98 55 103 56
rect 105 82 113 94
rect 105 78 108 82
rect 112 78 113 82
rect 105 72 113 78
rect 105 68 108 72
rect 112 68 113 72
rect 105 62 113 68
rect 105 58 108 62
rect 112 58 113 62
rect 105 55 113 58
<< metal1 >>
rect -2 92 122 100
rect -2 88 72 92
rect 76 88 96 92
rect 100 88 122 92
rect 72 82 76 88
rect 3 78 4 82
rect 8 78 28 82
rect 32 78 52 82
rect 56 78 57 82
rect 72 77 76 78
rect 84 82 88 83
rect 15 71 16 72
rect 8 68 16 71
rect 20 68 21 72
rect 8 67 20 68
rect 8 22 12 67
rect 18 42 22 63
rect 18 27 22 38
rect 28 42 32 73
rect 84 72 88 78
rect 39 68 40 72
rect 44 68 88 72
rect 96 82 100 88
rect 96 72 100 78
rect 96 67 100 68
rect 108 82 112 83
rect 108 72 112 78
rect 28 27 32 38
rect 38 52 42 63
rect 38 27 42 48
rect 48 52 52 63
rect 48 27 52 48
rect 78 52 82 63
rect 78 27 82 48
rect 88 52 92 63
rect 88 27 92 48
rect 108 62 112 68
rect 98 42 102 43
rect 98 22 102 38
rect 8 18 28 22
rect 32 18 76 22
rect 80 18 102 22
rect 108 22 112 58
rect 108 17 112 18
rect -2 8 8 12
rect 12 8 48 12
rect 52 10 96 12
rect 52 8 62 10
rect -2 6 62 8
rect 66 8 96 10
rect 100 8 122 12
rect 66 6 122 8
rect -2 0 122 6
<< ntransistor >>
rect 15 6 17 24
rect 23 6 25 24
rect 35 6 37 24
rect 43 6 45 24
rect 83 6 85 24
rect 91 6 93 24
rect 103 6 105 25
<< ptransistor >>
rect 11 56 13 94
rect 23 56 25 94
rect 35 56 37 94
rect 47 56 49 94
rect 79 56 81 94
rect 91 56 93 94
rect 103 55 105 94
<< polycontact >>
rect 38 48 42 52
rect 48 48 52 52
rect 78 48 82 52
rect 88 48 92 52
rect 18 38 22 42
rect 28 38 32 42
rect 98 38 102 42
<< ndcontact >>
rect 8 8 12 12
rect 28 18 32 22
rect 76 18 80 22
rect 48 8 52 12
rect 96 8 100 12
rect 108 18 112 22
<< pdcontact >>
rect 4 78 8 82
rect 16 68 20 72
rect 28 78 32 82
rect 40 68 44 72
rect 52 78 56 82
rect 72 88 76 92
rect 72 78 76 82
rect 84 78 88 82
rect 96 88 100 92
rect 96 78 100 82
rect 96 68 100 72
rect 108 78 112 82
rect 108 68 112 72
rect 108 58 112 62
<< psubstratepcontact >>
rect 62 6 66 10
<< psubstratepdiff >>
rect 61 10 67 16
rect 61 6 62 10
rect 66 6 67 10
rect 61 5 67 6
<< labels >>
rlabel metal1 20 45 20 45 6 i5
rlabel metal1 30 50 30 50 6 i4
rlabel metal1 40 45 40 45 6 i3
rlabel metal1 60 6 60 6 6 vss
rlabel metal1 50 45 50 45 6 i2
rlabel metal1 60 94 60 94 6 vdd
rlabel metal1 90 45 90 45 6 i0
rlabel metal1 80 45 80 45 6 i1
rlabel metal1 110 50 110 50 6 q
<< end >>
