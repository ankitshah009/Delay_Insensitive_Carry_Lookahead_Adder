magic
tech scmos
timestamp 1179385373
<< checkpaint >>
rect -22 -25 118 105
<< ab >>
rect 0 0 96 80
<< pwell >>
rect -4 -7 100 36
<< nwell >>
rect -4 36 100 87
<< polysilicon >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 39 70 41 74
rect 49 70 51 74
rect 59 70 61 74
rect 69 70 71 74
rect 79 70 81 74
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 9 38 21 39
rect 9 34 10 38
rect 14 34 21 38
rect 9 33 21 34
rect 25 38 31 39
rect 25 34 26 38
rect 30 35 31 38
rect 39 39 41 42
rect 49 39 51 42
rect 59 39 61 42
rect 69 39 71 42
rect 79 39 81 42
rect 39 38 45 39
rect 30 34 35 35
rect 25 33 35 34
rect 39 34 40 38
rect 44 34 45 38
rect 39 33 45 34
rect 49 38 63 39
rect 49 34 50 38
rect 54 34 58 38
rect 62 34 63 38
rect 49 33 63 34
rect 67 38 73 39
rect 67 34 68 38
rect 72 34 73 38
rect 67 33 73 34
rect 77 38 88 39
rect 77 34 83 38
rect 87 34 88 38
rect 77 33 88 34
rect 9 30 11 33
rect 19 30 21 33
rect 33 30 35 33
rect 41 30 43 33
rect 49 30 51 33
rect 61 30 63 33
rect 69 30 71 33
rect 77 30 79 33
rect 9 17 11 22
rect 19 17 21 22
rect 33 7 35 12
rect 41 7 43 12
rect 49 7 51 12
rect 61 7 63 12
rect 69 7 71 12
rect 77 7 79 12
<< ndiffusion >>
rect 2 27 9 30
rect 2 23 3 27
rect 7 23 9 27
rect 2 22 9 23
rect 11 29 19 30
rect 11 25 13 29
rect 17 25 19 29
rect 11 22 19 25
rect 21 22 33 30
rect 23 12 33 22
rect 35 12 41 30
rect 43 12 49 30
rect 51 22 61 30
rect 51 18 54 22
rect 58 18 61 22
rect 51 12 61 18
rect 63 12 69 30
rect 71 12 77 30
rect 79 17 87 30
rect 79 13 81 17
rect 85 13 87 17
rect 79 12 87 13
rect 23 8 25 12
rect 29 8 31 12
rect 23 7 31 8
<< pdiffusion >>
rect 4 64 9 70
rect 2 63 9 64
rect 2 59 3 63
rect 7 59 9 63
rect 2 58 9 59
rect 4 42 9 58
rect 11 54 19 70
rect 11 50 13 54
rect 17 50 19 54
rect 11 47 19 50
rect 11 43 13 47
rect 17 43 19 47
rect 11 42 19 43
rect 21 62 29 70
rect 21 58 23 62
rect 27 58 29 62
rect 21 55 29 58
rect 21 51 23 55
rect 27 51 29 55
rect 21 42 29 51
rect 31 69 39 70
rect 31 65 33 69
rect 37 65 39 69
rect 31 42 39 65
rect 41 62 49 70
rect 41 58 43 62
rect 47 58 49 62
rect 41 55 49 58
rect 41 51 43 55
rect 47 51 49 55
rect 41 42 49 51
rect 51 69 59 70
rect 51 65 53 69
rect 57 65 59 69
rect 51 62 59 65
rect 51 58 53 62
rect 57 58 59 62
rect 51 42 59 58
rect 61 61 69 70
rect 61 57 63 61
rect 67 57 69 61
rect 61 54 69 57
rect 61 50 63 54
rect 67 50 69 54
rect 61 42 69 50
rect 71 69 79 70
rect 71 65 73 69
rect 77 65 79 69
rect 71 62 79 65
rect 71 58 73 62
rect 77 58 79 62
rect 71 42 79 58
rect 81 55 86 70
rect 81 54 88 55
rect 81 50 83 54
rect 87 50 88 54
rect 81 47 88 50
rect 81 43 83 47
rect 87 43 88 47
rect 81 42 88 43
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect -2 69 98 78
rect -2 68 33 69
rect 37 68 53 69
rect 33 64 37 65
rect 52 65 53 68
rect 57 68 73 69
rect 57 65 58 68
rect 2 59 3 63
rect 7 62 27 63
rect 7 59 23 62
rect 23 55 27 58
rect 2 39 6 55
rect 12 50 13 54
rect 17 50 18 54
rect 43 62 47 63
rect 52 62 58 65
rect 72 65 73 68
rect 77 68 98 69
rect 77 65 78 68
rect 72 62 78 65
rect 52 58 53 62
rect 57 58 58 62
rect 63 61 67 62
rect 43 55 47 58
rect 27 51 43 54
rect 72 58 73 62
rect 77 58 78 62
rect 63 54 67 57
rect 47 51 63 54
rect 23 50 63 51
rect 67 50 83 54
rect 87 50 88 54
rect 12 47 18 50
rect 82 47 88 50
rect 12 43 13 47
rect 17 43 22 47
rect 2 38 14 39
rect 2 34 10 38
rect 2 33 14 34
rect 18 29 22 43
rect 39 42 73 46
rect 82 43 83 47
rect 87 43 88 47
rect 3 27 7 28
rect 12 25 13 29
rect 17 25 22 29
rect 26 38 30 39
rect 39 38 45 42
rect 67 38 73 42
rect 83 38 87 39
rect 39 34 40 38
rect 44 34 45 38
rect 49 34 50 38
rect 54 34 58 38
rect 62 34 63 38
rect 67 34 68 38
rect 72 34 79 38
rect 26 30 30 34
rect 83 30 87 34
rect 26 26 87 30
rect 3 12 7 23
rect 18 22 22 25
rect 18 18 54 22
rect 58 18 59 22
rect 66 17 70 26
rect 81 17 85 18
rect 81 12 85 13
rect -2 8 25 12
rect 29 8 98 12
rect -2 2 98 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
<< ntransistor >>
rect 9 22 11 30
rect 19 22 21 30
rect 33 12 35 30
rect 41 12 43 30
rect 49 12 51 30
rect 61 12 63 30
rect 69 12 71 30
rect 77 12 79 30
<< ptransistor >>
rect 9 42 11 70
rect 19 42 21 70
rect 29 42 31 70
rect 39 42 41 70
rect 49 42 51 70
rect 59 42 61 70
rect 69 42 71 70
rect 79 42 81 70
<< polycontact >>
rect 10 34 14 38
rect 26 34 30 38
rect 40 34 44 38
rect 50 34 54 38
rect 58 34 62 38
rect 68 34 72 38
rect 83 34 87 38
<< ndcontact >>
rect 3 23 7 27
rect 13 25 17 29
rect 54 18 58 22
rect 81 13 85 17
rect 25 8 29 12
<< pdcontact >>
rect 3 59 7 63
rect 13 50 17 54
rect 13 43 17 47
rect 23 58 27 62
rect 23 51 27 55
rect 33 65 37 69
rect 43 58 47 62
rect 43 51 47 55
rect 53 65 57 69
rect 53 58 57 62
rect 63 57 67 61
rect 63 50 67 54
rect 73 65 77 69
rect 73 58 77 62
rect 83 50 87 54
rect 83 43 87 47
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
rect 90 -2 94 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
rect 90 78 94 82
<< psubstratepdiff >>
rect 0 2 96 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 96 2
rect 0 -3 96 -2
<< nsubstratendiff >>
rect 0 82 96 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 96 82
rect 0 77 96 78
<< labels >>
rlabel metal1 4 44 4 44 6 b
rlabel polycontact 12 36 12 36 6 b
rlabel metal1 28 20 28 20 6 z
rlabel metal1 20 36 20 36 6 z
rlabel polycontact 28 36 28 36 6 a1
rlabel metal1 25 56 25 56 6 n3
rlabel metal1 14 61 14 61 6 n3
rlabel metal1 48 6 48 6 6 vss
rlabel metal1 36 20 36 20 6 z
rlabel metal1 36 28 36 28 6 a1
rlabel metal1 44 20 44 20 6 z
rlabel metal1 44 28 44 28 6 a1
rlabel metal1 52 20 52 20 6 z
rlabel metal1 52 28 52 28 6 a1
rlabel metal1 44 44 44 44 6 a2
rlabel polycontact 52 36 52 36 6 a3
rlabel metal1 52 44 52 44 6 a2
rlabel metal1 45 56 45 56 6 n3
rlabel metal1 48 74 48 74 6 vdd
rlabel metal1 60 28 60 28 6 a1
rlabel metal1 68 24 68 24 6 a1
rlabel metal1 76 28 76 28 6 a1
rlabel polycontact 60 36 60 36 6 a3
rlabel metal1 60 44 60 44 6 a2
rlabel metal1 68 44 68 44 6 a2
rlabel metal1 76 36 76 36 6 a2
rlabel metal1 65 56 65 56 6 n3
rlabel metal1 84 28 84 28 6 a1
rlabel metal1 85 48 85 48 6 n3
rlabel metal1 55 52 55 52 6 n3
<< end >>
