magic
tech scmos
timestamp 1185094639
<< checkpaint >>
rect -22 -22 112 122
<< ab >>
rect 0 0 90 100
<< pwell >>
rect -4 -4 94 48
<< nwell >>
rect -4 48 94 104
<< polysilicon >>
rect 15 94 17 98
rect 27 94 29 98
rect 39 94 41 98
rect 51 94 53 98
rect 63 94 65 98
rect 75 94 77 98
rect 15 52 17 55
rect 27 52 29 55
rect 39 52 41 55
rect 51 52 53 55
rect 63 52 65 55
rect 15 51 23 52
rect 15 49 18 51
rect 17 47 18 49
rect 22 47 23 51
rect 27 51 41 52
rect 27 50 36 51
rect 17 46 23 47
rect 35 47 36 50
rect 40 47 41 51
rect 35 46 41 47
rect 47 51 65 52
rect 47 47 48 51
rect 52 50 65 51
rect 52 47 53 50
rect 47 46 53 47
rect 75 48 77 55
rect 75 47 83 48
rect 37 39 39 46
rect 49 39 51 46
rect 75 44 78 47
rect 57 43 78 44
rect 82 43 83 47
rect 57 42 83 43
rect 57 39 59 42
rect 37 12 39 17
rect 49 2 51 6
rect 57 2 59 6
<< ndiffusion >>
rect 28 22 37 39
rect 28 18 30 22
rect 34 18 37 22
rect 28 17 37 18
rect 39 30 49 39
rect 39 26 42 30
rect 46 26 49 30
rect 39 22 49 26
rect 39 18 42 22
rect 46 18 49 22
rect 39 17 49 18
rect 44 6 49 17
rect 51 6 57 39
rect 59 21 68 39
rect 59 17 62 21
rect 66 17 68 21
rect 59 11 68 17
rect 59 7 62 11
rect 66 7 68 11
rect 59 6 68 7
<< pdiffusion >>
rect 6 92 15 94
rect 6 88 8 92
rect 12 88 15 92
rect 6 82 15 88
rect 6 78 8 82
rect 12 78 15 82
rect 6 55 15 78
rect 17 82 27 94
rect 17 78 20 82
rect 24 78 27 82
rect 17 55 27 78
rect 29 72 39 94
rect 29 68 32 72
rect 36 68 39 72
rect 29 55 39 68
rect 41 81 51 94
rect 41 77 44 81
rect 48 77 51 81
rect 41 73 51 77
rect 41 69 44 73
rect 48 69 51 73
rect 41 55 51 69
rect 53 92 63 94
rect 53 88 56 92
rect 60 88 63 92
rect 53 82 63 88
rect 53 78 56 82
rect 60 78 63 82
rect 53 55 63 78
rect 65 81 75 94
rect 65 77 68 81
rect 72 77 75 81
rect 65 73 75 77
rect 65 69 68 73
rect 72 69 75 73
rect 65 55 75 69
rect 77 92 86 94
rect 77 88 80 92
rect 84 88 86 92
rect 77 82 86 88
rect 77 78 80 82
rect 84 78 86 82
rect 77 72 86 78
rect 77 68 80 72
rect 84 68 86 72
rect 77 55 86 68
<< metal1 >>
rect -2 92 92 100
rect -2 88 8 92
rect 12 88 56 92
rect 60 88 80 92
rect 84 88 92 92
rect 8 82 12 88
rect 56 82 60 88
rect 80 82 84 88
rect 19 78 20 82
rect 24 81 48 82
rect 24 78 44 81
rect 8 77 12 78
rect 56 77 60 78
rect 68 81 72 82
rect 44 73 48 77
rect 8 72 37 73
rect 8 68 32 72
rect 36 68 37 72
rect 68 73 72 77
rect 48 69 68 72
rect 44 68 72 69
rect 80 72 84 78
rect 8 32 12 68
rect 80 67 84 68
rect 17 58 83 62
rect 17 51 23 58
rect 17 47 18 51
rect 22 47 23 51
rect 28 51 42 53
rect 28 47 36 51
rect 40 47 42 51
rect 47 51 62 53
rect 47 47 48 51
rect 52 47 62 51
rect 38 37 42 47
rect 8 30 46 32
rect 8 27 42 30
rect 58 27 62 47
rect 77 47 83 58
rect 77 43 78 47
rect 82 43 83 47
rect 77 38 83 43
rect 30 22 34 23
rect 30 12 34 18
rect 42 22 46 26
rect 42 17 46 18
rect 62 21 66 22
rect 62 12 66 17
rect -2 11 92 12
rect -2 8 62 11
rect -2 4 8 8
rect 12 4 18 8
rect 22 7 62 8
rect 66 7 92 11
rect 22 4 92 7
rect -2 0 92 4
<< ntransistor >>
rect 37 17 39 39
rect 49 6 51 39
rect 57 6 59 39
<< ptransistor >>
rect 15 55 17 94
rect 27 55 29 94
rect 39 55 41 94
rect 51 55 53 94
rect 63 55 65 94
rect 75 55 77 94
<< polycontact >>
rect 18 47 22 51
rect 36 47 40 51
rect 48 47 52 51
rect 78 43 82 47
<< ndcontact >>
rect 30 18 34 22
rect 42 26 46 30
rect 42 18 46 22
rect 62 17 66 21
rect 62 7 66 11
<< pdcontact >>
rect 8 88 12 92
rect 8 78 12 82
rect 20 78 24 82
rect 32 68 36 72
rect 44 77 48 81
rect 44 69 48 73
rect 56 88 60 92
rect 56 78 60 82
rect 68 77 72 81
rect 68 69 72 73
rect 80 88 84 92
rect 80 78 84 82
rect 80 68 84 72
<< psubstratepcontact >>
rect 8 4 12 8
rect 18 4 22 8
<< psubstratepdiff >>
rect 7 8 23 9
rect 7 4 8 8
rect 12 4 18 8
rect 22 4 23 8
rect 7 3 23 4
<< labels >>
rlabel metal1 10 50 10 50 6 z
rlabel metal1 20 30 20 30 6 z
rlabel metal1 30 30 30 30 6 z
rlabel metal1 20 55 20 55 6 a1
rlabel metal1 30 50 30 50 6 b
rlabel metal1 30 60 30 60 6 a1
rlabel metal1 20 70 20 70 6 z
rlabel metal1 30 70 30 70 6 z
rlabel metal1 45 6 45 6 6 vss
rlabel metal1 40 30 40 30 6 z
rlabel polycontact 50 50 50 50 6 a2
rlabel metal1 40 45 40 45 6 b
rlabel metal1 40 60 40 60 6 a1
rlabel metal1 50 60 50 60 6 a1
rlabel metal1 46 75 46 75 6 n2
rlabel metal1 33 80 33 80 6 n2
rlabel metal1 45 94 45 94 6 vdd
rlabel metal1 60 40 60 40 6 a2
rlabel metal1 60 60 60 60 6 a1
rlabel metal1 70 60 70 60 6 a1
rlabel metal1 70 75 70 75 6 n2
rlabel metal1 80 50 80 50 6 a1
<< end >>
