.subckt iv1_x05 a vdd vss z
*   SPICE3 file   created from iv1_x05.ext -      technology: scmos
m00 vdd    a      z      vdd p w=12u  l=2.3636u ad=108p     pd=42u      as=78p      ps=40u
m01 vss    a      z      vss n w=6u   l=2.3636u ad=54p      pd=30u      as=48p      ps=28u
C0  z      vdd    0.036f
C1  vss    z      0.093f
C2  z      a      0.162f
C3  a      vdd    0.025f
C4  vss    a      0.011f
C6  z      vss    0.025f
C7  a      vss    0.037f
.ends
