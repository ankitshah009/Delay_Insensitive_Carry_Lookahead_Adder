magic
tech scmos
timestamp 1179386672
<< checkpaint >>
rect -22 -22 70 94
<< ab >>
rect 0 0 48 72
<< pwell >>
rect -4 -4 52 32
<< nwell >>
rect -4 32 52 76
<< polysilicon >>
rect 12 66 14 70
rect 19 66 21 70
rect 33 54 35 59
rect 12 35 14 38
rect 9 34 15 35
rect 9 30 10 34
rect 14 30 15 34
rect 9 29 15 30
rect 11 18 13 29
rect 19 27 21 38
rect 33 35 35 38
rect 29 34 35 35
rect 29 30 30 34
rect 34 30 35 34
rect 29 29 35 30
rect 19 26 25 27
rect 33 26 35 29
rect 19 22 20 26
rect 24 22 25 26
rect 19 21 25 22
rect 21 18 23 21
rect 33 13 35 18
rect 11 4 13 10
rect 21 4 23 10
<< ndiffusion >>
rect 27 18 33 26
rect 35 25 42 26
rect 35 21 37 25
rect 41 21 42 25
rect 35 20 42 21
rect 35 18 40 20
rect 3 10 11 18
rect 13 17 21 18
rect 13 13 15 17
rect 19 13 21 17
rect 13 10 21 13
rect 23 16 31 18
rect 23 12 26 16
rect 30 12 31 16
rect 23 10 31 12
rect 3 8 9 10
rect 3 4 4 8
rect 8 4 9 8
rect 3 3 9 4
<< pdiffusion >>
rect 7 59 12 66
rect 5 58 12 59
rect 5 54 6 58
rect 10 54 12 58
rect 5 51 12 54
rect 5 47 6 51
rect 10 47 12 51
rect 5 46 12 47
rect 7 38 12 46
rect 14 38 19 66
rect 21 64 31 66
rect 21 60 26 64
rect 30 60 31 64
rect 21 54 31 60
rect 21 53 33 54
rect 21 49 26 53
rect 30 49 33 53
rect 21 38 33 49
rect 35 51 40 54
rect 35 50 42 51
rect 35 46 37 50
rect 41 46 42 50
rect 35 43 42 46
rect 35 39 37 43
rect 41 39 42 43
rect 35 38 42 39
<< metal1 >>
rect -2 68 50 72
rect -2 64 36 68
rect 40 64 50 68
rect 6 58 14 59
rect 10 54 14 58
rect 6 53 14 54
rect 26 53 30 60
rect 6 51 11 53
rect 2 18 6 51
rect 10 47 11 51
rect 18 43 22 51
rect 26 48 30 49
rect 37 50 42 51
rect 41 46 42 50
rect 37 43 42 46
rect 10 39 22 43
rect 10 34 14 39
rect 26 35 30 43
rect 41 39 42 43
rect 37 38 42 39
rect 10 29 14 30
rect 18 34 34 35
rect 18 30 30 34
rect 18 29 34 30
rect 19 22 20 26
rect 24 25 25 26
rect 38 25 42 38
rect 24 22 37 25
rect 19 21 37 22
rect 41 21 42 25
rect 2 17 23 18
rect 2 13 15 17
rect 19 13 23 17
rect 26 16 30 17
rect 26 8 30 12
rect -2 4 4 8
rect 8 4 36 8
rect 40 4 50 8
rect -2 0 50 4
<< ntransistor >>
rect 33 18 35 26
rect 11 10 13 18
rect 21 10 23 18
<< ptransistor >>
rect 12 38 14 66
rect 19 38 21 66
rect 33 38 35 54
<< polycontact >>
rect 10 30 14 34
rect 30 30 34 34
rect 20 22 24 26
<< ndcontact >>
rect 37 21 41 25
rect 15 13 19 17
rect 26 12 30 16
rect 4 4 8 8
<< pdcontact >>
rect 6 54 10 58
rect 6 47 10 51
rect 26 60 30 64
rect 26 49 30 53
rect 37 46 41 50
rect 37 39 41 43
<< psubstratepcontact >>
rect 36 4 40 8
<< nsubstratencontact >>
rect 36 64 40 68
<< psubstratepdiff >>
rect 35 8 41 11
rect 35 4 36 8
rect 40 4 41 8
rect 35 3 41 4
<< nsubstratendiff >>
rect 35 68 41 69
rect 35 64 36 68
rect 40 64 41 68
rect 35 61 41 64
<< labels >>
rlabel ntransistor 22 15 22 15 6 an
rlabel metal1 4 32 4 32 6 z
rlabel metal1 20 16 20 16 6 z
rlabel metal1 12 16 12 16 6 z
rlabel metal1 20 32 20 32 6 a
rlabel metal1 12 36 12 36 6 b
rlabel metal1 20 48 20 48 6 b
rlabel metal1 12 56 12 56 6 z
rlabel metal1 24 4 24 4 6 vss
rlabel metal1 28 36 28 36 6 a
rlabel metal1 24 68 24 68 6 vdd
rlabel metal1 30 23 30 23 6 an
rlabel metal1 39 44 39 44 6 an
<< end >>
