.subckt nr3abv0x05 a b c vdd vss z
*   SPICE3 file   created from nr3abv0x05.ext -      technology: scmos
m00 w1     c      z      vdd p w=20u  l=2.3636u ad=50p      pd=25u      as=126p     ps=54u
m01 vdd    nd     w1     vdd p w=20u  l=2.3636u ad=142.727p pd=55.4545u as=50p      ps=25u
m02 nd     a      vdd    vdd p w=12u  l=2.3636u ad=48p      pd=20u      as=85.6364p ps=33.2727u
m03 vdd    b      nd     vdd p w=12u  l=2.3636u ad=85.6364p pd=33.2727u as=48p      ps=20u
m04 z      c      vss    vss n w=6u   l=2.3636u ad=24p      pd=14u      as=47.4545p ps=22.3636u
m05 vss    nd     z      vss n w=6u   l=2.3636u ad=47.4545p pd=22.3636u as=24p      ps=14u
m06 w2     a      vss    vss n w=10u  l=2.3636u ad=25p      pd=15u      as=79.0909p ps=37.2727u
m07 nd     b      w2     vss n w=10u  l=2.3636u ad=62p      pd=34u      as=25p      ps=15u
C0  vss    c      0.016f
C1  a      vdd    0.014f
C2  b      nd     0.212f
C3  z      vdd    0.045f
C4  a      c      0.066f
C5  vdd    nd     0.047f
C6  z      c      0.221f
C7  vss    a      0.069f
C8  nd     c      0.223f
C9  vss    z      0.148f
C10 a      z      0.034f
C11 b      vdd    0.121f
C12 vss    nd     0.051f
C13 b      c      0.036f
C14 w1     vdd    0.004f
C15 a      nd     0.263f
C16 z      nd     0.048f
C17 w1     c      0.009f
C18 vss    b      0.008f
C19 vdd    c      0.065f
C20 b      a      0.085f
C21 b      z      0.021f
C22 vss    vdd    0.002f
C24 b      vss    0.025f
C25 a      vss    0.026f
C26 z      vss    0.014f
C28 nd     vss    0.039f
C29 c      vss    0.025f
.ends
