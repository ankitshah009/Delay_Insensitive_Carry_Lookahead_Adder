magic
tech scmos
timestamp 1179386900
<< checkpaint >>
rect -22 -22 134 94
<< ab >>
rect 0 0 112 72
<< pwell >>
rect -4 -4 116 32
<< nwell >>
rect -4 32 116 76
<< polysilicon >>
rect 13 66 15 70
rect 21 66 23 70
rect 29 66 31 70
rect 39 66 41 70
rect 46 66 48 70
rect 53 66 55 70
rect 63 66 65 70
rect 70 66 72 70
rect 77 66 79 70
rect 87 57 89 62
rect 94 57 96 61
rect 101 57 103 61
rect 13 35 15 38
rect 21 35 23 38
rect 29 35 31 38
rect 39 35 41 38
rect 9 34 15 35
rect 9 30 10 34
rect 14 30 15 34
rect 9 29 15 30
rect 19 34 25 35
rect 19 30 20 34
rect 24 30 25 34
rect 19 29 25 30
rect 29 34 41 35
rect 29 30 36 34
rect 40 30 41 34
rect 29 29 41 30
rect 9 26 11 29
rect 21 26 23 29
rect 31 26 33 29
rect 9 2 11 7
rect 46 19 48 38
rect 53 35 55 38
rect 63 35 65 38
rect 53 34 65 35
rect 53 33 60 34
rect 59 30 60 33
rect 64 30 65 34
rect 59 29 65 30
rect 70 19 72 38
rect 77 35 79 38
rect 87 35 89 38
rect 77 33 89 35
rect 77 26 83 33
rect 77 22 78 26
rect 82 22 83 26
rect 77 21 83 22
rect 94 19 96 38
rect 101 35 103 38
rect 101 34 107 35
rect 101 30 102 34
rect 106 30 107 34
rect 101 29 107 30
rect 46 18 52 19
rect 46 14 47 18
rect 51 14 52 18
rect 46 13 52 14
rect 66 18 72 19
rect 66 14 67 18
rect 71 14 72 18
rect 66 13 72 14
rect 89 18 96 19
rect 89 14 90 18
rect 94 14 96 18
rect 89 13 96 14
rect 21 2 23 7
rect 31 2 33 7
<< ndiffusion >>
rect 2 25 9 26
rect 2 21 3 25
rect 7 21 9 25
rect 2 18 9 21
rect 2 14 3 18
rect 7 14 9 18
rect 2 13 9 14
rect 4 7 9 13
rect 11 8 21 26
rect 11 7 14 8
rect 13 4 14 7
rect 18 7 21 8
rect 23 18 31 26
rect 23 14 25 18
rect 29 14 31 18
rect 23 7 31 14
rect 33 19 41 26
rect 33 15 35 19
rect 39 15 41 19
rect 33 12 41 15
rect 33 8 35 12
rect 39 8 41 12
rect 33 7 41 8
rect 18 4 19 7
rect 13 3 19 4
<< pdiffusion >>
rect 5 65 13 66
rect 5 61 7 65
rect 11 61 13 65
rect 5 58 13 61
rect 5 54 7 58
rect 11 54 13 58
rect 5 38 13 54
rect 15 38 21 66
rect 23 38 29 66
rect 31 58 39 66
rect 31 54 33 58
rect 37 54 39 58
rect 31 50 39 54
rect 31 46 33 50
rect 37 46 39 50
rect 31 38 39 46
rect 41 38 46 66
rect 48 38 53 66
rect 55 65 63 66
rect 55 61 57 65
rect 61 61 63 65
rect 55 58 63 61
rect 55 54 57 58
rect 61 54 63 58
rect 55 38 63 54
rect 65 38 70 66
rect 72 38 77 66
rect 79 57 84 66
rect 79 50 87 57
rect 79 46 81 50
rect 85 46 87 50
rect 79 43 87 46
rect 79 39 81 43
rect 85 39 87 43
rect 79 38 87 39
rect 89 38 94 57
rect 96 38 101 57
rect 103 56 110 57
rect 103 52 105 56
rect 109 52 110 56
rect 103 49 110 52
rect 103 45 105 49
rect 109 45 110 49
rect 103 38 110 45
<< metal1 >>
rect -2 68 114 72
rect -2 65 92 68
rect -2 64 7 65
rect 6 61 7 64
rect 11 64 57 65
rect 11 61 12 64
rect 6 58 12 61
rect 56 61 57 64
rect 61 64 92 65
rect 96 64 104 68
rect 108 64 114 68
rect 61 61 62 64
rect 6 54 7 58
rect 11 54 12 58
rect 33 58 38 59
rect 37 54 38 58
rect 56 58 62 61
rect 56 54 57 58
rect 61 54 62 58
rect 104 56 110 64
rect 33 50 38 54
rect 104 52 105 56
rect 109 52 110 56
rect 2 46 33 50
rect 37 46 81 50
rect 85 46 87 50
rect 2 25 6 46
rect 81 43 87 46
rect 104 49 110 52
rect 104 45 105 49
rect 109 45 110 49
rect 10 38 63 42
rect 85 42 87 43
rect 85 39 95 42
rect 81 38 95 39
rect 10 34 14 38
rect 59 34 63 38
rect 19 30 20 34
rect 24 30 31 34
rect 35 30 36 34
rect 40 30 55 34
rect 59 30 60 34
rect 64 30 102 34
rect 106 30 107 34
rect 10 29 14 30
rect 25 26 31 30
rect 51 26 55 30
rect 2 21 3 25
rect 7 21 8 25
rect 25 22 47 26
rect 51 22 78 26
rect 82 22 87 26
rect 2 18 8 21
rect 2 14 3 18
rect 7 14 25 18
rect 29 14 31 18
rect 34 15 35 19
rect 39 15 40 19
rect 34 12 40 15
rect 43 14 47 22
rect 51 14 67 18
rect 71 14 90 18
rect 94 14 95 18
rect 34 8 35 12
rect 39 8 40 12
rect -2 4 14 8
rect 18 4 48 8
rect 52 4 76 8
rect 80 4 104 8
rect 108 4 114 8
rect -2 0 114 4
<< ntransistor >>
rect 9 7 11 26
rect 21 7 23 26
rect 31 7 33 26
<< ptransistor >>
rect 13 38 15 66
rect 21 38 23 66
rect 29 38 31 66
rect 39 38 41 66
rect 46 38 48 66
rect 53 38 55 66
rect 63 38 65 66
rect 70 38 72 66
rect 77 38 79 66
rect 87 38 89 57
rect 94 38 96 57
rect 101 38 103 57
<< polycontact >>
rect 10 30 14 34
rect 20 30 24 34
rect 36 30 40 34
rect 60 30 64 34
rect 78 22 82 26
rect 102 30 106 34
rect 47 14 51 18
rect 67 14 71 18
rect 90 14 94 18
<< ndcontact >>
rect 3 21 7 25
rect 3 14 7 18
rect 14 4 18 8
rect 25 14 29 18
rect 35 15 39 19
rect 35 8 39 12
<< pdcontact >>
rect 7 61 11 65
rect 7 54 11 58
rect 33 54 37 58
rect 33 46 37 50
rect 57 61 61 65
rect 57 54 61 58
rect 81 46 85 50
rect 81 39 85 43
rect 105 52 109 56
rect 105 45 109 49
<< psubstratepcontact >>
rect 48 4 52 8
rect 76 4 80 8
rect 104 4 108 8
<< nsubstratencontact >>
rect 92 64 96 68
rect 104 64 108 68
<< psubstratepdiff >>
rect 47 8 109 9
rect 47 4 48 8
rect 52 4 76 8
rect 80 4 104 8
rect 108 4 109 8
rect 47 3 109 4
<< nsubstratendiff >>
rect 91 68 109 69
rect 91 64 92 68
rect 96 64 104 68
rect 108 64 109 68
rect 91 63 109 64
<< labels >>
rlabel metal1 12 16 12 16 6 z
rlabel metal1 4 32 4 32 6 z
rlabel polycontact 12 32 12 32 6 a
rlabel metal1 12 48 12 48 6 z
rlabel ndcontact 28 16 28 16 6 z
rlabel metal1 20 16 20 16 6 z
rlabel metal1 36 24 36 24 6 b
rlabel metal1 28 28 28 28 6 b
rlabel metal1 20 40 20 40 6 a
rlabel metal1 36 40 36 40 6 a
rlabel metal1 28 40 28 40 6 a
rlabel metal1 20 48 20 48 6 z
rlabel metal1 36 52 36 52 6 z
rlabel metal1 28 48 28 48 6 z
rlabel metal1 56 4 56 4 6 vss
rlabel metal1 60 16 60 16 6 b
rlabel metal1 52 16 52 16 6 b
rlabel metal1 44 24 44 24 6 b
rlabel metal1 60 24 60 24 6 c
rlabel metal1 52 32 52 32 6 c
rlabel metal1 44 32 44 32 6 c
rlabel metal1 44 40 44 40 6 a
rlabel metal1 60 40 60 40 6 a
rlabel metal1 52 40 52 40 6 a
rlabel metal1 44 48 44 48 6 z
rlabel metal1 60 48 60 48 6 z
rlabel metal1 52 48 52 48 6 z
rlabel metal1 56 68 56 68 6 vdd
rlabel metal1 84 16 84 16 6 b
rlabel metal1 76 16 76 16 6 b
rlabel polycontact 68 16 68 16 6 b
rlabel metal1 68 24 68 24 6 c
rlabel metal1 84 24 84 24 6 c
rlabel metal1 76 24 76 24 6 c
rlabel metal1 84 32 84 32 6 a
rlabel metal1 76 32 76 32 6 a
rlabel metal1 68 32 68 32 6 a
rlabel metal1 84 44 84 44 6 z
rlabel metal1 68 48 68 48 6 z
rlabel metal1 76 48 76 48 6 z
rlabel polycontact 92 16 92 16 6 b
rlabel metal1 100 32 100 32 6 a
rlabel metal1 92 32 92 32 6 a
rlabel metal1 92 40 92 40 6 z
<< end >>
