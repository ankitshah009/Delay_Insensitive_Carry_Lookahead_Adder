magic
tech scmos
timestamp 1185039127
<< checkpaint >>
rect -22 -24 122 124
<< ab >>
rect 0 0 100 100
<< pwell >>
rect -2 -4 102 49
<< nwell >>
rect -2 49 102 104
<< polysilicon >>
rect 35 95 37 98
rect 47 95 49 98
rect 57 95 59 98
rect 81 95 83 98
rect 11 84 13 87
rect 23 84 25 87
rect 11 43 13 55
rect 23 53 25 55
rect 35 53 37 55
rect 21 51 25 53
rect 33 51 37 53
rect 21 43 23 51
rect 33 43 35 51
rect 7 42 13 43
rect 7 38 8 42
rect 12 38 13 42
rect 7 37 13 38
rect 17 42 23 43
rect 17 38 18 42
rect 22 38 23 42
rect 17 37 23 38
rect 27 42 35 43
rect 27 38 28 42
rect 32 38 35 42
rect 47 43 49 55
rect 57 43 59 55
rect 81 53 83 55
rect 75 52 83 53
rect 75 48 76 52
rect 80 48 83 52
rect 75 47 83 48
rect 47 42 53 43
rect 47 39 48 42
rect 27 37 35 38
rect 11 35 13 37
rect 21 35 23 37
rect 33 35 35 37
rect 45 38 48 39
rect 52 38 53 42
rect 45 37 53 38
rect 57 42 63 43
rect 57 38 58 42
rect 62 38 63 42
rect 57 37 63 38
rect 45 35 47 37
rect 57 35 59 37
rect 81 35 83 47
rect 33 20 35 23
rect 45 20 47 23
rect 11 14 13 17
rect 21 14 23 17
rect 57 20 59 23
rect 81 12 83 15
<< ndiffusion >>
rect 3 17 11 35
rect 13 17 21 35
rect 23 23 33 35
rect 35 23 45 35
rect 47 23 57 35
rect 59 23 67 35
rect 23 22 31 23
rect 23 18 26 22
rect 30 18 31 22
rect 37 22 43 23
rect 23 17 31 18
rect 37 18 38 22
rect 42 18 43 22
rect 37 17 43 18
rect 3 12 9 17
rect 3 8 4 12
rect 8 8 9 12
rect 49 12 55 23
rect 61 22 67 23
rect 61 18 62 22
rect 66 18 67 22
rect 61 17 67 18
rect 73 32 81 35
rect 73 28 74 32
rect 78 28 81 32
rect 73 22 81 28
rect 73 18 74 22
rect 78 18 81 22
rect 73 15 81 18
rect 83 32 91 35
rect 83 28 86 32
rect 90 28 91 32
rect 83 22 91 28
rect 83 18 86 22
rect 90 18 91 22
rect 83 15 91 18
rect 3 7 9 8
rect 49 8 50 12
rect 54 8 55 12
rect 49 7 55 8
<< pdiffusion >>
rect 15 92 21 93
rect 15 88 16 92
rect 20 88 21 92
rect 15 84 21 88
rect 28 84 35 95
rect 3 82 11 84
rect 3 78 4 82
rect 8 78 11 82
rect 3 55 11 78
rect 13 55 23 84
rect 25 82 35 84
rect 25 78 28 82
rect 32 78 35 82
rect 25 55 35 78
rect 37 72 47 95
rect 37 68 40 72
rect 44 68 47 72
rect 37 55 47 68
rect 49 55 57 95
rect 59 82 67 95
rect 59 78 62 82
rect 66 78 67 82
rect 59 55 67 78
rect 73 92 81 95
rect 73 88 74 92
rect 78 88 81 92
rect 73 82 81 88
rect 73 78 74 82
rect 78 78 81 82
rect 73 55 81 78
rect 83 82 91 95
rect 83 78 86 82
rect 90 78 91 82
rect 83 72 91 78
rect 83 68 86 72
rect 90 68 91 72
rect 83 62 91 68
rect 83 58 86 62
rect 90 58 91 62
rect 83 55 91 58
<< metal1 >>
rect -2 92 102 101
rect -2 88 16 92
rect 20 88 74 92
rect 78 88 102 92
rect -2 87 102 88
rect 3 82 9 83
rect 27 82 33 83
rect 61 82 67 83
rect 3 78 4 82
rect 8 78 28 82
rect 32 78 62 82
rect 66 78 67 82
rect 3 77 9 78
rect 27 77 33 78
rect 61 77 67 78
rect 73 82 79 87
rect 73 78 74 82
rect 78 78 79 82
rect 73 77 79 78
rect 85 82 91 83
rect 85 78 86 82
rect 90 78 93 82
rect 85 77 93 78
rect 87 73 93 77
rect 39 72 45 73
rect 85 72 93 73
rect 7 42 13 72
rect 7 38 8 42
rect 12 38 13 42
rect 7 18 13 38
rect 17 42 23 72
rect 17 38 18 42
rect 22 38 23 42
rect 17 28 23 38
rect 27 42 33 72
rect 27 38 28 42
rect 32 38 33 42
rect 27 37 33 38
rect 38 68 40 72
rect 44 68 80 72
rect 38 67 45 68
rect 38 32 42 67
rect 28 28 42 32
rect 47 42 53 62
rect 47 38 48 42
rect 52 38 53 42
rect 47 28 53 38
rect 57 42 63 62
rect 76 53 80 68
rect 85 68 86 72
rect 90 68 93 72
rect 85 67 93 68
rect 87 63 93 67
rect 85 62 93 63
rect 85 58 86 62
rect 90 58 93 62
rect 85 57 93 58
rect 75 52 81 53
rect 75 48 76 52
rect 80 48 81 52
rect 75 47 81 48
rect 57 38 58 42
rect 62 38 63 42
rect 57 28 63 38
rect 87 33 93 57
rect 73 32 79 33
rect 73 28 74 32
rect 78 28 79 32
rect 28 23 32 28
rect 25 22 32 23
rect 25 18 26 22
rect 30 18 32 22
rect 37 22 43 23
rect 61 22 67 23
rect 37 18 38 22
rect 42 18 62 22
rect 66 18 67 22
rect 25 17 31 18
rect 37 17 43 18
rect 61 17 67 18
rect 73 22 79 28
rect 85 32 93 33
rect 85 28 86 32
rect 90 28 93 32
rect 85 27 93 28
rect 87 23 93 27
rect 73 18 74 22
rect 78 18 79 22
rect 73 13 79 18
rect 85 22 93 23
rect 85 18 86 22
rect 90 18 93 22
rect 85 17 91 18
rect -2 12 102 13
rect -2 8 4 12
rect 8 10 50 12
rect 8 8 22 10
rect -2 6 22 8
rect 26 6 30 10
rect 34 6 38 10
rect 42 8 50 10
rect 54 8 102 12
rect 42 6 84 8
rect -2 4 84 6
rect 88 4 92 8
rect 96 4 102 8
rect -2 -1 102 4
<< ntransistor >>
rect 11 17 13 35
rect 21 17 23 35
rect 33 23 35 35
rect 45 23 47 35
rect 57 23 59 35
rect 81 15 83 35
<< ptransistor >>
rect 11 55 13 84
rect 23 55 25 84
rect 35 55 37 95
rect 47 55 49 95
rect 57 55 59 95
rect 81 55 83 95
<< polycontact >>
rect 8 38 12 42
rect 18 38 22 42
rect 28 38 32 42
rect 76 48 80 52
rect 48 38 52 42
rect 58 38 62 42
<< ndcontact >>
rect 26 18 30 22
rect 38 18 42 22
rect 4 8 8 12
rect 62 18 66 22
rect 74 28 78 32
rect 74 18 78 22
rect 86 28 90 32
rect 86 18 90 22
rect 50 8 54 12
<< pdcontact >>
rect 16 88 20 92
rect 4 78 8 82
rect 28 78 32 82
rect 40 68 44 72
rect 62 78 66 82
rect 74 88 78 92
rect 74 78 78 82
rect 86 78 90 82
rect 86 68 90 72
rect 86 58 90 62
<< psubstratepcontact >>
rect 22 6 26 10
rect 30 6 34 10
rect 38 6 42 10
rect 84 4 88 8
rect 92 4 96 8
<< psubstratepdiff >>
rect 21 10 43 11
rect 21 6 22 10
rect 26 6 30 10
rect 34 6 38 10
rect 42 6 43 10
rect 83 8 97 9
rect 21 5 43 6
rect 83 4 84 8
rect 88 4 92 8
rect 96 4 97 8
rect 83 3 97 4
<< labels >>
rlabel metal1 10 45 10 45 6 i0
rlabel metal1 10 45 10 45 6 i0
rlabel metal1 20 50 20 50 6 i1
rlabel metal1 20 50 20 50 6 i1
rlabel metal1 30 55 30 55 6 i4
rlabel metal1 30 55 30 55 6 i4
rlabel metal1 50 6 50 6 6 vss
rlabel metal1 50 6 50 6 6 vss
rlabel metal1 50 45 50 45 6 i2
rlabel metal1 50 45 50 45 6 i2
rlabel metal1 50 94 50 94 6 vdd
rlabel metal1 50 94 50 94 6 vdd
rlabel metal1 60 45 60 45 6 i3
rlabel metal1 60 45 60 45 6 i3
rlabel metal1 90 50 90 50 6 q
rlabel metal1 90 50 90 50 6 q
<< end >>
