magic
tech scmos
timestamp 1179387229
<< checkpaint >>
rect -22 -22 94 94
<< ab >>
rect 0 0 72 72
<< pwell >>
rect -4 -4 76 32
<< nwell >>
rect -4 32 76 76
<< polysilicon >>
rect 9 66 11 70
rect 29 68 55 70
rect 22 60 24 65
rect 29 60 31 68
rect 36 60 38 64
rect 46 57 48 62
rect 53 57 55 68
rect 60 57 62 61
rect 9 35 11 38
rect 22 35 24 38
rect 9 34 15 35
rect 9 30 10 34
rect 14 30 15 34
rect 9 29 15 30
rect 19 34 25 35
rect 19 30 20 34
rect 24 30 25 34
rect 19 29 25 30
rect 9 26 11 29
rect 20 18 22 29
rect 29 27 31 38
rect 36 35 38 38
rect 46 35 48 38
rect 36 33 48 35
rect 53 33 55 38
rect 60 35 62 38
rect 60 34 67 35
rect 44 27 48 33
rect 60 30 62 34
rect 66 30 67 34
rect 60 29 67 30
rect 29 26 39 27
rect 29 22 34 26
rect 38 22 39 26
rect 29 21 39 22
rect 44 26 50 27
rect 44 22 45 26
rect 49 22 50 26
rect 44 21 50 22
rect 30 18 32 21
rect 44 18 46 21
rect 9 7 11 12
rect 20 5 22 10
rect 30 5 32 10
rect 44 5 46 10
<< ndiffusion >>
rect 2 25 9 26
rect 2 21 3 25
rect 7 21 9 25
rect 2 18 9 21
rect 2 14 3 18
rect 7 14 9 18
rect 2 12 9 14
rect 11 18 18 26
rect 11 16 20 18
rect 11 12 14 16
rect 18 12 20 16
rect 13 10 20 12
rect 22 17 30 18
rect 22 13 24 17
rect 28 13 30 17
rect 22 10 30 13
rect 32 10 44 18
rect 46 17 53 18
rect 46 13 48 17
rect 52 13 53 17
rect 46 12 53 13
rect 46 10 51 12
rect 34 8 42 10
rect 34 4 36 8
rect 40 4 42 8
rect 34 3 42 4
<< pdiffusion >>
rect 4 51 9 66
rect 2 50 9 51
rect 2 46 3 50
rect 7 46 9 50
rect 2 43 9 46
rect 2 39 3 43
rect 7 39 9 43
rect 2 38 9 39
rect 11 65 20 66
rect 11 61 15 65
rect 19 61 20 65
rect 11 60 20 61
rect 11 58 22 60
rect 11 54 15 58
rect 19 54 22 58
rect 11 38 22 54
rect 24 38 29 60
rect 31 38 36 60
rect 38 57 43 60
rect 38 56 46 57
rect 38 52 40 56
rect 44 52 46 56
rect 38 49 46 52
rect 38 45 40 49
rect 44 45 46 49
rect 38 38 46 45
rect 48 38 53 57
rect 55 38 60 57
rect 62 56 70 57
rect 62 52 64 56
rect 68 52 70 56
rect 62 49 70 52
rect 62 45 64 49
rect 68 45 70 49
rect 62 38 70 45
<< metal1 >>
rect -2 68 74 72
rect -2 65 64 68
rect -2 64 15 65
rect 14 61 15 64
rect 19 64 64 65
rect 68 64 74 68
rect 19 61 20 64
rect 14 58 20 61
rect 14 54 15 58
rect 19 54 20 58
rect 63 56 69 64
rect 39 52 40 56
rect 44 52 45 56
rect 2 50 14 51
rect 2 46 3 50
rect 7 46 14 50
rect 39 49 45 52
rect 2 45 14 46
rect 18 45 40 49
rect 44 45 45 49
rect 63 52 64 56
rect 68 52 69 56
rect 63 49 69 52
rect 63 45 64 49
rect 68 45 69 49
rect 2 43 7 45
rect 2 39 3 43
rect 18 42 22 45
rect 2 38 7 39
rect 10 38 22 42
rect 26 38 63 42
rect 2 26 6 38
rect 10 34 14 38
rect 26 35 30 38
rect 2 25 7 26
rect 2 21 3 25
rect 10 25 14 30
rect 20 34 30 35
rect 57 34 63 38
rect 24 30 30 34
rect 20 29 30 30
rect 34 30 47 34
rect 57 30 62 34
rect 66 30 67 34
rect 34 26 38 30
rect 10 21 27 25
rect 44 22 45 26
rect 49 22 63 26
rect 34 21 38 22
rect 2 18 7 21
rect 2 14 3 18
rect 23 17 27 21
rect 2 13 7 14
rect 13 12 14 16
rect 18 12 19 16
rect 23 13 24 17
rect 28 13 48 17
rect 52 13 53 17
rect 57 14 63 22
rect 13 8 19 12
rect -2 4 36 8
rect 40 4 64 8
rect 68 4 74 8
rect -2 0 74 4
<< ntransistor >>
rect 9 12 11 26
rect 20 10 22 18
rect 30 10 32 18
rect 44 10 46 18
<< ptransistor >>
rect 9 38 11 66
rect 22 38 24 60
rect 29 38 31 60
rect 36 38 38 60
rect 46 38 48 57
rect 53 38 55 57
rect 60 38 62 57
<< polycontact >>
rect 10 30 14 34
rect 20 30 24 34
rect 62 30 66 34
rect 34 22 38 26
rect 45 22 49 26
<< ndcontact >>
rect 3 21 7 25
rect 3 14 7 18
rect 14 12 18 16
rect 24 13 28 17
rect 48 13 52 17
rect 36 4 40 8
<< pdcontact >>
rect 3 46 7 50
rect 3 39 7 43
rect 15 61 19 65
rect 15 54 19 58
rect 40 52 44 56
rect 40 45 44 49
rect 64 52 68 56
rect 64 45 68 49
<< psubstratepcontact >>
rect 64 4 68 8
<< nsubstratencontact >>
rect 64 64 68 68
<< psubstratepdiff >>
rect 63 8 69 24
rect 63 4 64 8
rect 68 4 69 8
rect 63 3 69 4
<< nsubstratendiff >>
rect 63 68 69 69
rect 63 64 64 68
rect 68 64 69 68
rect 63 63 69 64
<< labels >>
rlabel polycontact 12 32 12 32 6 zn
rlabel metal1 4 32 4 32 6 z
rlabel polycontact 12 31 12 31 6 zn
rlabel metal1 12 48 12 48 6 z
rlabel metal1 28 32 28 32 6 a
rlabel metal1 36 4 36 4 6 vss
rlabel metal1 38 15 38 15 6 zn
rlabel polycontact 36 24 36 24 6 b
rlabel metal1 44 32 44 32 6 b
rlabel metal1 52 24 52 24 6 c
rlabel metal1 44 40 44 40 6 a
rlabel metal1 52 40 52 40 6 a
rlabel metal1 36 40 36 40 6 a
rlabel metal1 31 47 31 47 6 zn
rlabel metal1 42 50 42 50 6 zn
rlabel metal1 36 68 36 68 6 vdd
rlabel metal1 60 20 60 20 6 c
rlabel metal1 60 36 60 36 6 a
<< end >>
