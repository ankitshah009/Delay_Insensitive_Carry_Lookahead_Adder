magic
tech scmos
timestamp 1179386549
<< checkpaint >>
rect -22 -25 86 105
<< ab >>
rect 0 0 64 80
<< pwell >>
rect -4 -7 68 36
<< nwell >>
rect -4 36 68 87
<< polysilicon >>
rect 11 70 13 74
rect 21 70 23 74
rect 37 70 39 74
rect 49 70 51 74
rect 11 53 13 56
rect 21 53 23 56
rect 11 52 23 53
rect 11 51 18 52
rect 17 48 18 51
rect 22 48 23 52
rect 17 47 23 48
rect 9 38 15 39
rect 9 34 10 38
rect 14 34 15 38
rect 9 33 15 34
rect 12 30 14 33
rect 19 30 21 47
rect 37 39 39 42
rect 33 38 39 39
rect 33 35 34 38
rect 26 34 34 35
rect 38 34 39 38
rect 49 39 51 42
rect 49 38 55 39
rect 26 33 39 34
rect 26 30 28 33
rect 36 30 38 33
rect 43 30 45 35
rect 49 34 50 38
rect 54 34 55 38
rect 49 33 55 34
rect 50 30 52 33
rect 12 11 14 16
rect 19 8 21 16
rect 26 12 28 16
rect 36 12 38 16
rect 43 8 45 16
rect 50 11 52 16
rect 19 6 45 8
<< ndiffusion >>
rect 2 21 12 30
rect 2 17 3 21
rect 7 17 12 21
rect 2 16 12 17
rect 14 16 19 30
rect 21 16 26 30
rect 28 22 36 30
rect 28 18 30 22
rect 34 18 36 22
rect 28 16 36 18
rect 38 16 43 30
rect 45 16 50 30
rect 52 21 60 30
rect 52 17 54 21
rect 58 17 60 21
rect 52 16 60 17
<< pdiffusion >>
rect 3 69 11 70
rect 3 65 5 69
rect 9 65 11 69
rect 3 56 11 65
rect 13 62 21 70
rect 13 58 15 62
rect 19 58 21 62
rect 13 56 21 58
rect 23 69 37 70
rect 23 65 28 69
rect 32 65 37 69
rect 23 56 37 65
rect 25 42 37 56
rect 39 62 49 70
rect 39 58 42 62
rect 46 58 49 62
rect 39 54 49 58
rect 39 50 42 54
rect 46 50 49 54
rect 39 42 49 50
rect 51 69 59 70
rect 51 65 53 69
rect 57 65 59 69
rect 51 62 59 65
rect 51 58 53 62
rect 57 58 59 62
rect 51 42 59 58
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect -2 69 66 78
rect -2 68 5 69
rect 4 65 5 68
rect 9 68 28 69
rect 9 65 10 68
rect 27 65 28 68
rect 32 68 53 69
rect 32 65 33 68
rect 52 65 53 68
rect 57 68 66 69
rect 57 65 58 68
rect 52 62 58 65
rect 2 58 15 62
rect 19 58 42 62
rect 46 58 47 62
rect 52 58 53 62
rect 57 58 58 62
rect 2 29 6 58
rect 41 54 47 58
rect 17 52 23 54
rect 17 48 18 52
rect 22 48 23 52
rect 41 50 42 54
rect 46 50 47 54
rect 17 46 23 48
rect 17 42 31 46
rect 38 42 47 46
rect 10 38 16 39
rect 14 34 26 38
rect 33 34 34 38
rect 38 34 42 42
rect 49 34 50 38
rect 54 34 55 38
rect 10 33 26 34
rect 22 30 26 33
rect 49 30 55 34
rect 2 25 15 29
rect 22 26 55 30
rect 11 22 15 25
rect 3 21 7 22
rect 11 18 30 22
rect 34 18 35 22
rect 54 21 58 22
rect 3 12 7 17
rect 54 12 58 17
rect -2 2 66 12
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
<< ntransistor >>
rect 12 16 14 30
rect 19 16 21 30
rect 26 16 28 30
rect 36 16 38 30
rect 43 16 45 30
rect 50 16 52 30
<< ptransistor >>
rect 11 56 13 70
rect 21 56 23 70
rect 37 42 39 70
rect 49 42 51 70
<< polycontact >>
rect 18 48 22 52
rect 10 34 14 38
rect 34 34 38 38
rect 50 34 54 38
<< ndcontact >>
rect 3 17 7 21
rect 30 18 34 22
rect 54 17 58 21
<< pdcontact >>
rect 5 65 9 69
rect 15 58 19 62
rect 28 65 32 69
rect 42 58 46 62
rect 42 50 46 54
rect 53 65 57 69
rect 53 58 57 62
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
<< psubstratepdiff >>
rect 0 2 64 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 64 2
rect 0 -3 64 -2
<< nsubstratendiff >>
rect 0 82 64 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 64 82
rect 0 77 64 78
<< labels >>
rlabel metal1 4 40 4 40 6 z
rlabel metal1 20 20 20 20 6 z
rlabel metal1 20 36 20 36 6 a
rlabel metal1 20 48 20 48 6 b
rlabel metal1 12 60 12 60 6 z
rlabel metal1 20 60 20 60 6 z
rlabel metal1 32 6 32 6 6 vss
rlabel metal1 28 20 28 20 6 z
rlabel metal1 28 28 28 28 6 a
rlabel metal1 36 28 36 28 6 a
rlabel metal1 28 44 28 44 6 b
rlabel metal1 28 60 28 60 6 z
rlabel metal1 36 60 36 60 6 z
rlabel metal1 32 74 32 74 6 vdd
rlabel metal1 44 28 44 28 6 a
rlabel metal1 44 44 44 44 6 c
rlabel metal1 44 56 44 56 6 z
rlabel metal1 52 32 52 32 6 a
<< end >>
