.subckt nr3v1x05 a b c vdd vss z
*   SPICE3 file   created from nr3v1x05.ext -      technology: scmos
m00 w1     c      z      vdd p w=28u  l=2.3636u ad=70p      pd=33u      as=166p     ps=70u
m01 w2     b      w1     vdd p w=28u  l=2.3636u ad=70p      pd=33u      as=70p      ps=33u
m02 vdd    a      w2     vdd p w=28u  l=2.3636u ad=280p     pd=76u      as=70p      ps=33u
m03 vss    c      z      vss n w=10u  l=2.3636u ad=70p      pd=32.6667u as=47.3333p ps=23.3333u
m04 z      b      vss    vss n w=10u  l=2.3636u ad=47.3333p pd=23.3333u as=70p      ps=32.6667u
m05 vss    a      z      vss n w=10u  l=2.3636u ad=70p      pd=32.6667u as=47.3333p ps=23.3333u
C0  vdd    a      0.086f
C1  vss    b      0.030f
C2  vdd    c      0.025f
C3  z      b      0.104f
C4  w1     c      0.016f
C5  vss    vdd    0.003f
C6  a      c      0.089f
C7  vdd    w2     0.005f
C8  vdd    z      0.049f
C9  vss    a      0.021f
C10 vss    c      0.014f
C11 w2     a      0.003f
C12 vdd    b      0.015f
C13 z      a      0.031f
C14 w2     c      0.010f
C15 a      b      0.117f
C16 z      c      0.175f
C17 b      c      0.139f
C18 vss    z      0.162f
C19 vdd    w1     0.005f
C22 z      vss    0.014f
C23 a      vss    0.024f
C24 b      vss    0.021f
C25 c      vss    0.015f
.ends
