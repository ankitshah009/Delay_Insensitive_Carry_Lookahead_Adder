magic
tech scmos
timestamp 1180640195
<< checkpaint >>
rect -24 -26 94 126
<< ab >>
rect 0 0 70 100
<< pwell >>
rect -4 -6 74 49
<< nwell >>
rect -4 49 74 106
<< polysilicon >>
rect 13 94 15 98
rect 21 94 23 98
rect 33 94 35 98
rect 45 94 47 98
rect 57 94 59 98
rect 13 48 15 57
rect 21 54 23 57
rect 33 54 35 57
rect 21 52 27 54
rect 33 52 41 54
rect 25 48 27 52
rect 35 51 41 52
rect 13 47 21 48
rect 13 45 16 47
rect 11 43 16 45
rect 20 43 21 47
rect 11 42 21 43
rect 25 47 31 48
rect 25 43 26 47
rect 30 43 31 47
rect 35 47 36 51
rect 40 47 41 51
rect 35 46 41 47
rect 25 42 31 43
rect 45 42 47 57
rect 57 53 59 57
rect 51 52 59 53
rect 51 48 52 52
rect 56 48 59 52
rect 51 47 59 48
rect 11 33 13 42
rect 25 38 27 42
rect 45 41 53 42
rect 45 38 48 41
rect 23 36 27 38
rect 35 37 48 38
rect 52 37 53 41
rect 35 36 53 37
rect 23 33 25 36
rect 35 33 37 36
rect 57 33 59 47
rect 11 12 13 17
rect 23 12 25 17
rect 35 12 37 17
rect 57 12 59 17
<< ndiffusion >>
rect 6 23 11 33
rect 3 22 11 23
rect 3 18 4 22
rect 8 18 11 22
rect 3 17 11 18
rect 13 30 23 33
rect 13 26 16 30
rect 20 26 23 30
rect 13 17 23 26
rect 25 32 35 33
rect 25 28 28 32
rect 32 28 35 32
rect 25 17 35 28
rect 37 17 57 33
rect 59 32 67 33
rect 59 28 62 32
rect 66 28 67 32
rect 59 24 67 28
rect 59 20 62 24
rect 66 20 67 24
rect 59 19 67 20
rect 59 17 64 19
rect 39 12 55 17
rect 39 8 40 12
rect 44 8 50 12
rect 54 8 55 12
rect 39 7 55 8
<< pdiffusion >>
rect 4 92 13 94
rect 4 88 6 92
rect 10 88 13 92
rect 4 57 13 88
rect 15 57 21 94
rect 23 82 33 94
rect 23 78 26 82
rect 30 78 33 82
rect 23 57 33 78
rect 35 82 45 94
rect 35 78 38 82
rect 42 78 45 82
rect 35 74 45 78
rect 35 70 38 74
rect 42 70 45 74
rect 35 57 45 70
rect 47 92 57 94
rect 47 88 50 92
rect 54 88 57 92
rect 47 82 57 88
rect 47 78 50 82
rect 54 78 57 82
rect 47 72 57 78
rect 47 68 50 72
rect 54 68 57 72
rect 47 57 57 68
rect 59 71 64 94
rect 59 70 67 71
rect 59 66 62 70
rect 66 66 67 70
rect 59 62 67 66
rect 59 58 62 62
rect 66 58 67 62
rect 59 57 67 58
<< metal1 >>
rect -2 92 72 100
rect -2 88 6 92
rect 10 88 50 92
rect 54 88 72 92
rect 8 82 33 83
rect 8 78 26 82
rect 30 78 33 82
rect 38 82 42 83
rect 8 30 12 78
rect 38 74 42 78
rect 18 70 38 72
rect 18 68 42 70
rect 50 82 54 88
rect 50 72 54 78
rect 18 48 22 68
rect 50 67 54 68
rect 62 70 66 71
rect 62 62 66 66
rect 16 47 22 48
rect 20 43 22 47
rect 16 42 22 43
rect 26 58 62 62
rect 26 47 30 58
rect 26 42 30 43
rect 36 51 52 52
rect 40 48 52 51
rect 56 48 57 52
rect 40 47 42 48
rect 18 38 22 42
rect 18 34 32 38
rect 36 37 42 47
rect 47 41 53 42
rect 47 37 48 41
rect 52 37 53 41
rect 28 32 32 34
rect 47 32 53 37
rect 8 26 16 30
rect 20 26 21 30
rect 37 28 53 32
rect 62 32 66 58
rect 28 27 32 28
rect 62 24 66 28
rect 3 18 4 22
rect 8 20 62 22
rect 8 18 66 20
rect -2 8 40 12
rect 44 8 50 12
rect 54 8 72 12
rect -2 0 72 8
<< ntransistor >>
rect 11 17 13 33
rect 23 17 25 33
rect 35 17 37 33
rect 57 17 59 33
<< ptransistor >>
rect 13 57 15 94
rect 21 57 23 94
rect 33 57 35 94
rect 45 57 47 94
rect 57 57 59 94
<< polycontact >>
rect 16 43 20 47
rect 26 43 30 47
rect 36 47 40 51
rect 52 48 56 52
rect 48 37 52 41
<< ndcontact >>
rect 4 18 8 22
rect 16 26 20 30
rect 28 28 32 32
rect 62 28 66 32
rect 62 20 66 24
rect 40 8 44 12
rect 50 8 54 12
<< pdcontact >>
rect 6 88 10 92
rect 26 78 30 82
rect 38 78 42 82
rect 38 70 42 74
rect 50 88 54 92
rect 50 78 54 82
rect 50 68 54 72
rect 62 66 66 70
rect 62 58 66 62
<< psubstratepcontact >>
rect 8 4 12 8
rect 18 4 22 8
<< psubstratepdiff >>
rect 7 8 23 9
rect 7 4 8 8
rect 12 4 18 8
rect 22 4 23 8
rect 7 3 23 4
<< labels >>
rlabel polycontact 28 45 28 45 6 bn
rlabel metal1 10 55 10 55 6 z
rlabel metal1 10 55 10 55 6 z
rlabel metal1 30 32 30 32 6 an
rlabel metal1 28 52 28 52 6 bn
rlabel metal1 20 53 20 53 6 an
rlabel metal1 20 80 20 80 6 z
rlabel metal1 20 80 20 80 6 z
rlabel metal1 30 80 30 80 6 z
rlabel metal1 30 80 30 80 6 z
rlabel metal1 35 6 35 6 6 vss
rlabel metal1 35 6 35 6 6 vss
rlabel metal1 50 35 50 35 6 a
rlabel metal1 40 45 40 45 6 b
rlabel metal1 40 30 40 30 6 a
rlabel metal1 40 45 40 45 6 b
rlabel metal1 50 35 50 35 6 a
rlabel metal1 40 30 40 30 6 a
rlabel metal1 50 50 50 50 6 b
rlabel metal1 50 50 50 50 6 b
rlabel metal1 40 75 40 75 6 an
rlabel metal1 35 94 35 94 6 vdd
rlabel metal1 35 94 35 94 6 vdd
rlabel metal1 34 20 34 20 6 bn
rlabel metal1 64 44 64 44 6 bn
<< end >>
