magic
tech scmos
timestamp 1179385216
<< checkpaint >>
rect -22 -25 78 105
<< ab >>
rect 0 0 56 80
<< pwell >>
rect -4 -7 60 36
<< nwell >>
rect -4 36 60 87
<< polysilicon >>
rect 12 70 14 74
rect 19 70 21 74
rect 29 70 31 74
rect 39 70 41 74
rect 12 32 14 43
rect 19 40 21 43
rect 29 40 31 43
rect 39 40 41 43
rect 19 39 25 40
rect 19 35 20 39
rect 24 35 25 39
rect 19 34 25 35
rect 29 39 35 40
rect 29 35 30 39
rect 34 35 35 39
rect 29 34 35 35
rect 39 39 47 40
rect 39 35 42 39
rect 46 35 47 39
rect 39 34 47 35
rect 9 31 15 32
rect 9 27 10 31
rect 14 27 15 31
rect 9 26 15 27
rect 10 23 12 26
rect 20 23 22 34
rect 32 26 34 34
rect 39 26 41 34
rect 10 12 12 17
rect 20 12 22 17
rect 32 12 34 17
rect 39 12 41 17
<< ndiffusion >>
rect 24 23 32 26
rect 2 17 10 23
rect 12 22 20 23
rect 12 18 14 22
rect 18 18 20 22
rect 12 17 20 18
rect 22 17 32 23
rect 34 17 39 26
rect 41 23 46 26
rect 41 22 48 23
rect 41 18 43 22
rect 47 18 48 22
rect 41 17 48 18
rect 2 12 8 17
rect 24 12 30 17
rect 2 8 3 12
rect 7 8 8 12
rect 2 7 8 8
rect 24 8 25 12
rect 29 8 30 12
rect 24 7 30 8
<< pdiffusion >>
rect 7 64 12 70
rect 5 63 12 64
rect 5 59 6 63
rect 10 59 12 63
rect 5 55 12 59
rect 5 51 6 55
rect 10 51 12 55
rect 5 50 12 51
rect 7 43 12 50
rect 14 43 19 70
rect 21 62 29 70
rect 21 58 23 62
rect 27 58 29 62
rect 21 43 29 58
rect 31 69 39 70
rect 31 65 33 69
rect 37 65 39 69
rect 31 43 39 65
rect 41 63 46 70
rect 41 62 48 63
rect 41 58 43 62
rect 47 58 48 62
rect 41 57 48 58
rect 41 43 46 57
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect -2 69 58 78
rect -2 68 33 69
rect 32 65 33 68
rect 37 68 58 69
rect 37 65 38 68
rect 2 22 6 63
rect 10 59 11 63
rect 22 58 23 62
rect 27 58 43 62
rect 47 58 48 62
rect 10 51 11 55
rect 18 49 30 55
rect 34 49 46 55
rect 10 31 14 47
rect 18 41 24 49
rect 20 39 24 41
rect 42 39 46 49
rect 29 35 30 39
rect 34 35 38 39
rect 20 34 24 35
rect 33 30 38 35
rect 42 34 46 35
rect 14 27 23 30
rect 10 26 23 27
rect 33 26 47 30
rect 2 18 14 22
rect 18 18 43 22
rect 47 18 48 22
rect -2 8 3 12
rect 7 8 25 12
rect 29 8 58 12
rect -2 2 58 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
<< ntransistor >>
rect 10 17 12 23
rect 20 17 22 23
rect 32 17 34 26
rect 39 17 41 26
<< ptransistor >>
rect 12 43 14 70
rect 19 43 21 70
rect 29 43 31 70
rect 39 43 41 70
<< polycontact >>
rect 20 35 24 39
rect 30 35 34 39
rect 42 35 46 39
rect 10 27 14 31
<< ndcontact >>
rect 14 18 18 22
rect 43 18 47 22
rect 3 8 7 12
rect 25 8 29 12
<< pdcontact >>
rect 6 59 10 63
rect 6 51 10 55
rect 23 58 27 62
rect 33 65 37 69
rect 43 58 47 62
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
<< psubstratepdiff >>
rect 0 2 56 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 56 2
rect 0 -3 56 -2
<< nsubstratendiff >>
rect 0 82 56 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 56 82
rect 0 77 56 78
<< labels >>
rlabel metal1 4 44 4 44 6 z
rlabel metal1 12 20 12 20 6 z
rlabel metal1 12 40 12 40 6 c
rlabel metal1 28 6 28 6 6 vss
rlabel metal1 20 28 20 28 6 c
rlabel metal1 20 20 20 20 6 z
rlabel metal1 28 20 28 20 6 z
rlabel metal1 28 52 28 52 6 b
rlabel metal1 20 48 20 48 6 b
rlabel metal1 28 74 28 74 6 vdd
rlabel metal1 36 20 36 20 6 z
rlabel metal1 44 28 44 28 6 a1
rlabel ndcontact 44 20 44 20 6 z
rlabel metal1 36 32 36 32 6 a1
rlabel metal1 44 48 44 48 6 a2
rlabel metal1 36 52 36 52 6 a2
rlabel metal1 35 60 35 60 6 n1
<< end >>
