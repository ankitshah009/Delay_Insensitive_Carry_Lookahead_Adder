magic
tech scmos
timestamp 1179386407
<< checkpaint >>
rect -22 -25 78 105
<< ab >>
rect 0 0 56 80
<< pwell >>
rect -4 -7 60 36
<< nwell >>
rect -4 36 60 87
<< polysilicon >>
rect 14 69 16 74
rect 24 69 26 74
rect 35 61 37 66
rect 45 61 47 65
rect 14 39 16 42
rect 24 39 26 42
rect 35 39 37 42
rect 45 39 47 42
rect 9 38 26 39
rect 9 34 10 38
rect 14 34 26 38
rect 9 33 26 34
rect 24 30 26 33
rect 31 38 47 39
rect 31 34 42 38
rect 46 34 47 38
rect 31 33 47 34
rect 31 30 33 33
rect 24 6 26 11
rect 31 6 33 11
<< ndiffusion >>
rect 17 29 24 30
rect 17 25 18 29
rect 22 25 24 29
rect 17 22 24 25
rect 17 18 18 22
rect 22 18 24 22
rect 17 17 24 18
rect 19 11 24 17
rect 26 11 31 30
rect 33 23 41 30
rect 33 19 35 23
rect 39 19 41 23
rect 33 16 41 19
rect 33 12 35 16
rect 39 12 41 16
rect 33 11 41 12
<< pdiffusion >>
rect 6 68 14 69
rect 6 64 8 68
rect 12 64 14 68
rect 6 61 14 64
rect 6 57 8 61
rect 12 57 14 61
rect 6 42 14 57
rect 16 54 24 69
rect 16 50 18 54
rect 22 50 24 54
rect 16 47 24 50
rect 16 43 18 47
rect 22 43 24 47
rect 16 42 24 43
rect 26 68 33 69
rect 26 64 28 68
rect 32 64 33 68
rect 26 61 33 64
rect 26 57 28 61
rect 32 57 35 61
rect 26 42 35 57
rect 37 54 45 61
rect 37 50 39 54
rect 43 50 45 54
rect 37 47 45 50
rect 37 43 39 47
rect 43 43 45 47
rect 37 42 45 43
rect 47 60 54 61
rect 47 56 49 60
rect 53 56 54 60
rect 47 53 54 56
rect 47 49 49 53
rect 53 49 54 53
rect 47 42 54 49
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect -2 68 58 78
rect 8 61 12 64
rect 8 56 12 57
rect 28 61 32 64
rect 28 56 32 57
rect 49 60 53 68
rect 18 54 22 55
rect 18 47 22 50
rect 2 39 6 47
rect 39 54 43 55
rect 39 47 43 50
rect 49 53 53 56
rect 49 48 53 49
rect 22 43 39 46
rect 18 42 43 43
rect 2 38 14 39
rect 2 34 10 38
rect 2 33 14 34
rect 18 29 22 42
rect 41 34 42 38
rect 46 34 54 38
rect 50 25 54 34
rect 18 22 22 25
rect 18 17 22 18
rect 35 23 39 24
rect 35 16 39 19
rect -2 2 58 12
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
<< ntransistor >>
rect 24 11 26 30
rect 31 11 33 30
<< ptransistor >>
rect 14 42 16 69
rect 24 42 26 69
rect 35 42 37 61
rect 45 42 47 61
<< polycontact >>
rect 10 34 14 38
rect 42 34 46 38
<< ndcontact >>
rect 18 25 22 29
rect 18 18 22 22
rect 35 19 39 23
rect 35 12 39 16
<< pdcontact >>
rect 8 64 12 68
rect 8 57 12 61
rect 18 50 22 54
rect 18 43 22 47
rect 28 64 32 68
rect 28 57 32 61
rect 39 50 43 54
rect 39 43 43 47
rect 49 56 53 60
rect 49 49 53 53
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
<< psubstratepdiff >>
rect 0 2 56 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 56 2
rect 0 -3 56 -2
<< nsubstratendiff >>
rect 0 82 56 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 56 82
rect 0 77 56 78
<< labels >>
rlabel metal1 4 40 4 40 6 b
rlabel polycontact 12 36 12 36 6 b
rlabel metal1 20 36 20 36 6 z
rlabel metal1 28 6 28 6 6 vss
rlabel metal1 36 44 36 44 6 z
rlabel metal1 28 44 28 44 6 z
rlabel metal1 28 74 28 74 6 vdd
rlabel polycontact 44 36 44 36 6 a
rlabel metal1 52 28 52 28 6 a
<< end >>
