magic
tech scmos
timestamp 1179387663
<< checkpaint >>
rect -22 -25 182 105
<< ab >>
rect 0 0 160 80
<< pwell >>
rect -4 -7 164 36
<< nwell >>
rect -4 36 164 87
<< polysilicon >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 39 70 41 74
rect 49 70 71 72
rect 49 67 51 70
rect 59 67 61 70
rect 69 67 71 70
rect 79 67 81 72
rect 89 67 91 72
rect 119 67 121 72
rect 129 67 131 72
rect 139 67 141 72
rect 149 67 151 72
rect 99 61 101 65
rect 109 61 111 65
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 39 39 41 42
rect 9 38 41 39
rect 49 38 51 42
rect 59 38 61 42
rect 69 39 71 42
rect 79 39 81 42
rect 89 39 91 42
rect 99 39 101 42
rect 109 39 111 42
rect 119 39 121 42
rect 129 39 131 42
rect 139 39 141 42
rect 149 39 151 42
rect 66 38 72 39
rect 9 34 10 38
rect 14 37 41 38
rect 14 34 32 37
rect 66 34 67 38
rect 71 34 72 38
rect 9 33 32 34
rect 20 30 22 33
rect 30 30 32 33
rect 50 30 52 34
rect 60 30 62 34
rect 66 33 72 34
rect 70 30 72 33
rect 77 38 94 39
rect 77 34 78 38
rect 82 34 85 38
rect 89 34 94 38
rect 77 33 94 34
rect 77 30 79 33
rect 92 30 94 33
rect 99 38 111 39
rect 99 34 100 38
rect 104 34 111 38
rect 99 33 111 34
rect 115 38 121 39
rect 115 34 116 38
rect 120 34 121 38
rect 115 33 121 34
rect 128 38 151 39
rect 128 34 146 38
rect 150 34 151 38
rect 128 33 151 34
rect 99 30 101 33
rect 109 30 111 33
rect 116 30 118 33
rect 128 30 130 33
rect 138 30 140 33
rect 20 6 22 11
rect 30 8 32 11
rect 50 8 52 11
rect 60 8 62 11
rect 30 6 62 8
rect 70 6 72 10
rect 77 6 79 10
rect 92 8 94 16
rect 99 12 101 16
rect 109 12 111 16
rect 116 8 118 16
rect 92 6 118 8
rect 128 6 130 11
rect 138 6 140 11
<< ndiffusion >>
rect 13 24 20 30
rect 13 20 14 24
rect 18 20 20 24
rect 13 16 20 20
rect 13 12 14 16
rect 18 12 20 16
rect 13 11 20 12
rect 22 29 30 30
rect 22 25 24 29
rect 28 25 30 29
rect 22 22 30 25
rect 22 18 24 22
rect 28 18 30 22
rect 22 11 30 18
rect 32 24 39 30
rect 32 20 34 24
rect 38 20 39 24
rect 45 23 50 30
rect 32 16 39 20
rect 43 22 50 23
rect 43 18 44 22
rect 48 18 50 22
rect 43 17 50 18
rect 32 12 34 16
rect 38 12 39 16
rect 32 11 39 12
rect 45 11 50 17
rect 52 29 60 30
rect 52 25 54 29
rect 58 25 60 29
rect 52 11 60 25
rect 62 22 70 30
rect 62 18 64 22
rect 68 18 70 22
rect 62 11 70 18
rect 65 10 70 11
rect 72 10 77 30
rect 79 16 92 30
rect 94 16 99 30
rect 101 22 109 30
rect 101 18 103 22
rect 107 18 109 22
rect 101 16 109 18
rect 111 16 116 30
rect 118 21 128 30
rect 118 17 120 21
rect 124 17 128 21
rect 118 16 128 17
rect 79 12 90 16
rect 79 10 83 12
rect 81 8 83 10
rect 87 8 90 12
rect 81 7 90 8
rect 120 11 128 16
rect 130 29 138 30
rect 130 25 132 29
rect 136 25 138 29
rect 130 22 138 25
rect 130 18 132 22
rect 136 18 138 22
rect 130 11 138 18
rect 140 24 147 30
rect 140 20 142 24
rect 146 20 147 24
rect 140 16 147 20
rect 140 12 142 16
rect 146 12 147 16
rect 140 11 147 12
<< pdiffusion >>
rect 4 55 9 70
rect 2 54 9 55
rect 2 50 3 54
rect 7 50 9 54
rect 2 47 9 50
rect 2 43 3 47
rect 7 43 9 47
rect 2 42 9 43
rect 11 69 19 70
rect 11 65 13 69
rect 17 65 19 69
rect 11 62 19 65
rect 11 58 13 62
rect 17 58 19 62
rect 11 42 19 58
rect 21 54 29 70
rect 21 50 23 54
rect 27 50 29 54
rect 21 47 29 50
rect 21 43 23 47
rect 27 43 29 47
rect 21 42 29 43
rect 31 69 39 70
rect 31 65 33 69
rect 37 65 39 69
rect 31 62 39 65
rect 31 58 33 62
rect 37 58 39 62
rect 31 42 39 58
rect 41 67 46 70
rect 41 61 49 67
rect 41 57 43 61
rect 47 57 49 61
rect 41 54 49 57
rect 41 50 43 54
rect 47 50 49 54
rect 41 42 49 50
rect 51 63 59 67
rect 51 59 53 63
rect 57 59 59 63
rect 51 47 59 59
rect 51 43 53 47
rect 57 43 59 47
rect 51 42 59 43
rect 61 54 69 67
rect 61 50 63 54
rect 67 50 69 54
rect 61 47 69 50
rect 61 43 63 47
rect 67 43 69 47
rect 61 42 69 43
rect 71 63 79 67
rect 71 59 73 63
rect 77 59 79 63
rect 71 56 79 59
rect 71 52 73 56
rect 77 52 79 56
rect 71 42 79 52
rect 81 54 89 67
rect 81 50 83 54
rect 87 50 89 54
rect 81 47 89 50
rect 81 43 83 47
rect 87 43 89 47
rect 81 42 89 43
rect 91 61 96 67
rect 114 61 119 67
rect 91 56 99 61
rect 91 52 93 56
rect 97 52 99 56
rect 91 42 99 52
rect 101 47 109 61
rect 101 43 103 47
rect 107 43 109 47
rect 101 42 109 43
rect 111 55 119 61
rect 111 51 113 55
rect 117 51 119 55
rect 111 42 119 51
rect 121 54 129 67
rect 121 50 123 54
rect 127 50 129 54
rect 121 47 129 50
rect 121 43 123 47
rect 127 43 129 47
rect 121 42 129 43
rect 131 66 139 67
rect 131 62 133 66
rect 137 62 139 66
rect 131 58 139 62
rect 131 54 133 58
rect 137 54 139 58
rect 131 42 139 54
rect 141 54 149 67
rect 141 50 143 54
rect 147 50 149 54
rect 141 47 149 50
rect 141 43 143 47
rect 147 43 149 47
rect 141 42 149 43
rect 151 66 158 67
rect 151 62 153 66
rect 157 62 158 66
rect 151 58 158 62
rect 151 54 153 58
rect 157 54 158 58
rect 151 42 158 54
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect 118 78 122 82
rect 126 78 130 82
rect 134 78 138 82
rect 142 78 146 82
rect 150 78 154 82
rect 158 78 162 82
rect -2 69 162 78
rect -2 68 13 69
rect 12 65 13 68
rect 17 68 33 69
rect 17 65 18 68
rect 12 62 18 65
rect 12 58 13 62
rect 17 58 18 62
rect 32 65 33 68
rect 37 68 162 69
rect 37 65 38 68
rect 32 62 38 65
rect 133 66 137 68
rect 32 58 33 62
rect 37 58 38 62
rect 43 61 47 62
rect 52 59 53 63
rect 57 59 73 63
rect 77 59 97 63
rect 43 54 47 57
rect 73 56 77 59
rect 2 50 3 54
rect 7 50 23 54
rect 27 50 43 54
rect 47 50 63 54
rect 67 50 68 54
rect 93 56 97 59
rect 73 51 77 52
rect 82 54 87 55
rect 2 47 7 50
rect 2 43 3 47
rect 2 42 7 43
rect 23 47 28 50
rect 62 47 68 50
rect 82 50 83 54
rect 133 58 137 62
rect 97 52 113 55
rect 93 51 113 52
rect 117 51 118 55
rect 123 54 127 55
rect 82 47 87 50
rect 153 66 157 68
rect 153 58 157 62
rect 133 53 137 54
rect 143 54 147 55
rect 123 47 127 50
rect 27 43 28 47
rect 52 46 53 47
rect 23 42 28 43
rect 2 38 14 39
rect 2 34 10 38
rect 2 33 14 34
rect 2 25 6 33
rect 24 29 28 42
rect 42 43 53 46
rect 57 43 58 47
rect 62 43 63 47
rect 67 43 78 47
rect 82 43 83 47
rect 87 43 98 47
rect 102 43 103 47
rect 107 43 117 47
rect 42 42 58 43
rect 14 24 18 25
rect 14 16 18 20
rect 24 22 28 25
rect 24 17 28 18
rect 34 24 38 25
rect 34 16 38 20
rect 42 22 46 42
rect 67 38 71 39
rect 74 34 78 43
rect 94 38 98 43
rect 113 38 117 43
rect 153 53 157 54
rect 143 47 147 50
rect 127 43 143 46
rect 123 42 147 43
rect 82 34 85 38
rect 89 34 90 38
rect 94 34 100 38
rect 104 34 105 38
rect 113 34 116 38
rect 120 34 121 38
rect 67 30 71 34
rect 94 30 98 34
rect 132 30 136 42
rect 154 38 158 47
rect 145 34 146 38
rect 150 34 158 38
rect 145 33 158 34
rect 53 29 136 30
rect 53 25 54 29
rect 58 26 132 29
rect 58 25 59 26
rect 132 22 136 25
rect 42 18 44 22
rect 48 18 64 22
rect 68 18 103 22
rect 107 18 108 22
rect 120 21 124 22
rect 132 17 136 18
rect 142 24 146 25
rect 120 12 124 17
rect 142 16 146 20
rect -2 8 83 12
rect 87 8 162 12
rect -2 2 162 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 122 2
rect 126 -2 130 2
rect 134 -2 138 2
rect 142 -2 146 2
rect 150 -2 154 2
rect 158 -2 162 2
<< ntransistor >>
rect 20 11 22 30
rect 30 11 32 30
rect 50 11 52 30
rect 60 11 62 30
rect 70 10 72 30
rect 77 10 79 30
rect 92 16 94 30
rect 99 16 101 30
rect 109 16 111 30
rect 116 16 118 30
rect 128 11 130 30
rect 138 11 140 30
<< ptransistor >>
rect 9 42 11 70
rect 19 42 21 70
rect 29 42 31 70
rect 39 42 41 70
rect 49 42 51 67
rect 59 42 61 67
rect 69 42 71 67
rect 79 42 81 67
rect 89 42 91 67
rect 99 42 101 61
rect 109 42 111 61
rect 119 42 121 67
rect 129 42 131 67
rect 139 42 141 67
rect 149 42 151 67
<< polycontact >>
rect 10 34 14 38
rect 67 34 71 38
rect 78 34 82 38
rect 85 34 89 38
rect 100 34 104 38
rect 116 34 120 38
rect 146 34 150 38
<< ndcontact >>
rect 14 20 18 24
rect 14 12 18 16
rect 24 25 28 29
rect 24 18 28 22
rect 34 20 38 24
rect 44 18 48 22
rect 34 12 38 16
rect 54 25 58 29
rect 64 18 68 22
rect 103 18 107 22
rect 120 17 124 21
rect 83 8 87 12
rect 132 25 136 29
rect 132 18 136 22
rect 142 20 146 24
rect 142 12 146 16
<< pdcontact >>
rect 3 50 7 54
rect 3 43 7 47
rect 13 65 17 69
rect 13 58 17 62
rect 23 50 27 54
rect 23 43 27 47
rect 33 65 37 69
rect 33 58 37 62
rect 43 57 47 61
rect 43 50 47 54
rect 53 59 57 63
rect 53 43 57 47
rect 63 50 67 54
rect 63 43 67 47
rect 73 59 77 63
rect 73 52 77 56
rect 83 50 87 54
rect 83 43 87 47
rect 93 52 97 56
rect 103 43 107 47
rect 113 51 117 55
rect 123 50 127 54
rect 123 43 127 47
rect 133 62 137 66
rect 133 54 137 58
rect 143 50 147 54
rect 143 43 147 47
rect 153 62 157 66
rect 153 54 157 58
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
rect 90 -2 94 2
rect 98 -2 102 2
rect 106 -2 110 2
rect 114 -2 118 2
rect 122 -2 126 2
rect 130 -2 134 2
rect 138 -2 142 2
rect 146 -2 150 2
rect 154 -2 158 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
rect 90 78 94 82
rect 98 78 102 82
rect 106 78 110 82
rect 114 78 118 82
rect 122 78 126 82
rect 130 78 134 82
rect 138 78 142 82
rect 146 78 150 82
rect 154 78 158 82
<< psubstratepdiff >>
rect 0 2 160 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 122 2
rect 126 -2 130 2
rect 134 -2 138 2
rect 142 -2 146 2
rect 150 -2 154 2
rect 158 -2 160 2
rect 0 -3 160 -2
<< nsubstratendiff >>
rect 0 82 160 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect 118 78 122 82
rect 126 78 130 82
rect 134 78 138 82
rect 142 78 146 82
rect 150 78 154 82
rect 158 78 160 82
rect 0 77 160 78
<< labels >>
rlabel ptransistor 70 52 70 52 6 an
rlabel polysilicon 105 36 105 36 6 an
rlabel ntransistor 117 22 117 22 6 bn
rlabel metal1 4 32 4 32 6 b
rlabel polycontact 12 36 12 36 6 b
rlabel metal1 4 48 4 48 6 bn
rlabel metal1 26 35 26 35 6 bn
rlabel metal1 60 20 60 20 6 z
rlabel metal1 52 20 52 20 6 z
rlabel metal1 44 32 44 32 6 z
rlabel metal1 52 44 52 44 6 z
rlabel metal1 45 56 45 56 6 bn
rlabel metal1 80 6 80 6 6 vss
rlabel metal1 84 20 84 20 6 z
rlabel metal1 92 20 92 20 6 z
rlabel metal1 76 20 76 20 6 z
rlabel metal1 68 20 68 20 6 z
rlabel metal1 69 32 69 32 6 an
rlabel metal1 70 45 70 45 6 bn
rlabel metal1 82 36 82 36 6 bn
rlabel metal1 84 49 84 49 6 an
rlabel metal1 35 52 35 52 6 bn
rlabel metal1 80 74 80 74 6 vdd
rlabel metal1 100 20 100 20 6 z
rlabel metal1 90 45 90 45 6 an
rlabel metal1 99 36 99 36 6 an
rlabel metal1 115 40 115 40 6 bn
rlabel metal1 109 45 109 45 6 bn
rlabel metal1 125 48 125 48 6 an
rlabel metal1 94 28 94 28 6 an
rlabel metal1 134 31 134 31 6 an
rlabel metal1 156 40 156 40 6 a
rlabel polycontact 148 36 148 36 6 a
rlabel metal1 145 48 145 48 6 an
<< end >>
