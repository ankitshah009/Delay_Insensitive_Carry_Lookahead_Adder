magic
tech scmos
timestamp 1179387404
<< checkpaint >>
rect -22 -25 102 105
<< ab >>
rect 0 0 80 80
<< pwell >>
rect -4 -7 84 36
<< nwell >>
rect -4 36 84 87
<< polysilicon >>
rect 28 66 30 71
rect 38 70 40 74
rect 45 70 47 74
rect 55 70 57 74
rect 65 70 67 74
rect 9 58 11 63
rect 9 39 11 42
rect 28 39 30 50
rect 38 44 40 50
rect 9 38 30 39
rect 34 43 40 44
rect 34 39 35 43
rect 39 39 40 43
rect 34 38 40 39
rect 9 34 10 38
rect 14 37 30 38
rect 14 34 15 37
rect 9 33 15 34
rect 25 30 27 37
rect 35 30 37 38
rect 45 30 47 50
rect 55 47 57 50
rect 55 46 61 47
rect 55 42 56 46
rect 60 42 61 46
rect 55 41 61 42
rect 55 30 57 41
rect 65 39 67 50
rect 65 38 71 39
rect 65 35 66 38
rect 62 34 66 35
rect 70 34 71 38
rect 62 33 71 34
rect 62 30 64 33
rect 9 27 15 28
rect 9 23 10 27
rect 14 23 15 27
rect 9 22 15 23
rect 13 11 15 22
rect 25 15 27 20
rect 35 15 37 20
rect 45 11 47 20
rect 55 15 57 20
rect 62 15 64 20
rect 13 9 47 11
<< ndiffusion >>
rect 17 20 25 30
rect 27 27 35 30
rect 27 23 29 27
rect 33 23 35 27
rect 27 20 35 23
rect 37 29 45 30
rect 37 25 39 29
rect 43 25 45 29
rect 37 20 45 25
rect 47 29 55 30
rect 47 25 49 29
rect 53 25 55 29
rect 47 20 55 25
rect 57 20 62 30
rect 64 20 73 30
rect 17 16 18 20
rect 22 16 23 20
rect 17 15 23 16
rect 66 16 67 20
rect 71 16 73 20
rect 66 15 73 16
<< pdiffusion >>
rect 33 66 38 70
rect 23 63 28 66
rect 21 62 28 63
rect 21 58 22 62
rect 26 58 28 62
rect 2 57 9 58
rect 2 53 3 57
rect 7 53 9 57
rect 2 49 9 53
rect 2 45 3 49
rect 7 45 9 49
rect 2 42 9 45
rect 11 48 16 58
rect 21 57 28 58
rect 23 50 28 57
rect 30 55 38 66
rect 30 51 32 55
rect 36 51 38 55
rect 30 50 38 51
rect 40 50 45 70
rect 47 69 55 70
rect 47 65 49 69
rect 53 65 55 69
rect 47 50 55 65
rect 57 62 65 70
rect 57 58 59 62
rect 63 58 65 62
rect 57 50 65 58
rect 67 69 74 70
rect 67 65 69 69
rect 73 65 74 69
rect 67 62 74 65
rect 67 58 69 62
rect 73 58 74 62
rect 67 50 74 58
rect 11 47 18 48
rect 11 43 13 47
rect 17 43 18 47
rect 11 42 18 43
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect -2 69 82 78
rect -2 68 49 69
rect 3 57 7 68
rect 48 65 49 68
rect 53 68 69 69
rect 53 65 54 68
rect 68 65 69 68
rect 73 68 82 69
rect 73 65 74 68
rect 68 62 74 65
rect 21 58 22 62
rect 26 58 59 62
rect 63 58 64 62
rect 68 58 69 62
rect 73 58 74 62
rect 3 49 7 53
rect 26 51 32 55
rect 36 51 38 55
rect 26 49 38 51
rect 3 44 7 45
rect 12 43 13 47
rect 17 43 22 47
rect 2 38 14 39
rect 2 34 10 38
rect 2 33 14 34
rect 2 17 6 33
rect 18 27 22 43
rect 26 35 30 49
rect 42 43 46 58
rect 50 49 62 55
rect 56 46 62 49
rect 34 39 35 43
rect 39 39 51 43
rect 60 42 62 46
rect 56 41 62 42
rect 26 31 41 35
rect 37 29 41 31
rect 47 29 51 39
rect 66 38 70 39
rect 66 31 70 34
rect 9 23 10 27
rect 14 23 29 27
rect 33 23 34 27
rect 37 25 39 29
rect 43 25 44 29
rect 47 25 49 29
rect 53 25 54 29
rect 58 25 70 31
rect 67 20 71 21
rect 17 16 18 20
rect 22 16 23 20
rect 17 12 23 16
rect 67 12 71 16
rect -2 2 82 12
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
<< ntransistor >>
rect 25 20 27 30
rect 35 20 37 30
rect 45 20 47 30
rect 55 20 57 30
rect 62 20 64 30
<< ptransistor >>
rect 9 42 11 58
rect 28 50 30 66
rect 38 50 40 70
rect 45 50 47 70
rect 55 50 57 70
rect 65 50 67 70
<< polycontact >>
rect 35 39 39 43
rect 10 34 14 38
rect 56 42 60 46
rect 66 34 70 38
rect 10 23 14 27
<< ndcontact >>
rect 29 23 33 27
rect 39 25 43 29
rect 49 25 53 29
rect 18 16 22 20
rect 67 16 71 20
<< pdcontact >>
rect 22 58 26 62
rect 3 53 7 57
rect 3 45 7 49
rect 32 51 36 55
rect 49 65 53 69
rect 59 58 63 62
rect 69 65 73 69
rect 69 58 73 62
rect 13 43 17 47
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
<< psubstratepdiff >>
rect 0 2 80 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 80 2
rect 0 -3 80 -2
<< nsubstratendiff >>
rect 0 82 80 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 80 82
rect 0 77 80 78
<< labels >>
rlabel polycontact 12 25 12 25 6 bn
rlabel polycontact 37 41 37 41 6 an
rlabel metal1 4 28 4 28 6 b
rlabel polycontact 12 36 12 36 6 b
rlabel metal1 17 45 17 45 6 bn
rlabel metal1 28 44 28 44 6 z
rlabel metal1 40 6 40 6 6 vss
rlabel metal1 21 25 21 25 6 bn
rlabel metal1 36 52 36 52 6 z
rlabel metal1 40 74 40 74 6 vdd
rlabel metal1 60 28 60 28 6 a1
rlabel metal1 49 34 49 34 6 an
rlabel metal1 42 41 42 41 6 an
rlabel metal1 60 48 60 48 6 a2
rlabel metal1 52 52 52 52 6 a2
rlabel metal1 42 60 42 60 6 an
rlabel metal1 68 32 68 32 6 a1
<< end >>
