magic
tech scmos
timestamp 1179387314
<< checkpaint >>
rect -22 -22 86 94
<< ab >>
rect 0 0 64 72
<< pwell >>
rect -4 -4 68 32
<< nwell >>
rect -4 32 68 76
<< polysilicon >>
rect 28 58 30 63
rect 35 58 37 63
rect 42 58 44 63
rect 49 58 51 63
rect 9 51 11 56
rect 28 43 30 46
rect 19 42 30 43
rect 9 36 11 39
rect 19 38 20 42
rect 24 41 30 42
rect 24 38 25 41
rect 19 37 25 38
rect 9 35 15 36
rect 9 31 10 35
rect 14 31 15 35
rect 9 30 15 31
rect 9 26 11 30
rect 19 26 21 37
rect 35 35 37 46
rect 29 34 37 35
rect 29 30 30 34
rect 34 32 37 34
rect 34 30 35 32
rect 29 29 35 30
rect 29 26 31 29
rect 42 27 44 46
rect 49 43 51 46
rect 49 42 55 43
rect 49 38 50 42
rect 54 38 55 42
rect 49 37 55 38
rect 39 26 45 27
rect 9 15 11 20
rect 19 15 21 20
rect 29 15 31 20
rect 39 22 40 26
rect 44 22 45 26
rect 39 21 45 22
rect 39 18 41 21
rect 49 18 51 37
rect 39 7 41 12
rect 49 7 51 12
<< ndiffusion >>
rect 2 25 9 26
rect 2 21 3 25
rect 7 21 9 25
rect 2 20 9 21
rect 11 20 19 26
rect 21 25 29 26
rect 21 21 23 25
rect 27 21 29 25
rect 21 20 29 21
rect 31 20 37 26
rect 13 13 17 20
rect 33 18 37 20
rect 33 13 39 18
rect 13 12 19 13
rect 13 8 14 12
rect 18 8 19 12
rect 13 7 19 8
rect 31 12 39 13
rect 41 17 49 18
rect 41 13 43 17
rect 47 13 49 17
rect 41 12 49 13
rect 51 12 59 18
rect 31 8 37 12
rect 31 4 32 8
rect 36 4 37 8
rect 53 8 59 12
rect 31 3 37 4
rect 53 4 54 8
rect 58 4 59 8
rect 53 3 59 4
<< pdiffusion >>
rect 53 68 59 69
rect 53 64 54 68
rect 58 64 59 68
rect 13 61 19 62
rect 13 57 14 61
rect 18 57 19 61
rect 53 58 59 64
rect 13 56 19 57
rect 13 51 17 56
rect 23 52 28 58
rect 2 50 9 51
rect 2 46 3 50
rect 7 46 9 50
rect 2 45 9 46
rect 4 39 9 45
rect 11 39 17 51
rect 21 51 28 52
rect 21 47 22 51
rect 26 47 28 51
rect 21 46 28 47
rect 30 46 35 58
rect 37 46 42 58
rect 44 46 49 58
rect 51 46 59 58
<< metal1 >>
rect -2 68 66 72
rect -2 64 4 68
rect 8 64 54 68
rect 58 64 66 68
rect 14 61 18 64
rect 14 56 18 57
rect 2 50 7 51
rect 2 46 3 50
rect 2 45 7 46
rect 10 47 22 51
rect 26 47 27 51
rect 2 26 6 45
rect 10 35 14 47
rect 34 42 38 59
rect 42 53 54 59
rect 17 38 20 42
rect 24 38 38 42
rect 42 34 46 43
rect 50 42 54 53
rect 50 37 54 38
rect 14 31 25 34
rect 10 30 25 31
rect 29 30 30 34
rect 34 30 46 34
rect 2 25 16 26
rect 2 21 3 25
rect 7 21 16 25
rect 21 25 25 30
rect 21 21 23 25
rect 27 21 29 25
rect 39 22 40 26
rect 44 22 62 26
rect 25 17 29 21
rect 25 13 43 17
rect 47 13 48 17
rect 58 13 62 22
rect 14 12 18 13
rect -2 4 4 8
rect 8 4 32 8
rect 36 4 54 8
rect 58 4 66 8
rect -2 0 66 4
<< ntransistor >>
rect 9 20 11 26
rect 19 20 21 26
rect 29 20 31 26
rect 39 12 41 18
rect 49 12 51 18
<< ptransistor >>
rect 9 39 11 51
rect 28 46 30 58
rect 35 46 37 58
rect 42 46 44 58
rect 49 46 51 58
<< polycontact >>
rect 20 38 24 42
rect 10 31 14 35
rect 30 30 34 34
rect 50 38 54 42
rect 40 22 44 26
<< ndcontact >>
rect 3 21 7 25
rect 23 21 27 25
rect 14 8 18 12
rect 43 13 47 17
rect 32 4 36 8
rect 54 4 58 8
<< pdcontact >>
rect 54 64 58 68
rect 14 57 18 61
rect 3 46 7 50
rect 22 47 26 51
<< psubstratepcontact >>
rect 4 4 8 8
<< nsubstratencontact >>
rect 4 64 8 68
<< psubstratepdiff >>
rect 3 8 9 13
rect 3 4 4 8
rect 8 4 9 8
rect 3 3 9 4
<< nsubstratendiff >>
rect 3 68 9 69
rect 3 64 4 68
rect 8 64 9 68
rect 3 58 9 64
<< labels >>
rlabel polycontact 12 33 12 33 6 zn
rlabel metal1 12 24 12 24 6 z
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 40 12 40 6 zn
rlabel metal1 20 40 20 40 6 d
rlabel metal1 28 40 28 40 6 d
rlabel metal1 18 49 18 49 6 zn
rlabel metal1 32 4 32 4 6 vss
rlabel metal1 36 15 36 15 6 zn
rlabel metal1 36 32 36 32 6 c
rlabel metal1 44 24 44 24 6 b
rlabel metal1 44 40 44 40 6 c
rlabel metal1 36 52 36 52 6 d
rlabel metal1 44 56 44 56 6 a
rlabel metal1 32 68 32 68 6 vdd
rlabel metal1 60 16 60 16 6 b
rlabel metal1 52 24 52 24 6 b
rlabel metal1 52 48 52 48 6 a
<< end >>
