.subckt na2_x1 i0 i1 nq vdd vss
*   SPICE3 file   created from na2_x1.ext -      technology: scmos
m00 nq     i0     vdd    vdd p w=20u  l=2.3636u ad=100p     pd=30u      as=208p     ps=72u
m01 vdd    i1     nq     vdd p w=20u  l=2.3636u ad=208p     pd=72u      as=100p     ps=30u
m02 w1     i0     vss    vss n w=20u  l=2.3636u ad=60p      pd=26u      as=208p     ps=72u
m03 nq     i1     w1     vss n w=20u  l=2.3636u ad=160p     pd=56u      as=60p      ps=26u
C0  nq     vdd    0.046f
C1  i1     i0     0.184f
C2  i0     vdd    0.074f
C3  w1     nq     0.028f
C4  vss    i1     0.015f
C5  nq     i0     0.485f
C6  i1     vdd    0.074f
C7  vss    nq     0.111f
C8  vss    i0     0.074f
C9  nq     i1     0.456f
C11 nq     vss    0.021f
C12 i1     vss    0.044f
C13 i0     vss    0.040f
.ends
