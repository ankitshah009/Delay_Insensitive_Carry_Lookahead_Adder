magic
tech scmos
timestamp 1185094780
<< checkpaint >>
rect -22 -22 72 122
<< ab >>
rect 0 0 50 100
<< pwell >>
rect -4 -4 54 48
<< nwell >>
rect -4 48 54 104
<< polysilicon >>
rect 25 84 27 89
rect 33 84 35 89
rect 13 73 15 78
rect 13 53 15 61
rect 13 52 21 53
rect 13 48 16 52
rect 20 48 21 52
rect 13 47 21 48
rect 13 27 15 47
rect 25 43 27 61
rect 33 53 35 61
rect 33 52 43 53
rect 33 51 38 52
rect 37 48 38 51
rect 42 48 43 52
rect 37 47 43 48
rect 25 42 33 43
rect 25 38 28 42
rect 32 38 33 42
rect 25 37 33 38
rect 25 27 27 37
rect 37 27 39 47
rect 13 12 15 17
rect 25 12 27 17
rect 37 12 39 17
<< ndiffusion >>
rect 8 23 13 27
rect 5 22 13 23
rect 5 18 6 22
rect 10 18 13 22
rect 5 17 13 18
rect 15 22 25 27
rect 15 18 18 22
rect 22 18 25 22
rect 15 17 25 18
rect 27 17 37 27
rect 39 23 44 27
rect 39 22 47 23
rect 39 18 42 22
rect 46 18 47 22
rect 39 17 47 18
rect 29 12 35 17
rect 29 8 30 12
rect 34 8 35 12
rect 29 7 35 8
<< pdiffusion >>
rect 20 73 25 84
rect 5 72 13 73
rect 5 68 6 72
rect 10 68 13 72
rect 5 61 13 68
rect 15 72 25 73
rect 15 68 18 72
rect 22 68 25 72
rect 15 61 25 68
rect 27 61 33 84
rect 35 82 43 84
rect 35 78 38 82
rect 42 78 43 82
rect 35 61 43 78
<< metal1 >>
rect -2 96 52 100
rect -2 92 8 96
rect 12 92 18 96
rect 22 92 52 96
rect -2 88 52 92
rect 6 72 10 88
rect 38 82 42 88
rect 38 77 42 78
rect 6 67 10 68
rect 18 72 22 73
rect 27 68 42 73
rect 18 63 22 68
rect 8 57 22 63
rect 8 23 12 57
rect 16 52 22 53
rect 20 48 22 52
rect 16 47 22 48
rect 18 32 22 47
rect 28 42 32 63
rect 38 52 42 68
rect 38 47 42 48
rect 32 38 43 42
rect 28 37 43 38
rect 18 27 33 32
rect 5 22 12 23
rect 5 18 6 22
rect 10 18 12 22
rect 17 18 18 22
rect 22 18 42 22
rect 46 18 47 22
rect 5 17 12 18
rect -2 8 30 12
rect 34 8 52 12
rect -2 4 8 8
rect 12 4 18 8
rect 22 4 52 8
rect -2 0 52 4
<< ntransistor >>
rect 13 17 15 27
rect 25 17 27 27
rect 37 17 39 27
<< ptransistor >>
rect 13 61 15 73
rect 25 61 27 84
rect 33 61 35 84
<< polycontact >>
rect 16 48 20 52
rect 38 48 42 52
rect 28 38 32 42
<< ndcontact >>
rect 6 18 10 22
rect 18 18 22 22
rect 42 18 46 22
rect 30 8 34 12
<< pdcontact >>
rect 6 68 10 72
rect 18 68 22 72
rect 38 78 42 82
<< psubstratepcontact >>
rect 8 4 12 8
rect 18 4 22 8
<< nsubstratencontact >>
rect 8 92 12 96
rect 18 92 22 96
<< psubstratepdiff >>
rect 7 8 23 9
rect 7 4 8 8
rect 12 4 18 8
rect 22 4 23 8
rect 7 3 23 4
<< nsubstratendiff >>
rect 7 96 23 97
rect 7 92 8 96
rect 12 92 18 96
rect 22 92 23 96
rect 7 91 23 92
<< labels >>
rlabel metal1 10 40 10 40 6 z
rlabel metal1 20 40 20 40 6 b
rlabel metal1 20 65 20 65 6 z
rlabel metal1 25 6 25 6 6 vss
rlabel metal1 30 30 30 30 6 b
rlabel metal1 30 50 30 50 6 a2
rlabel metal1 30 70 30 70 6 a1
rlabel metal1 25 94 25 94 6 vdd
rlabel metal1 32 20 32 20 6 n2
rlabel metal1 40 40 40 40 6 a2
rlabel metal1 40 60 40 60 6 a1
<< end >>
