magic
tech scmos
timestamp 1179385630
<< checkpaint >>
rect -22 -25 110 105
<< ab >>
rect 0 0 88 80
<< pwell >>
rect -4 -7 92 36
<< nwell >>
rect -4 36 92 87
<< polysilicon >>
rect 9 62 11 67
rect 19 62 21 67
rect 39 63 41 68
rect 46 63 48 68
rect 56 63 58 68
rect 66 63 68 68
rect 76 67 78 72
rect 9 39 11 42
rect 19 39 21 46
rect 39 39 41 47
rect 46 39 48 47
rect 56 39 58 47
rect 66 39 68 47
rect 76 39 78 47
rect 5 38 11 39
rect 5 34 6 38
rect 10 34 11 38
rect 5 33 11 34
rect 17 38 23 39
rect 17 34 18 38
rect 22 34 23 38
rect 17 33 23 34
rect 32 38 42 39
rect 32 34 33 38
rect 37 34 42 38
rect 46 36 49 39
rect 32 33 42 34
rect 9 26 11 33
rect 19 23 21 33
rect 40 30 42 33
rect 47 30 49 36
rect 55 38 61 39
rect 55 34 56 38
rect 60 34 61 38
rect 55 33 61 34
rect 65 38 71 39
rect 65 34 66 38
rect 70 34 71 38
rect 65 33 71 34
rect 76 38 86 39
rect 76 34 81 38
rect 85 34 86 38
rect 76 33 86 34
rect 57 30 59 33
rect 67 30 69 33
rect 77 30 79 33
rect 9 11 11 16
rect 19 11 21 16
rect 40 18 42 23
rect 47 14 49 23
rect 57 18 59 23
rect 67 20 69 23
rect 63 18 69 20
rect 63 14 65 18
rect 47 12 65 14
rect 77 15 79 20
<< ndiffusion >>
rect 2 25 9 26
rect 2 21 3 25
rect 7 21 9 25
rect 2 20 9 21
rect 4 16 9 20
rect 11 23 16 26
rect 32 23 40 30
rect 42 23 47 30
rect 49 29 57 30
rect 49 25 51 29
rect 55 25 57 29
rect 49 23 57 25
rect 59 28 67 30
rect 59 24 61 28
rect 65 24 67 28
rect 59 23 67 24
rect 69 23 77 30
rect 11 21 19 23
rect 11 17 13 21
rect 17 17 19 21
rect 11 16 19 17
rect 21 21 28 23
rect 21 17 23 21
rect 27 17 28 21
rect 21 16 28 17
rect 32 12 38 23
rect 71 20 77 23
rect 79 29 86 30
rect 79 25 81 29
rect 85 25 86 29
rect 79 24 86 25
rect 79 20 84 24
rect 71 16 75 20
rect 69 15 75 16
rect 32 8 33 12
rect 37 8 38 12
rect 69 11 70 15
rect 74 11 75 15
rect 69 10 75 11
rect 32 7 38 8
<< pdiffusion >>
rect 70 63 76 67
rect 32 62 39 63
rect 2 61 9 62
rect 2 57 3 61
rect 7 57 9 61
rect 2 54 9 57
rect 2 50 3 54
rect 7 50 9 54
rect 2 49 9 50
rect 4 42 9 49
rect 11 61 19 62
rect 11 57 13 61
rect 17 57 19 61
rect 11 46 19 57
rect 21 61 28 62
rect 21 57 23 61
rect 27 57 28 61
rect 21 54 28 57
rect 21 50 23 54
rect 27 50 28 54
rect 21 49 28 50
rect 32 58 33 62
rect 37 58 39 62
rect 21 46 26 49
rect 32 47 39 58
rect 41 47 46 63
rect 48 53 56 63
rect 48 49 50 53
rect 54 49 56 53
rect 48 47 56 49
rect 58 62 66 63
rect 58 58 60 62
rect 64 58 66 62
rect 58 47 66 58
rect 68 62 76 63
rect 68 58 70 62
rect 74 58 76 62
rect 68 47 76 58
rect 78 63 83 67
rect 78 62 85 63
rect 78 58 80 62
rect 84 58 85 62
rect 78 55 85 58
rect 78 51 80 55
rect 84 51 85 55
rect 78 50 85 51
rect 78 47 83 50
rect 11 42 17 46
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect -2 68 90 78
rect 12 61 18 68
rect 32 62 38 68
rect 69 62 75 68
rect 2 57 3 61
rect 7 57 8 61
rect 12 57 13 61
rect 17 57 18 61
rect 22 57 23 61
rect 27 57 28 61
rect 32 58 33 62
rect 37 58 38 62
rect 42 58 60 62
rect 64 58 65 62
rect 69 58 70 62
rect 74 58 75 62
rect 80 62 84 63
rect 2 54 8 57
rect 22 54 28 57
rect 42 54 46 58
rect 80 55 84 58
rect 2 50 3 54
rect 7 50 17 54
rect 22 50 23 54
rect 27 50 46 54
rect 50 53 54 55
rect 13 47 17 50
rect 50 47 54 49
rect 2 39 6 47
rect 13 43 22 47
rect 2 38 14 39
rect 2 34 6 38
rect 10 34 14 38
rect 2 33 14 34
rect 18 38 22 43
rect 42 43 54 47
rect 22 34 33 38
rect 37 34 38 38
rect 18 29 22 34
rect 3 25 22 29
rect 42 29 46 43
rect 58 39 62 55
rect 50 38 62 39
rect 50 34 56 38
rect 60 34 62 38
rect 50 33 62 34
rect 66 51 80 54
rect 66 50 84 51
rect 66 38 70 50
rect 74 41 86 47
rect 81 38 86 41
rect 70 34 76 37
rect 66 33 76 34
rect 85 34 86 38
rect 81 33 86 34
rect 72 29 76 33
rect 42 25 51 29
rect 55 25 56 29
rect 61 28 65 29
rect 72 25 81 29
rect 85 25 86 29
rect 61 21 65 24
rect 3 20 7 21
rect 12 17 13 21
rect 17 17 18 21
rect 22 17 23 21
rect 27 17 65 21
rect 12 12 18 17
rect 70 15 74 16
rect -2 8 33 12
rect 37 11 70 12
rect 74 11 90 12
rect 37 8 90 11
rect -2 2 90 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
<< ntransistor >>
rect 9 16 11 26
rect 40 23 42 30
rect 47 23 49 30
rect 57 23 59 30
rect 67 23 69 30
rect 19 16 21 23
rect 77 20 79 30
<< ptransistor >>
rect 9 42 11 62
rect 19 46 21 62
rect 39 47 41 63
rect 46 47 48 63
rect 56 47 58 63
rect 66 47 68 63
rect 76 47 78 67
<< polycontact >>
rect 6 34 10 38
rect 18 34 22 38
rect 33 34 37 38
rect 56 34 60 38
rect 66 34 70 38
rect 81 34 85 38
<< ndcontact >>
rect 3 21 7 25
rect 51 25 55 29
rect 61 24 65 28
rect 13 17 17 21
rect 23 17 27 21
rect 81 25 85 29
rect 33 8 37 12
rect 70 11 74 15
<< pdcontact >>
rect 3 57 7 61
rect 3 50 7 54
rect 13 57 17 61
rect 23 57 27 61
rect 23 50 27 54
rect 33 58 37 62
rect 50 49 54 53
rect 60 58 64 62
rect 70 58 74 62
rect 80 58 84 62
rect 80 51 84 55
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
<< psubstratepdiff >>
rect 0 2 88 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 88 2
rect 0 -3 88 -2
<< nsubstratendiff >>
rect 0 82 88 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 88 82
rect 0 77 88 78
<< labels >>
rlabel polysilicon 20 39 20 39 6 an
rlabel polysilicon 37 36 37 36 6 an
rlabel polycontact 68 36 68 36 6 bn
rlabel ndcontact 5 24 5 24 6 an
rlabel metal1 4 40 4 40 6 a
rlabel metal1 12 36 12 36 6 a
rlabel metal1 5 55 5 55 6 an
rlabel metal1 25 55 25 55 6 n1
rlabel metal1 9 52 9 52 6 an
rlabel metal1 44 6 44 6 6 vss
rlabel metal1 28 36 28 36 6 an
rlabel metal1 44 36 44 36 6 z
rlabel metal1 34 52 34 52 6 n1
rlabel metal1 44 74 44 74 6 vdd
rlabel metal1 43 19 43 19 6 n3
rlabel metal1 63 23 63 23 6 n3
rlabel metal1 52 36 52 36 6 c
rlabel metal1 60 44 60 44 6 c
rlabel pdcontact 52 52 52 52 6 z
rlabel metal1 68 43 68 43 6 bn
rlabel metal1 53 60 53 60 6 n1
rlabel metal1 79 27 79 27 6 bn
rlabel metal1 84 40 84 40 6 b
rlabel metal1 76 44 76 44 6 b
rlabel metal1 82 56 82 56 6 bn
<< end >>
