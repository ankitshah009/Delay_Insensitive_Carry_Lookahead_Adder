magic
tech scmos
timestamp 1179385487
<< checkpaint >>
rect -22 -25 62 105
<< ab >>
rect 0 0 40 80
<< pwell >>
rect -4 -7 44 36
<< nwell >>
rect -4 36 44 87
<< polysilicon >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 69 31 74
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 9 38 22 39
rect 9 34 17 38
rect 21 34 22 38
rect 9 33 22 34
rect 26 38 32 39
rect 26 34 27 38
rect 31 34 32 38
rect 26 33 32 34
rect 9 30 11 33
rect 19 30 21 33
rect 29 30 31 33
rect 9 11 11 16
rect 19 11 21 16
rect 29 10 31 15
<< ndiffusion >>
rect 2 28 9 30
rect 2 24 3 28
rect 7 24 9 28
rect 2 21 9 24
rect 2 17 3 21
rect 7 17 9 21
rect 2 16 9 17
rect 11 22 19 30
rect 11 18 13 22
rect 17 18 19 22
rect 11 16 19 18
rect 21 21 29 30
rect 21 17 23 21
rect 27 17 29 21
rect 21 16 29 17
rect 23 15 29 16
rect 31 29 38 30
rect 31 25 33 29
rect 37 25 38 29
rect 31 22 38 25
rect 31 18 33 22
rect 37 18 38 22
rect 31 17 38 18
rect 31 15 36 17
<< pdiffusion >>
rect 2 69 9 70
rect 2 65 3 69
rect 7 65 9 69
rect 2 62 9 65
rect 2 58 3 62
rect 7 58 9 62
rect 2 42 9 58
rect 11 62 19 70
rect 11 58 13 62
rect 17 58 19 62
rect 11 55 19 58
rect 11 51 13 55
rect 17 51 19 55
rect 11 42 19 51
rect 21 69 27 70
rect 21 68 29 69
rect 21 64 23 68
rect 27 64 29 68
rect 21 61 29 64
rect 21 57 23 61
rect 27 57 29 61
rect 21 42 29 57
rect 31 62 36 69
rect 31 61 38 62
rect 31 57 33 61
rect 37 57 38 61
rect 31 54 38 57
rect 31 50 33 54
rect 37 50 38 54
rect 31 49 38 50
rect 31 42 36 49
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect -2 69 42 78
rect -2 68 3 69
rect 2 65 3 68
rect 7 68 42 69
rect 7 65 8 68
rect 2 62 8 65
rect 2 58 3 62
rect 7 58 8 62
rect 13 62 17 63
rect 13 55 17 58
rect 23 61 27 64
rect 23 56 27 57
rect 33 61 38 62
rect 37 57 38 61
rect 2 51 13 54
rect 2 50 17 51
rect 33 54 38 57
rect 37 50 38 54
rect 2 37 6 50
rect 33 49 38 50
rect 17 42 31 46
rect 17 38 21 39
rect 2 33 14 37
rect 3 28 7 29
rect 3 21 7 24
rect 10 23 14 33
rect 17 30 21 34
rect 26 38 31 42
rect 26 34 27 38
rect 26 33 31 34
rect 34 30 38 49
rect 17 29 38 30
rect 17 26 33 29
rect 37 26 38 29
rect 10 22 17 23
rect 33 22 37 25
rect 10 18 13 22
rect 10 17 17 18
rect 23 21 27 22
rect 33 17 37 18
rect 3 12 7 17
rect 23 12 27 17
rect -2 2 42 12
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
<< ntransistor >>
rect 9 16 11 30
rect 19 16 21 30
rect 29 15 31 30
<< ptransistor >>
rect 9 42 11 70
rect 19 42 21 70
rect 29 42 31 69
<< polycontact >>
rect 17 34 21 38
rect 27 34 31 38
<< ndcontact >>
rect 3 24 7 28
rect 3 17 7 21
rect 13 18 17 22
rect 23 17 27 21
rect 33 25 37 29
rect 33 18 37 22
<< pdcontact >>
rect 3 65 7 69
rect 3 58 7 62
rect 13 58 17 62
rect 13 51 17 55
rect 23 64 27 68
rect 23 57 27 61
rect 33 57 37 61
rect 33 50 37 54
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
<< psubstratepdiff >>
rect 0 2 40 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 40 2
rect 0 -3 40 -2
<< nsubstratendiff >>
rect 0 82 40 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 40 82
rect 0 77 40 78
<< labels >>
rlabel polysilicon 15 36 15 36 6 an
rlabel metal1 4 40 4 40 6 z
rlabel metal1 12 24 12 24 6 z
rlabel metal1 12 52 12 52 6 z
rlabel metal1 20 6 20 6 6 vss
rlabel metal1 19 32 19 32 6 an
rlabel metal1 28 40 28 40 6 a
rlabel metal1 20 44 20 44 6 a
rlabel metal1 20 74 20 74 6 vdd
rlabel metal1 35 23 35 23 6 an
rlabel metal1 36 44 36 44 6 an
<< end >>
