magic
tech scmos
timestamp 1180600761
<< checkpaint >>
rect -22 -22 102 122
<< ab >>
rect 0 0 80 100
<< pwell >>
rect -4 -4 84 48
<< nwell >>
rect -4 48 84 104
<< polysilicon >>
rect 11 94 13 98
rect 23 94 25 98
rect 35 94 37 98
rect 47 94 49 98
rect 11 41 13 55
rect 23 53 25 56
rect 35 53 37 56
rect 67 75 69 79
rect 23 52 43 53
rect 23 51 38 52
rect 37 48 38 51
rect 42 48 43 52
rect 37 47 43 48
rect 17 42 23 43
rect 17 41 18 42
rect 11 39 18 41
rect 11 25 13 39
rect 17 38 18 39
rect 22 41 23 42
rect 47 41 49 55
rect 67 43 69 55
rect 22 39 49 41
rect 22 38 23 39
rect 17 37 23 38
rect 37 32 43 33
rect 37 29 38 32
rect 23 28 38 29
rect 42 28 43 32
rect 23 27 43 28
rect 23 24 25 27
rect 35 24 37 27
rect 47 25 49 39
rect 57 42 69 43
rect 57 38 58 42
rect 62 38 69 42
rect 57 37 69 38
rect 67 25 69 37
rect 67 11 69 15
rect 11 2 13 6
rect 23 2 25 6
rect 35 2 37 6
rect 47 2 49 6
<< ndiffusion >>
rect 3 22 11 25
rect 3 18 4 22
rect 8 18 11 22
rect 3 12 11 18
rect 3 8 4 12
rect 8 8 11 12
rect 3 6 11 8
rect 13 24 18 25
rect 42 24 47 25
rect 13 6 23 24
rect 25 22 35 24
rect 25 18 28 22
rect 32 18 35 22
rect 25 6 35 18
rect 37 6 47 24
rect 49 15 67 25
rect 69 22 77 25
rect 69 18 72 22
rect 76 18 77 22
rect 69 15 77 18
rect 49 12 65 15
rect 49 8 52 12
rect 56 8 60 12
rect 64 8 65 12
rect 49 6 65 8
<< pdiffusion >>
rect 3 92 11 94
rect 3 88 4 92
rect 8 88 11 92
rect 3 82 11 88
rect 3 78 4 82
rect 8 78 11 82
rect 3 72 11 78
rect 3 68 4 72
rect 8 68 11 72
rect 3 62 11 68
rect 3 58 4 62
rect 8 58 11 62
rect 3 55 11 58
rect 13 56 23 94
rect 25 82 35 94
rect 25 78 28 82
rect 32 78 35 82
rect 25 72 35 78
rect 25 68 28 72
rect 32 68 35 72
rect 25 62 35 68
rect 25 58 28 62
rect 32 58 35 62
rect 25 56 35 58
rect 37 56 47 94
rect 13 55 18 56
rect 42 55 47 56
rect 49 92 65 94
rect 49 88 52 92
rect 56 88 60 92
rect 64 88 65 92
rect 49 75 65 88
rect 49 55 67 75
rect 69 72 77 75
rect 69 68 72 72
rect 76 68 77 72
rect 69 62 77 68
rect 69 58 72 62
rect 76 58 77 62
rect 69 55 77 58
<< metal1 >>
rect -2 96 82 100
rect -2 92 72 96
rect 76 92 82 96
rect -2 88 4 92
rect 8 88 52 92
rect 56 88 60 92
rect 64 88 82 92
rect 4 82 8 88
rect 4 72 8 78
rect 4 62 8 68
rect 4 57 8 58
rect 18 42 22 83
rect 4 22 8 23
rect 4 12 8 18
rect 18 17 22 38
rect 28 82 32 83
rect 28 72 32 78
rect 28 62 32 68
rect 28 22 32 58
rect 38 78 76 82
rect 38 52 42 78
rect 38 47 42 48
rect 58 42 62 73
rect 58 32 62 38
rect 37 28 38 32
rect 42 28 62 32
rect 28 17 32 18
rect 58 17 62 28
rect 72 72 76 78
rect 72 62 76 68
rect 72 22 76 58
rect 72 17 76 18
rect -2 8 4 12
rect 8 8 52 12
rect 56 8 60 12
rect 64 8 82 12
rect -2 0 82 8
<< ntransistor >>
rect 11 6 13 25
rect 23 6 25 24
rect 35 6 37 24
rect 47 6 49 25
rect 67 15 69 25
<< ptransistor >>
rect 11 55 13 94
rect 23 56 25 94
rect 35 56 37 94
rect 47 55 49 94
rect 67 55 69 75
<< polycontact >>
rect 38 48 42 52
rect 18 38 22 42
rect 38 28 42 32
rect 58 38 62 42
<< ndcontact >>
rect 4 18 8 22
rect 4 8 8 12
rect 28 18 32 22
rect 72 18 76 22
rect 52 8 56 12
rect 60 8 64 12
<< pdcontact >>
rect 4 88 8 92
rect 4 78 8 82
rect 4 68 8 72
rect 4 58 8 62
rect 28 78 32 82
rect 28 68 32 72
rect 28 58 32 62
rect 52 88 56 92
rect 60 88 64 92
rect 72 68 76 72
rect 72 58 76 62
<< nsubstratencontact >>
rect 72 92 76 96
<< nsubstratendiff >>
rect 71 96 77 97
rect 71 92 72 96
rect 76 92 77 96
rect 71 86 77 92
<< labels >>
rlabel metal1 30 50 30 50 6 nq
rlabel metal1 20 50 20 50 6 i
rlabel metal1 40 6 40 6 6 vss
rlabel polycontact 40 30 40 30 6 cmd
rlabel metal1 50 30 50 30 6 cmd
rlabel metal1 40 94 40 94 6 vdd
rlabel metal1 60 45 60 45 6 cmd
<< end >>
