magic
tech scmos
timestamp 1179387604
<< checkpaint >>
rect -22 -25 118 105
<< ab >>
rect 0 0 96 80
<< pwell >>
rect -4 -7 100 36
<< nwell >>
rect -4 36 100 87
<< polysilicon >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 69 31 74
rect 36 72 64 74
rect 36 69 38 72
rect 55 64 57 68
rect 62 64 64 72
rect 74 70 76 74
rect 9 39 11 42
rect 19 39 21 42
rect 9 38 15 39
rect 9 34 10 38
rect 14 34 15 38
rect 9 33 15 34
rect 19 38 25 39
rect 19 34 20 38
rect 24 34 25 38
rect 19 33 25 34
rect 29 34 31 42
rect 36 38 38 42
rect 55 39 57 42
rect 51 38 57 39
rect 51 34 52 38
rect 56 34 57 38
rect 10 24 12 33
rect 19 29 21 33
rect 29 32 57 34
rect 62 38 64 42
rect 74 39 76 42
rect 74 38 81 39
rect 62 37 70 38
rect 62 33 65 37
rect 69 33 70 37
rect 62 32 70 33
rect 74 34 76 38
rect 80 34 81 38
rect 74 33 81 34
rect 17 27 21 29
rect 37 28 39 32
rect 62 29 64 32
rect 74 29 76 33
rect 17 24 19 27
rect 27 24 29 28
rect 37 12 39 16
rect 62 12 64 16
rect 10 6 12 11
rect 17 6 19 11
rect 27 8 29 11
rect 74 8 76 16
rect 27 6 76 8
<< ndiffusion >>
rect 55 28 62 29
rect 32 24 37 28
rect 2 12 10 24
rect 2 8 3 12
rect 7 11 10 12
rect 12 11 17 24
rect 19 22 27 24
rect 19 18 21 22
rect 25 18 27 22
rect 19 11 27 18
rect 29 23 37 24
rect 29 19 31 23
rect 35 19 37 23
rect 29 16 37 19
rect 39 21 46 28
rect 39 17 41 21
rect 45 17 46 21
rect 39 16 46 17
rect 55 24 56 28
rect 60 24 62 28
rect 55 21 62 24
rect 55 17 56 21
rect 60 17 62 21
rect 55 16 62 17
rect 64 21 74 29
rect 64 17 68 21
rect 72 17 74 21
rect 64 16 74 17
rect 76 22 81 29
rect 76 21 83 22
rect 76 17 78 21
rect 82 17 83 21
rect 76 16 83 17
rect 29 11 34 16
rect 7 8 8 11
rect 2 7 8 8
<< pdiffusion >>
rect 4 64 9 70
rect 2 63 9 64
rect 2 59 3 63
rect 7 59 9 63
rect 2 58 9 59
rect 4 42 9 58
rect 11 54 19 70
rect 11 50 13 54
rect 17 50 19 54
rect 11 42 19 50
rect 21 69 26 70
rect 21 54 29 69
rect 21 50 23 54
rect 27 50 29 54
rect 21 47 29 50
rect 21 43 23 47
rect 27 43 29 47
rect 21 42 29 43
rect 31 42 36 69
rect 38 68 46 69
rect 38 64 40 68
rect 44 64 46 68
rect 66 69 74 70
rect 66 65 68 69
rect 72 65 74 69
rect 66 64 74 65
rect 38 54 46 64
rect 38 42 44 54
rect 50 48 55 64
rect 48 47 55 48
rect 48 43 49 47
rect 53 43 55 47
rect 48 42 55 43
rect 57 42 62 64
rect 64 42 74 64
rect 76 63 81 70
rect 76 62 83 63
rect 76 58 78 62
rect 82 58 83 62
rect 76 57 83 58
rect 76 42 81 57
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect -2 69 98 78
rect -2 68 68 69
rect 67 65 68 68
rect 72 68 98 69
rect 72 65 73 68
rect 40 63 44 64
rect 2 59 3 63
rect 7 59 36 63
rect 50 59 78 62
rect 32 58 78 59
rect 82 58 89 62
rect 32 55 54 58
rect 23 54 27 55
rect 2 50 13 54
rect 17 50 18 54
rect 2 22 6 50
rect 23 47 27 50
rect 10 43 23 46
rect 10 42 27 43
rect 10 38 14 42
rect 32 38 36 55
rect 19 34 20 38
rect 24 34 36 38
rect 42 43 49 47
rect 53 43 54 47
rect 10 30 14 34
rect 10 29 35 30
rect 42 29 46 43
rect 58 39 62 55
rect 66 49 78 55
rect 50 38 62 39
rect 66 38 70 39
rect 50 34 52 38
rect 56 34 62 38
rect 50 33 62 34
rect 65 37 70 38
rect 69 33 70 37
rect 74 38 78 49
rect 74 34 76 38
rect 80 34 81 38
rect 65 32 70 33
rect 66 30 70 32
rect 10 28 61 29
rect 10 26 56 28
rect 31 25 56 26
rect 31 23 35 25
rect 2 18 21 22
rect 25 18 26 22
rect 55 24 56 25
rect 60 24 61 28
rect 66 25 79 30
rect 55 21 61 24
rect 85 21 89 58
rect 31 18 35 19
rect 40 17 41 21
rect 45 17 46 21
rect 55 17 56 21
rect 60 17 61 21
rect 67 17 68 21
rect 72 17 73 21
rect 77 17 78 21
rect 82 17 89 21
rect 40 12 46 17
rect 67 12 73 17
rect -2 8 3 12
rect 7 8 98 12
rect -2 2 98 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
<< ntransistor >>
rect 10 11 12 24
rect 17 11 19 24
rect 27 11 29 24
rect 37 16 39 28
rect 62 16 64 29
rect 74 16 76 29
<< ptransistor >>
rect 9 42 11 70
rect 19 42 21 70
rect 29 42 31 69
rect 36 42 38 69
rect 55 42 57 64
rect 62 42 64 64
rect 74 42 76 70
<< polycontact >>
rect 10 34 14 38
rect 20 34 24 38
rect 52 34 56 38
rect 65 33 69 37
rect 76 34 80 38
<< ndcontact >>
rect 3 8 7 12
rect 21 18 25 22
rect 31 19 35 23
rect 41 17 45 21
rect 56 24 60 28
rect 56 17 60 21
rect 68 17 72 21
rect 78 17 82 21
<< pdcontact >>
rect 3 59 7 63
rect 13 50 17 54
rect 23 50 27 54
rect 23 43 27 47
rect 40 64 44 68
rect 68 65 72 69
rect 49 43 53 47
rect 78 58 82 62
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
rect 90 -2 94 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
rect 90 78 94 82
<< psubstratepdiff >>
rect 0 2 96 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 96 2
rect 0 -3 96 -2
<< nsubstratendiff >>
rect 0 82 96 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 96 82
rect 0 77 96 78
<< labels >>
rlabel polycontact 22 36 22 36 6 bn
rlabel polycontact 12 36 12 36 6 an
rlabel metal1 12 20 12 20 6 z
rlabel polycontact 12 36 12 36 6 an
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 52 12 52 6 z
rlabel metal1 20 20 20 20 6 z
rlabel metal1 33 24 33 24 6 an
rlabel metal1 27 36 27 36 6 bn
rlabel metal1 25 48 25 48 6 an
rlabel metal1 19 61 19 61 6 bn
rlabel metal1 48 6 48 6 6 vss
rlabel metal1 48 45 48 45 6 an
rlabel metal1 52 36 52 36 6 a2
rlabel metal1 48 74 48 74 6 vdd
rlabel metal1 58 23 58 23 6 an
rlabel metal1 76 28 76 28 6 a1
rlabel metal1 68 32 68 32 6 a1
rlabel metal1 60 44 60 44 6 a2
rlabel metal1 68 52 68 52 6 b
rlabel metal1 76 48 76 48 6 b
rlabel metal1 83 19 83 19 6 bn
rlabel metal1 69 60 69 60 6 bn
<< end >>
