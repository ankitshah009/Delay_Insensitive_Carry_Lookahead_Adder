magic
tech scmos
timestamp 1179386329
<< checkpaint >>
rect -22 -25 94 105
<< ab >>
rect 0 0 72 80
<< pwell >>
rect -4 -7 76 36
<< nwell >>
rect -4 36 76 87
<< polysilicon >>
rect 9 66 11 71
rect 19 69 21 74
rect 29 69 31 74
rect 39 66 41 71
rect 49 66 51 71
rect 59 60 61 65
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 39 39 41 42
rect 49 39 51 42
rect 59 39 61 42
rect 9 38 15 39
rect 9 34 10 38
rect 14 34 15 38
rect 9 33 15 34
rect 19 38 33 39
rect 19 34 26 38
rect 30 34 33 38
rect 19 33 33 34
rect 12 30 14 33
rect 19 30 21 33
rect 31 30 33 33
rect 38 38 51 39
rect 38 34 42 38
rect 46 34 51 38
rect 38 33 51 34
rect 55 38 63 39
rect 55 34 58 38
rect 62 34 63 38
rect 55 33 63 34
rect 38 30 40 33
rect 48 30 50 33
rect 55 30 57 33
rect 12 6 14 10
rect 19 6 21 10
rect 31 6 33 10
rect 38 6 40 10
rect 48 6 50 10
rect 55 6 57 10
<< ndiffusion >>
rect 5 29 12 30
rect 5 25 6 29
rect 10 25 12 29
rect 5 22 12 25
rect 5 18 6 22
rect 10 18 12 22
rect 5 17 12 18
rect 7 10 12 17
rect 14 10 19 30
rect 21 15 31 30
rect 21 11 24 15
rect 28 11 31 15
rect 21 10 31 11
rect 33 10 38 30
rect 40 22 48 30
rect 40 18 42 22
rect 46 18 48 22
rect 40 10 48 18
rect 50 10 55 30
rect 57 15 65 30
rect 57 11 59 15
rect 63 11 65 15
rect 57 10 65 11
<< pdiffusion >>
rect 14 66 19 69
rect 2 65 9 66
rect 2 61 3 65
rect 7 61 9 65
rect 2 57 9 61
rect 2 53 3 57
rect 7 53 9 57
rect 2 42 9 53
rect 11 54 19 66
rect 11 50 13 54
rect 17 50 19 54
rect 11 47 19 50
rect 11 43 13 47
rect 17 43 19 47
rect 11 42 19 43
rect 21 68 29 69
rect 21 64 23 68
rect 27 64 29 68
rect 21 61 29 64
rect 21 57 23 61
rect 27 57 29 61
rect 21 42 29 57
rect 31 66 36 69
rect 31 62 39 66
rect 31 58 33 62
rect 37 58 39 62
rect 31 54 39 58
rect 31 50 33 54
rect 37 50 39 54
rect 31 42 39 50
rect 41 65 49 66
rect 41 61 43 65
rect 47 61 49 65
rect 41 42 49 61
rect 51 60 56 66
rect 51 54 59 60
rect 51 50 53 54
rect 57 50 59 54
rect 51 42 59 50
rect 61 59 68 60
rect 61 55 63 59
rect 67 55 68 59
rect 61 42 68 55
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect -2 68 74 78
rect 3 65 7 68
rect 3 57 7 61
rect 22 64 23 68
rect 27 64 28 68
rect 22 61 28 64
rect 43 65 47 68
rect 22 57 23 61
rect 27 57 28 61
rect 33 62 38 63
rect 37 58 38 62
rect 43 60 47 61
rect 33 54 38 58
rect 63 59 67 68
rect 63 54 67 55
rect 3 52 7 53
rect 12 50 13 54
rect 17 50 33 54
rect 37 50 53 54
rect 57 50 58 54
rect 12 47 18 50
rect 2 43 13 47
rect 17 43 18 47
rect 2 25 6 43
rect 25 42 63 46
rect 10 38 21 39
rect 14 34 21 38
rect 25 38 31 42
rect 57 38 63 42
rect 25 34 26 38
rect 30 34 31 38
rect 41 34 42 38
rect 46 34 47 38
rect 57 34 58 38
rect 62 34 63 38
rect 10 33 21 34
rect 17 30 21 33
rect 41 30 47 34
rect 10 25 11 29
rect 17 26 47 30
rect 5 22 11 25
rect 5 18 6 22
rect 10 18 42 22
rect 46 18 47 22
rect 23 12 24 15
rect -2 11 24 12
rect 28 12 29 15
rect 58 12 59 15
rect 28 11 59 12
rect 63 12 64 15
rect 63 11 74 12
rect -2 2 74 11
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
<< ntransistor >>
rect 12 10 14 30
rect 19 10 21 30
rect 31 10 33 30
rect 38 10 40 30
rect 48 10 50 30
rect 55 10 57 30
<< ptransistor >>
rect 9 42 11 66
rect 19 42 21 69
rect 29 42 31 69
rect 39 42 41 66
rect 49 42 51 66
rect 59 42 61 60
<< polycontact >>
rect 10 34 14 38
rect 26 34 30 38
rect 42 34 46 38
rect 58 34 62 38
<< ndcontact >>
rect 6 25 10 29
rect 6 18 10 22
rect 24 11 28 15
rect 42 18 46 22
rect 59 11 63 15
<< pdcontact >>
rect 3 61 7 65
rect 3 53 7 57
rect 13 50 17 54
rect 13 43 17 47
rect 23 64 27 68
rect 23 57 27 61
rect 33 58 37 62
rect 33 50 37 54
rect 43 61 47 65
rect 53 50 57 54
rect 63 55 67 59
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
<< psubstratepdiff >>
rect 0 2 72 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 72 2
rect 0 -3 72 -2
<< nsubstratendiff >>
rect 0 82 72 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 72 82
rect 0 77 72 78
<< labels >>
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 20 12 20 6 z
rlabel metal1 20 28 20 28 6 b
rlabel metal1 20 20 20 20 6 z
rlabel polycontact 12 36 12 36 6 b
rlabel metal1 20 52 20 52 6 z
rlabel metal1 36 6 36 6 6 vss
rlabel metal1 28 28 28 28 6 b
rlabel metal1 28 20 28 20 6 z
rlabel metal1 36 28 36 28 6 b
rlabel metal1 36 20 36 20 6 z
rlabel metal1 28 40 28 40 6 a
rlabel metal1 36 44 36 44 6 a
rlabel metal1 28 52 28 52 6 z
rlabel metal1 36 56 36 56 6 z
rlabel metal1 36 74 36 74 6 vdd
rlabel ndcontact 44 20 44 20 6 z
rlabel metal1 44 32 44 32 6 b
rlabel metal1 44 44 44 44 6 a
rlabel metal1 52 44 52 44 6 a
rlabel metal1 52 52 52 52 6 z
rlabel metal1 44 52 44 52 6 z
rlabel metal1 60 40 60 40 6 a
<< end >>
