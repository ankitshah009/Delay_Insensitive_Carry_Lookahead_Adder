.subckt oai22v0x2 a1 a2 b1 b2 vdd vss z
*   SPICE3 file   created from oai22v0x2.ext -      technology: scmos
m00 w1     b1     vdd    vdd p w=28u  l=2.3636u ad=70p      pd=33u      as=215.25p  ps=58u
m01 z      b2     w1     vdd p w=28u  l=2.3636u ad=112p     pd=36u      as=70p      ps=33u
m02 w2     b2     z      vdd p w=28u  l=2.3636u ad=70p      pd=33u      as=112p     ps=36u
m03 vdd    b1     w2     vdd p w=28u  l=2.3636u ad=215.25p  pd=58u      as=70p      ps=33u
m04 w3     a1     vdd    vdd p w=28u  l=2.3636u ad=70p      pd=33u      as=215.25p  ps=58u
m05 z      a2     w3     vdd p w=28u  l=2.3636u ad=112p     pd=36u      as=70p      ps=33u
m06 w4     a2     z      vdd p w=28u  l=2.3636u ad=70p      pd=33u      as=112p     ps=36u
m07 vdd    a1     w4     vdd p w=28u  l=2.3636u ad=215.25p  pd=58u      as=70p      ps=33u
m08 z      b1     n3     vss n w=14u  l=2.3636u ad=56p      pd=22u      as=63.1373p ps=28.2745u
m09 n3     b2     z      vss n w=14u  l=2.3636u ad=63.1373p pd=28.2745u as=56p      ps=22u
m10 z      b2     n3     vss n w=14u  l=2.3636u ad=56p      pd=22u      as=63.1373p ps=28.2745u
m11 n3     b1     z      vss n w=14u  l=2.3636u ad=63.1373p pd=28.2745u as=56p      ps=22u
m12 vss    a1     n3     vss n w=14u  l=2.3636u ad=87.0435p pd=33.4783u as=63.1373p ps=28.2745u
m13 n3     a2     vss    vss n w=14u  l=2.3636u ad=63.1373p pd=28.2745u as=87.0435p ps=33.4783u
m14 vss    a2     n3     vss n w=9u   l=2.3636u ad=55.9565p pd=21.5217u as=40.5882p ps=18.1765u
m15 n3     a1     vss    vss n w=9u   l=2.3636u ad=40.5882p pd=18.1765u as=55.9565p ps=21.5217u
C0  w2     z      0.010f
C1  vss    vdd    0.003f
C2  a1     b1     0.135f
C3  z      w1     0.010f
C4  w2     vdd    0.005f
C5  n3     a2     0.102f
C6  vss    a1     0.046f
C7  w4     vdd    0.005f
C8  z      a2     0.028f
C9  w1     vdd    0.005f
C10 vss    b1     0.047f
C11 n3     b2     0.043f
C12 w4     a1     0.016f
C13 w2     b1     0.007f
C14 vdd    a2     0.021f
C15 z      b2     0.152f
C16 vdd    b2     0.022f
C17 a2     a1     0.298f
C18 w1     b1     0.007f
C19 w3     z      0.010f
C20 n3     z      0.430f
C21 a1     b2     0.033f
C22 a2     b1     0.031f
C23 w3     vdd    0.005f
C24 vss    a2     0.036f
C25 n3     vdd    0.032f
C26 b2     b1     0.341f
C27 w3     a1     0.007f
C28 z      vdd    0.409f
C29 n3     a1     0.107f
C30 vss    b2     0.024f
C31 z      a1     0.176f
C32 n3     b1     0.093f
C33 vss    n3     0.574f
C34 z      b1     0.476f
C35 vdd    a1     0.147f
C36 vss    z      0.134f
C37 a2     b2     0.027f
C38 vdd    b1     0.068f
C40 n3     vss    0.006f
C41 z      vss    0.010f
C43 a2     vss    0.033f
C44 a1     vss    0.032f
C45 b2     vss    0.029f
C46 b1     vss    0.033f
.ends
