magic
tech scmos
timestamp 1185039097
<< checkpaint >>
rect -22 -24 92 124
<< ab >>
rect 0 0 70 100
<< pwell >>
rect -2 -4 72 49
<< nwell >>
rect -2 49 72 104
<< polysilicon >>
rect 45 95 47 98
rect 57 95 59 98
rect 11 85 13 88
rect 19 85 21 88
rect 27 85 29 88
rect 11 33 13 55
rect 19 43 21 55
rect 27 53 29 55
rect 27 52 33 53
rect 27 48 28 52
rect 32 48 33 52
rect 27 47 33 48
rect 17 42 23 43
rect 17 38 18 42
rect 22 38 23 42
rect 17 37 23 38
rect 7 32 13 33
rect 7 28 8 32
rect 12 28 13 32
rect 7 27 13 28
rect 19 29 21 37
rect 31 29 33 47
rect 45 43 47 55
rect 57 43 59 55
rect 37 42 59 43
rect 37 38 38 42
rect 42 38 59 42
rect 37 37 59 38
rect 19 27 25 29
rect 31 27 37 29
rect 11 25 13 27
rect 23 25 25 27
rect 35 25 37 27
rect 45 25 47 37
rect 57 25 59 37
rect 11 12 13 15
rect 23 12 25 15
rect 35 12 37 15
rect 45 2 47 5
rect 57 2 59 5
<< ndiffusion >>
rect 3 22 11 25
rect 3 18 4 22
rect 8 18 11 22
rect 3 15 11 18
rect 13 15 23 25
rect 25 22 35 25
rect 25 18 28 22
rect 32 18 35 22
rect 25 15 35 18
rect 37 15 45 25
rect 15 12 21 15
rect 15 8 16 12
rect 20 8 21 12
rect 39 9 45 15
rect 15 7 21 8
rect 37 8 45 9
rect 37 4 38 8
rect 42 5 45 8
rect 47 22 57 25
rect 47 18 50 22
rect 54 18 57 22
rect 47 5 57 18
rect 59 22 67 25
rect 59 18 62 22
rect 66 18 67 22
rect 59 12 67 18
rect 59 8 62 12
rect 66 8 67 12
rect 59 5 67 8
rect 42 4 43 5
rect 37 3 43 4
<< pdiffusion >>
rect 31 92 45 95
rect 31 88 38 92
rect 42 88 45 92
rect 31 85 45 88
rect 3 82 11 85
rect 3 78 4 82
rect 8 78 11 82
rect 3 55 11 78
rect 13 55 19 85
rect 21 55 27 85
rect 29 55 45 85
rect 47 82 57 95
rect 47 78 50 82
rect 54 78 57 82
rect 47 72 57 78
rect 47 68 50 72
rect 54 68 57 72
rect 47 62 57 68
rect 47 58 50 62
rect 54 58 57 62
rect 47 55 57 58
rect 59 92 67 95
rect 59 88 62 92
rect 66 88 67 92
rect 59 82 67 88
rect 59 78 62 82
rect 66 78 67 82
rect 59 72 67 78
rect 59 68 62 72
rect 66 68 67 72
rect 59 62 67 68
rect 59 58 62 62
rect 66 58 67 62
rect 59 55 67 58
<< metal1 >>
rect -2 96 72 101
rect -2 92 4 96
rect 8 92 20 96
rect 24 92 72 96
rect -2 88 38 92
rect 42 88 62 92
rect 66 88 72 92
rect -2 87 72 88
rect 3 82 9 83
rect 49 82 55 83
rect 3 78 4 82
rect 8 78 42 82
rect 3 77 9 78
rect 7 32 13 72
rect 7 28 8 32
rect 12 28 13 32
rect 17 42 23 72
rect 17 38 18 42
rect 22 38 23 42
rect 17 28 23 38
rect 27 52 33 72
rect 27 48 28 52
rect 32 48 33 52
rect 27 28 33 48
rect 38 43 42 78
rect 47 78 50 82
rect 54 78 55 82
rect 47 77 55 78
rect 61 82 67 87
rect 61 78 62 82
rect 66 78 67 82
rect 47 73 53 77
rect 47 72 55 73
rect 47 68 50 72
rect 54 68 55 72
rect 47 67 55 68
rect 61 72 67 78
rect 61 68 62 72
rect 66 68 67 72
rect 47 63 53 67
rect 47 62 55 63
rect 47 58 50 62
rect 54 58 55 62
rect 47 57 55 58
rect 61 62 67 68
rect 61 58 62 62
rect 66 58 67 62
rect 61 57 67 58
rect 37 42 43 43
rect 37 38 38 42
rect 42 38 43 42
rect 37 37 43 38
rect 7 27 13 28
rect 3 22 9 23
rect 27 22 33 23
rect 38 22 42 37
rect 3 18 4 22
rect 8 18 28 22
rect 32 18 42 22
rect 47 23 53 57
rect 47 22 55 23
rect 47 18 50 22
rect 54 18 55 22
rect 3 17 9 18
rect 27 17 33 18
rect 49 17 55 18
rect 61 22 67 23
rect 61 18 62 22
rect 66 18 67 22
rect 61 13 67 18
rect -2 12 72 13
rect -2 8 16 12
rect 20 8 62 12
rect 66 8 72 12
rect -2 4 38 8
rect 42 4 72 8
rect -2 -1 72 4
<< ntransistor >>
rect 11 15 13 25
rect 23 15 25 25
rect 35 15 37 25
rect 45 5 47 25
rect 57 5 59 25
<< ptransistor >>
rect 11 55 13 85
rect 19 55 21 85
rect 27 55 29 85
rect 45 55 47 95
rect 57 55 59 95
<< polycontact >>
rect 28 48 32 52
rect 18 38 22 42
rect 8 28 12 32
rect 38 38 42 42
<< ndcontact >>
rect 4 18 8 22
rect 28 18 32 22
rect 16 8 20 12
rect 38 4 42 8
rect 50 18 54 22
rect 62 18 66 22
rect 62 8 66 12
<< pdcontact >>
rect 38 88 42 92
rect 4 78 8 82
rect 50 78 54 82
rect 50 68 54 72
rect 50 58 54 62
rect 62 88 66 92
rect 62 78 66 82
rect 62 68 66 72
rect 62 58 66 62
<< nsubstratencontact >>
rect 4 92 8 96
rect 20 92 24 96
<< nsubstratendiff >>
rect 3 96 25 97
rect 3 92 4 96
rect 8 92 20 96
rect 24 92 25 96
rect 3 91 25 92
<< labels >>
rlabel metal1 10 50 10 50 6 i2
rlabel metal1 10 50 10 50 6 i2
rlabel polycontact 30 50 30 50 6 i0
rlabel metal1 20 50 20 50 6 i1
rlabel metal1 20 50 20 50 6 i1
rlabel polycontact 30 50 30 50 6 i0
rlabel metal1 35 6 35 6 6 vss
rlabel metal1 35 6 35 6 6 vss
rlabel metal1 50 50 50 50 6 q
rlabel metal1 50 50 50 50 6 q
rlabel metal1 35 94 35 94 6 vdd
rlabel metal1 35 94 35 94 6 vdd
<< end >>
