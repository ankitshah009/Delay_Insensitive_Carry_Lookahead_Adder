magic
tech scmos
timestamp 1179386284
<< checkpaint >>
rect -22 -22 54 94
<< ab >>
rect 0 0 32 72
<< pwell >>
rect -4 -4 36 32
<< nwell >>
rect -4 32 36 76
<< polysilicon >>
rect 10 58 16 59
rect 10 54 11 58
rect 15 54 16 58
rect 10 53 16 54
rect 10 46 12 53
rect 20 46 22 51
rect 10 35 12 38
rect 20 35 22 38
rect 9 32 12 35
rect 16 34 23 35
rect 9 26 11 32
rect 16 30 18 34
rect 22 30 23 34
rect 16 29 23 30
rect 16 26 18 29
rect 9 14 11 19
rect 16 14 18 19
<< ndiffusion >>
rect 2 25 9 26
rect 2 21 3 25
rect 7 21 9 25
rect 2 19 9 21
rect 11 19 16 26
rect 18 19 27 26
rect 20 17 27 19
rect 20 13 21 17
rect 25 13 27 17
rect 20 12 27 13
<< pdiffusion >>
rect 2 68 8 69
rect 2 64 3 68
rect 7 64 8 68
rect 2 46 8 64
rect 2 38 10 46
rect 12 43 20 46
rect 12 39 14 43
rect 18 39 20 43
rect 12 38 20 39
rect 22 45 30 46
rect 22 41 25 45
rect 29 41 30 45
rect 22 38 30 41
<< metal1 >>
rect -2 68 34 72
rect -2 64 3 68
rect 7 64 16 68
rect 20 64 24 68
rect 28 64 34 68
rect 2 58 16 59
rect 2 54 11 58
rect 15 54 16 58
rect 2 45 6 54
rect 25 45 29 64
rect 10 40 14 43
rect 2 36 14 40
rect 18 39 19 43
rect 25 40 29 41
rect 2 26 6 36
rect 18 34 30 35
rect 22 30 30 34
rect 18 29 30 30
rect 2 25 7 26
rect 2 21 3 25
rect 26 21 30 29
rect 2 20 7 21
rect 20 13 21 17
rect 25 13 26 17
rect 20 8 26 13
rect -2 4 4 8
rect 8 4 11 8
rect 15 4 34 8
rect -2 0 34 4
<< ntransistor >>
rect 9 19 11 26
rect 16 19 18 26
<< ptransistor >>
rect 10 38 12 46
rect 20 38 22 46
<< polycontact >>
rect 11 54 15 58
rect 18 30 22 34
<< ndcontact >>
rect 3 21 7 25
rect 21 13 25 17
<< pdcontact >>
rect 3 64 7 68
rect 14 39 18 43
rect 25 41 29 45
<< psubstratepcontact >>
rect 4 4 8 8
rect 11 4 15 8
<< nsubstratencontact >>
rect 16 64 20 68
rect 24 64 28 68
<< psubstratepdiff >>
rect 3 8 16 9
rect 3 4 4 8
rect 8 4 11 8
rect 15 4 16 8
rect 3 3 16 4
<< nsubstratendiff >>
rect 15 68 29 69
rect 15 64 16 68
rect 20 64 24 68
rect 28 64 29 68
rect 15 63 29 64
<< labels >>
rlabel metal1 4 28 4 28 6 z
rlabel metal1 4 52 4 52 6 b
rlabel metal1 12 40 12 40 6 z
rlabel polycontact 12 56 12 56 6 b
rlabel metal1 16 4 16 4 6 vss
rlabel polycontact 20 32 20 32 6 a
rlabel metal1 16 68 16 68 6 vdd
rlabel metal1 28 28 28 28 6 a
<< end >>
