magic
tech scmos
timestamp 1179386276
<< checkpaint >>
rect -22 -22 134 94
<< ab >>
rect 0 0 112 72
<< pwell >>
rect -4 -4 116 32
<< nwell >>
rect -4 32 116 76
<< polysilicon >>
rect 9 64 11 69
rect 19 64 21 69
rect 29 64 31 69
rect 39 64 41 69
rect 49 64 51 69
rect 59 64 61 69
rect 69 56 71 61
rect 79 56 81 61
rect 91 60 93 65
rect 101 60 103 65
rect 9 35 11 38
rect 19 35 21 38
rect 29 35 31 38
rect 39 35 41 38
rect 9 34 15 35
rect 9 30 10 34
rect 14 30 15 34
rect 9 29 15 30
rect 19 34 31 35
rect 19 30 26 34
rect 30 30 31 34
rect 19 29 31 30
rect 35 34 41 35
rect 35 30 36 34
rect 40 31 41 34
rect 49 31 51 38
rect 59 35 61 38
rect 69 35 71 38
rect 59 34 71 35
rect 40 30 54 31
rect 35 29 54 30
rect 12 26 14 29
rect 19 26 21 29
rect 29 26 31 29
rect 36 26 38 29
rect 52 26 54 29
rect 59 30 60 34
rect 64 30 71 34
rect 79 35 81 38
rect 91 35 93 38
rect 101 35 103 38
rect 79 34 87 35
rect 79 31 82 34
rect 59 29 71 30
rect 59 26 61 29
rect 69 26 71 29
rect 76 30 82 31
rect 86 30 87 34
rect 76 29 87 30
rect 91 34 103 35
rect 91 30 98 34
rect 102 30 103 34
rect 91 29 103 30
rect 76 26 78 29
rect 91 26 93 29
rect 101 26 103 29
rect 91 10 93 15
rect 101 11 103 15
rect 12 2 14 6
rect 19 2 21 6
rect 29 2 31 6
rect 36 2 38 6
rect 52 2 54 6
rect 59 2 61 6
rect 69 2 71 6
rect 76 2 78 6
<< ndiffusion >>
rect 4 11 12 26
rect 4 7 6 11
rect 10 7 12 11
rect 4 6 12 7
rect 14 6 19 26
rect 21 18 29 26
rect 21 14 23 18
rect 27 14 29 18
rect 21 6 29 14
rect 31 6 36 26
rect 38 11 52 26
rect 38 7 43 11
rect 47 7 52 11
rect 38 6 52 7
rect 54 6 59 26
rect 61 18 69 26
rect 61 14 63 18
rect 67 14 69 18
rect 61 6 69 14
rect 71 6 76 26
rect 78 18 91 26
rect 78 14 82 18
rect 86 15 91 18
rect 93 25 101 26
rect 93 21 95 25
rect 99 21 101 25
rect 93 15 101 21
rect 103 20 110 26
rect 103 16 105 20
rect 109 16 110 20
rect 103 15 110 16
rect 86 14 89 15
rect 78 11 89 14
rect 78 7 82 11
rect 86 7 89 11
rect 78 6 89 7
<< pdiffusion >>
rect 2 63 9 64
rect 2 59 3 63
rect 7 59 9 63
rect 2 38 9 59
rect 11 57 19 64
rect 11 53 13 57
rect 17 53 19 57
rect 11 50 19 53
rect 11 46 13 50
rect 17 46 19 50
rect 11 38 19 46
rect 21 63 29 64
rect 21 59 23 63
rect 27 59 29 63
rect 21 38 29 59
rect 31 58 39 64
rect 31 54 33 58
rect 37 54 39 58
rect 31 50 39 54
rect 31 46 33 50
rect 37 46 39 50
rect 31 38 39 46
rect 41 63 49 64
rect 41 59 43 63
rect 47 59 49 63
rect 41 38 49 59
rect 51 50 59 64
rect 51 46 53 50
rect 57 46 59 50
rect 51 43 59 46
rect 51 39 53 43
rect 57 39 59 43
rect 51 38 59 39
rect 61 56 67 64
rect 83 56 91 60
rect 61 55 69 56
rect 61 51 63 55
rect 67 51 69 55
rect 61 38 69 51
rect 71 50 79 56
rect 71 46 73 50
rect 77 46 79 50
rect 71 43 79 46
rect 71 39 73 43
rect 77 39 79 43
rect 71 38 79 39
rect 81 55 91 56
rect 81 51 83 55
rect 87 51 91 55
rect 81 38 91 51
rect 93 50 101 60
rect 93 46 95 50
rect 99 46 101 50
rect 93 43 101 46
rect 93 39 95 43
rect 99 39 101 43
rect 93 38 101 39
rect 103 59 110 60
rect 103 55 105 59
rect 109 55 110 59
rect 103 38 110 55
<< metal1 >>
rect -2 68 114 72
rect -2 64 73 68
rect 77 64 114 68
rect 3 63 7 64
rect 3 58 7 59
rect 23 63 27 64
rect 43 63 47 64
rect 23 58 27 59
rect 33 58 38 59
rect 43 58 47 59
rect 13 57 17 58
rect 13 51 17 53
rect 2 50 17 51
rect 37 54 38 58
rect 33 50 38 54
rect 63 55 67 64
rect 83 55 87 64
rect 104 59 110 64
rect 104 55 105 59
rect 109 55 110 59
rect 63 50 67 51
rect 73 50 78 51
rect 83 50 87 51
rect 95 50 99 51
rect 2 46 13 50
rect 17 46 33 50
rect 37 46 53 50
rect 57 46 58 50
rect 2 18 6 46
rect 53 43 58 46
rect 25 38 49 42
rect 57 42 58 43
rect 77 46 78 50
rect 73 43 78 46
rect 57 39 73 42
rect 77 39 78 43
rect 95 43 99 46
rect 53 38 78 39
rect 82 39 95 42
rect 82 38 99 39
rect 10 34 14 35
rect 25 34 31 38
rect 45 34 49 38
rect 82 34 86 38
rect 106 34 110 51
rect 25 30 26 34
rect 30 30 31 34
rect 35 30 36 34
rect 40 30 41 34
rect 45 30 60 34
rect 64 30 71 34
rect 97 30 98 34
rect 102 30 110 34
rect 10 26 14 30
rect 35 26 41 30
rect 82 26 86 30
rect 10 25 100 26
rect 10 22 95 25
rect 94 21 95 22
rect 99 21 100 25
rect 105 20 109 21
rect 2 14 23 18
rect 27 14 63 18
rect 67 14 71 18
rect 81 14 82 18
rect 86 14 87 18
rect 81 11 87 14
rect 5 8 6 11
rect -2 7 6 8
rect 10 8 11 11
rect 42 8 43 11
rect 10 7 43 8
rect 47 8 48 11
rect 81 8 82 11
rect 47 7 82 8
rect 86 8 87 11
rect 105 8 109 16
rect 86 7 96 8
rect -2 4 96 7
rect 100 4 104 8
rect 108 4 114 8
rect -2 0 114 4
<< ntransistor >>
rect 12 6 14 26
rect 19 6 21 26
rect 29 6 31 26
rect 36 6 38 26
rect 52 6 54 26
rect 59 6 61 26
rect 69 6 71 26
rect 76 6 78 26
rect 91 15 93 26
rect 101 15 103 26
<< ptransistor >>
rect 9 38 11 64
rect 19 38 21 64
rect 29 38 31 64
rect 39 38 41 64
rect 49 38 51 64
rect 59 38 61 64
rect 69 38 71 56
rect 79 38 81 56
rect 91 38 93 60
rect 101 38 103 60
<< polycontact >>
rect 10 30 14 34
rect 26 30 30 34
rect 36 30 40 34
rect 60 30 64 34
rect 82 30 86 34
rect 98 30 102 34
<< ndcontact >>
rect 6 7 10 11
rect 23 14 27 18
rect 43 7 47 11
rect 63 14 67 18
rect 82 14 86 18
rect 95 21 99 25
rect 105 16 109 20
rect 82 7 86 11
<< pdcontact >>
rect 3 59 7 63
rect 13 53 17 57
rect 13 46 17 50
rect 23 59 27 63
rect 33 54 37 58
rect 33 46 37 50
rect 43 59 47 63
rect 53 46 57 50
rect 53 39 57 43
rect 63 51 67 55
rect 73 46 77 50
rect 73 39 77 43
rect 83 51 87 55
rect 95 46 99 50
rect 95 39 99 43
rect 105 55 109 59
<< psubstratepcontact >>
rect 96 4 100 8
rect 104 4 108 8
<< nsubstratencontact >>
rect 73 64 77 68
<< psubstratepdiff >>
rect 95 8 109 9
rect 95 4 96 8
rect 100 4 104 8
rect 108 4 109 8
rect 95 3 109 4
<< nsubstratendiff >>
rect 72 68 78 69
rect 72 64 73 68
rect 77 64 78 68
rect 72 63 78 64
<< labels >>
rlabel ntransistor 13 18 13 18 6 an
rlabel ntransistor 37 18 37 18 6 an
rlabel polycontact 83 32 83 32 6 an
rlabel metal1 12 16 12 16 6 z
rlabel metal1 12 28 12 28 6 an
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 48 12 48 6 z
rlabel metal1 28 16 28 16 6 z
rlabel metal1 36 16 36 16 6 z
rlabel metal1 20 16 20 16 6 z
rlabel metal1 38 28 38 28 6 an
rlabel metal1 36 40 36 40 6 b
rlabel metal1 28 36 28 36 6 b
rlabel metal1 20 48 20 48 6 z
rlabel metal1 36 52 36 52 6 z
rlabel metal1 28 48 28 48 6 z
rlabel metal1 56 4 56 4 6 vss
rlabel metal1 52 16 52 16 6 z
rlabel metal1 60 16 60 16 6 z
rlabel metal1 44 16 44 16 6 z
rlabel metal1 52 32 52 32 6 b
rlabel metal1 60 32 60 32 6 b
rlabel metal1 44 40 44 40 6 b
rlabel metal1 60 40 60 40 6 z
rlabel metal1 44 48 44 48 6 z
rlabel metal1 52 48 52 48 6 z
rlabel metal1 56 68 56 68 6 vdd
rlabel metal1 68 16 68 16 6 z
rlabel polycontact 84 32 84 32 6 an
rlabel metal1 68 32 68 32 6 b
rlabel metal1 68 40 68 40 6 z
rlabel pdcontact 76 48 76 48 6 z
rlabel ndcontact 97 23 97 23 6 an
rlabel polycontact 100 32 100 32 6 a
rlabel metal1 108 44 108 44 6 a
rlabel metal1 97 44 97 44 6 an
<< end >>
