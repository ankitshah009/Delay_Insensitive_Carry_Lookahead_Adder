magic
tech scmos
timestamp 1179387045
<< checkpaint >>
rect -22 -25 126 105
<< ab >>
rect 0 0 104 80
<< pwell >>
rect -4 -7 108 36
<< nwell >>
rect -4 36 108 87
<< polysilicon >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 36 70 38 74
rect 46 70 48 74
rect 53 70 55 74
rect 63 70 65 74
rect 70 70 72 74
rect 80 62 82 67
rect 87 62 89 67
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 9 38 21 39
rect 9 34 10 38
rect 14 34 21 38
rect 9 33 21 34
rect 25 38 31 39
rect 25 34 26 38
rect 30 34 31 38
rect 25 33 31 34
rect 36 33 38 42
rect 46 33 48 42
rect 53 39 55 42
rect 63 39 65 42
rect 70 39 72 42
rect 80 39 82 42
rect 53 38 65 39
rect 53 37 56 38
rect 55 34 56 37
rect 60 37 65 38
rect 69 38 82 39
rect 60 34 61 37
rect 55 33 61 34
rect 9 30 11 33
rect 19 30 21 33
rect 36 31 51 33
rect 39 28 41 31
rect 49 28 51 31
rect 59 28 61 33
rect 69 34 70 38
rect 74 37 82 38
rect 87 39 89 42
rect 87 38 95 39
rect 74 34 75 37
rect 69 33 75 34
rect 87 34 90 38
rect 94 34 95 38
rect 87 33 95 34
rect 69 28 71 33
rect 79 31 95 33
rect 79 28 81 31
rect 91 28 93 31
rect 29 22 31 27
rect 59 12 61 16
rect 9 6 11 11
rect 19 8 21 11
rect 29 8 31 11
rect 19 6 31 8
rect 39 6 41 11
rect 49 8 51 11
rect 69 8 71 16
rect 49 6 71 8
rect 79 6 81 11
rect 91 6 93 11
<< ndiffusion >>
rect 2 29 9 30
rect 2 25 3 29
rect 7 25 9 29
rect 2 22 9 25
rect 2 18 3 22
rect 7 18 9 22
rect 2 17 9 18
rect 4 11 9 17
rect 11 29 19 30
rect 11 25 13 29
rect 17 25 19 29
rect 11 11 19 25
rect 21 22 26 30
rect 34 22 39 28
rect 21 21 29 22
rect 21 17 23 21
rect 27 17 29 21
rect 21 11 29 17
rect 31 21 39 22
rect 31 17 33 21
rect 37 17 39 21
rect 31 11 39 17
rect 41 16 49 28
rect 41 12 43 16
rect 47 12 49 16
rect 41 11 49 12
rect 51 26 59 28
rect 51 22 53 26
rect 57 22 59 26
rect 51 16 59 22
rect 61 21 69 28
rect 61 17 63 21
rect 67 17 69 21
rect 61 16 69 17
rect 71 26 79 28
rect 71 22 73 26
rect 77 22 79 26
rect 71 16 79 22
rect 51 11 56 16
rect 74 11 79 16
rect 81 12 91 28
rect 81 11 84 12
rect 83 8 84 11
rect 88 11 91 12
rect 93 22 98 28
rect 93 21 100 22
rect 93 17 95 21
rect 99 17 100 21
rect 93 16 100 17
rect 93 11 98 16
rect 88 8 89 11
rect 83 7 89 8
<< pdiffusion >>
rect 2 69 9 70
rect 2 65 3 69
rect 7 65 9 69
rect 2 62 9 65
rect 2 58 3 62
rect 7 58 9 62
rect 2 42 9 58
rect 11 61 19 70
rect 11 57 13 61
rect 17 57 19 61
rect 11 54 19 57
rect 11 50 13 54
rect 17 50 19 54
rect 11 42 19 50
rect 21 69 29 70
rect 21 65 23 69
rect 27 65 29 69
rect 21 62 29 65
rect 21 58 23 62
rect 27 58 29 62
rect 21 42 29 58
rect 31 42 36 70
rect 38 61 46 70
rect 38 57 40 61
rect 44 57 46 61
rect 38 54 46 57
rect 38 50 40 54
rect 44 50 46 54
rect 38 42 46 50
rect 48 42 53 70
rect 55 69 63 70
rect 55 65 57 69
rect 61 65 63 69
rect 55 62 63 65
rect 55 58 57 62
rect 61 58 63 62
rect 55 42 63 58
rect 65 42 70 70
rect 72 62 77 70
rect 72 61 80 62
rect 72 57 74 61
rect 78 57 80 61
rect 72 54 80 57
rect 72 50 74 54
rect 78 50 80 54
rect 72 42 80 50
rect 82 42 87 62
rect 89 61 97 62
rect 89 57 91 61
rect 95 57 97 61
rect 89 54 97 57
rect 89 50 91 54
rect 95 50 97 54
rect 89 42 97 50
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect -2 69 106 78
rect -2 68 3 69
rect 2 65 3 68
rect 7 68 23 69
rect 7 65 8 68
rect 2 62 8 65
rect 22 65 23 68
rect 27 68 57 69
rect 27 65 28 68
rect 22 62 28 65
rect 56 65 57 68
rect 61 68 106 69
rect 61 65 62 68
rect 2 58 3 62
rect 7 58 8 62
rect 13 61 17 62
rect 22 58 23 62
rect 27 58 28 62
rect 40 61 46 63
rect 13 54 17 57
rect 44 57 46 61
rect 56 62 62 65
rect 56 58 57 62
rect 61 58 62 62
rect 73 61 79 63
rect 40 54 46 57
rect 73 57 74 61
rect 78 57 79 61
rect 73 54 79 57
rect 2 50 13 54
rect 17 50 40 54
rect 44 50 74 54
rect 78 50 79 54
rect 90 61 96 68
rect 90 57 91 61
rect 95 57 96 61
rect 90 54 96 57
rect 90 50 91 54
rect 95 50 96 54
rect 2 29 6 50
rect 10 42 23 46
rect 57 42 95 46
rect 10 38 14 42
rect 57 38 61 42
rect 89 38 95 42
rect 25 34 26 38
rect 30 34 56 38
rect 60 34 61 38
rect 65 34 70 38
rect 74 34 85 38
rect 89 34 90 38
rect 94 34 95 38
rect 10 33 14 34
rect 81 30 85 34
rect 2 25 3 29
rect 7 25 8 29
rect 12 25 13 29
rect 17 26 77 29
rect 81 26 95 30
rect 17 25 53 26
rect 2 22 8 25
rect 2 18 3 22
rect 7 21 8 22
rect 33 21 37 25
rect 57 25 73 26
rect 53 21 57 22
rect 73 21 77 22
rect 7 18 23 21
rect 2 17 23 18
rect 27 17 28 21
rect 62 17 63 21
rect 67 17 68 21
rect 73 17 95 21
rect 99 17 100 21
rect 33 16 37 17
rect 43 16 47 17
rect 62 12 68 17
rect -2 8 84 12
rect 88 8 106 12
rect -2 2 106 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
<< ntransistor >>
rect 9 11 11 30
rect 19 11 21 30
rect 29 11 31 22
rect 39 11 41 28
rect 49 11 51 28
rect 59 16 61 28
rect 69 16 71 28
rect 79 11 81 28
rect 91 11 93 28
<< ptransistor >>
rect 9 42 11 70
rect 19 42 21 70
rect 29 42 31 70
rect 36 42 38 70
rect 46 42 48 70
rect 53 42 55 70
rect 63 42 65 70
rect 70 42 72 70
rect 80 42 82 62
rect 87 42 89 62
<< polycontact >>
rect 10 34 14 38
rect 26 34 30 38
rect 56 34 60 38
rect 70 34 74 38
rect 90 34 94 38
<< ndcontact >>
rect 3 25 7 29
rect 3 18 7 22
rect 13 25 17 29
rect 23 17 27 21
rect 33 17 37 21
rect 43 12 47 16
rect 53 22 57 26
rect 63 17 67 21
rect 73 22 77 26
rect 84 8 88 12
rect 95 17 99 21
<< pdcontact >>
rect 3 65 7 69
rect 3 58 7 62
rect 13 57 17 61
rect 13 50 17 54
rect 23 65 27 69
rect 23 58 27 62
rect 40 57 44 61
rect 40 50 44 54
rect 57 65 61 69
rect 57 58 61 62
rect 74 57 78 61
rect 74 50 78 54
rect 91 57 95 61
rect 91 50 95 54
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
rect 90 -2 94 2
rect 98 -2 102 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
rect 90 78 94 82
rect 98 78 102 82
<< psubstratepdiff >>
rect 0 2 104 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 104 2
rect 0 -3 104 -2
<< nsubstratendiff >>
rect 0 82 104 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 104 82
rect 0 77 104 78
<< labels >>
rlabel metal1 4 32 4 32 6 z
rlabel polycontact 12 36 12 36 6 b
rlabel metal1 12 52 12 52 6 z
rlabel metal1 35 22 35 22 6 n1
rlabel metal1 20 44 20 44 6 b
rlabel polycontact 28 36 28 36 6 a1
rlabel metal1 36 36 36 36 6 a1
rlabel metal1 28 52 28 52 6 z
rlabel metal1 36 52 36 52 6 z
rlabel metal1 20 52 20 52 6 z
rlabel metal1 52 6 52 6 6 vss
rlabel metal1 44 36 44 36 6 a1
rlabel metal1 52 36 52 36 6 a1
rlabel metal1 60 44 60 44 6 a1
rlabel metal1 52 52 52 52 6 z
rlabel metal1 60 52 60 52 6 z
rlabel metal1 44 56 44 56 6 z
rlabel metal1 52 74 52 74 6 vdd
rlabel metal1 44 27 44 27 6 n1
rlabel ndcontact 75 23 75 23 6 n1
rlabel metal1 68 36 68 36 6 a2
rlabel metal1 68 44 68 44 6 a1
rlabel metal1 76 36 76 36 6 a2
rlabel metal1 76 44 76 44 6 a1
rlabel metal1 68 52 68 52 6 z
rlabel metal1 76 56 76 56 6 z
rlabel metal1 84 28 84 28 6 a2
rlabel metal1 86 19 86 19 6 n1
rlabel metal1 92 28 92 28 6 a2
rlabel metal1 84 44 84 44 6 a1
rlabel metal1 92 40 92 40 6 a1
<< end >>
