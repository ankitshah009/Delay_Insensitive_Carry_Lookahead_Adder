.subckt no3_x4 i0 i1 i2 nq vdd vss
*   SPICE3 file   created from no3_x4.ext -      technology: scmos
m00 w1     i2     w2     vdd p w=40u  l=2.3636u ad=120p     pd=46u      as=320p     ps=96u
m01 w3     i1     w1     vdd p w=40u  l=2.3636u ad=120p     pd=46u      as=120p     ps=46u
m02 vdd    i0     w3     vdd p w=40u  l=2.3636u ad=262.857p pd=59.4286u as=120p     ps=46u
m03 nq     w4     vdd    vdd p w=40u  l=2.3636u ad=200p     pd=50u      as=262.857p ps=59.4286u
m04 vdd    w4     nq     vdd p w=40u  l=2.3636u ad=262.857p pd=59.4286u as=200p     ps=50u
m05 w4     w2     vdd    vdd p w=20u  l=2.3636u ad=160p     pd=56u      as=131.429p ps=29.7143u
m06 vss    i2     w2     vss n w=10u  l=2.3636u ad=58.5p    pd=23u      as=60p      ps=25.3333u
m07 w2     i1     vss    vss n w=10u  l=2.3636u ad=60p      pd=25.3333u as=58.5p    ps=23u
m08 vss    i0     w2     vss n w=10u  l=2.3636u ad=58.5p    pd=23u      as=60p      ps=25.3333u
m09 nq     w4     vss    vss n w=20u  l=2.3636u ad=100p     pd=30u      as=117p     ps=46u
m10 vss    w4     nq     vss n w=20u  l=2.3636u ad=117p     pd=46u      as=100p     ps=30u
m11 w4     w2     vss    vss n w=10u  l=2.3636u ad=80p      pd=36u      as=58.5p    ps=23u
C0  w4     i1     0.043f
C1  vdd    i2     0.017f
C2  nq     w2     0.486f
C3  i0     i2     0.127f
C4  w1     w2     0.012f
C5  nq     w4     0.155f
C6  vss    i0     0.015f
C7  w3     vdd    0.014f
C8  vss    i2     0.015f
C9  nq     i1     0.056f
C10 w2     vdd    0.538f
C11 w3     i0     0.009f
C12 vdd    w4     0.019f
C13 w2     i0     0.389f
C14 w1     i1     0.018f
C15 vdd    i1     0.017f
C16 w4     i0     0.124f
C17 w2     i2     0.163f
C18 vss    w2     0.298f
C19 w4     i2     0.024f
C20 i0     i1     0.398f
C21 w3     w2     0.012f
C22 nq     vdd    0.036f
C23 vss    w4     0.074f
C24 i1     i2     0.436f
C25 nq     i0     0.095f
C26 vss    i1     0.015f
C27 w1     vdd    0.014f
C28 w2     w4     0.322f
C29 nq     i2     0.040f
C30 w3     i1     0.018f
C31 vss    nq     0.084f
C32 w1     i2     0.009f
C33 vdd    i0     0.044f
C34 w2     i1     0.185f
C36 nq     vss    0.018f
C37 w2     vss    0.039f
C39 w4     vss    0.069f
C40 i0     vss    0.037f
C41 i1     vss    0.032f
C42 i2     vss    0.031f
.ends
