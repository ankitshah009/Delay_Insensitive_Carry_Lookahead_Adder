magic
tech scmos
timestamp 1179387115
<< checkpaint >>
rect -22 -22 94 94
<< ab >>
rect 0 0 72 72
<< pwell >>
rect -4 -4 76 32
<< nwell >>
rect -4 32 76 76
<< polysilicon >>
rect 22 66 24 70
rect 29 66 31 70
rect 36 66 38 70
rect 46 66 48 70
rect 53 66 55 70
rect 60 66 62 70
rect 9 57 11 61
rect 9 35 11 38
rect 22 37 24 40
rect 19 36 25 37
rect 9 34 15 35
rect 9 30 10 34
rect 14 30 15 34
rect 9 29 15 30
rect 19 32 20 36
rect 24 32 25 36
rect 19 31 25 32
rect 29 31 31 40
rect 36 37 38 40
rect 46 37 48 40
rect 36 36 48 37
rect 36 35 41 36
rect 40 32 41 35
rect 45 35 48 36
rect 45 32 46 35
rect 40 31 46 32
rect 53 31 55 40
rect 60 37 62 40
rect 60 36 70 37
rect 60 35 65 36
rect 64 32 65 35
rect 69 32 70 36
rect 64 31 70 32
rect 9 26 11 29
rect 19 26 21 31
rect 29 30 35 31
rect 29 26 30 30
rect 34 26 35 30
rect 29 25 35 26
rect 40 22 42 31
rect 50 30 56 31
rect 50 26 51 30
rect 55 26 56 30
rect 50 25 56 26
rect 50 22 52 25
rect 9 5 11 10
rect 19 5 21 10
rect 40 2 42 6
rect 50 2 52 6
<< ndiffusion >>
rect 2 25 9 26
rect 2 21 3 25
rect 7 21 9 25
rect 2 18 9 21
rect 2 14 3 18
rect 7 14 9 18
rect 2 13 9 14
rect 4 10 9 13
rect 11 25 19 26
rect 11 21 13 25
rect 17 21 19 25
rect 11 18 19 21
rect 11 14 13 18
rect 17 14 19 18
rect 11 10 19 14
rect 21 22 26 26
rect 21 10 40 22
rect 23 8 40 10
rect 23 4 24 8
rect 28 4 33 8
rect 37 6 40 8
rect 42 17 50 22
rect 42 13 44 17
rect 48 13 50 17
rect 42 6 50 13
rect 52 18 59 22
rect 52 14 54 18
rect 58 14 59 18
rect 52 11 59 14
rect 52 7 54 11
rect 58 7 59 11
rect 52 6 59 7
rect 37 4 38 6
rect 23 3 38 4
<< pdiffusion >>
rect 13 65 22 66
rect 13 61 15 65
rect 19 61 22 65
rect 13 57 22 61
rect 2 56 9 57
rect 2 52 3 56
rect 7 52 9 56
rect 2 49 9 52
rect 2 45 3 49
rect 7 45 9 49
rect 2 44 9 45
rect 4 38 9 44
rect 11 40 22 57
rect 24 40 29 66
rect 31 40 36 66
rect 38 58 46 66
rect 38 54 40 58
rect 44 54 46 58
rect 38 40 46 54
rect 48 40 53 66
rect 55 40 60 66
rect 62 65 70 66
rect 62 61 64 65
rect 68 61 70 65
rect 62 58 70 61
rect 62 54 64 58
rect 68 54 70 58
rect 62 40 70 54
rect 11 38 16 40
<< metal1 >>
rect -2 68 74 72
rect -2 64 4 68
rect 8 65 74 68
rect 8 64 15 65
rect 14 61 15 64
rect 19 64 64 65
rect 19 61 20 64
rect 63 61 64 64
rect 68 64 74 65
rect 68 61 69 64
rect 63 58 69 61
rect 2 56 40 58
rect 2 52 3 56
rect 7 54 40 56
rect 44 54 47 58
rect 63 54 64 58
rect 68 54 69 58
rect 2 49 7 52
rect 2 45 3 49
rect 2 44 7 45
rect 10 46 23 50
rect 31 46 70 50
rect 2 25 6 44
rect 10 34 14 46
rect 31 42 35 46
rect 10 29 14 30
rect 18 38 35 42
rect 41 38 55 42
rect 18 36 24 38
rect 18 32 20 36
rect 18 29 24 32
rect 41 36 47 38
rect 45 32 47 36
rect 30 30 34 31
rect 41 30 47 32
rect 65 36 70 46
rect 69 32 70 36
rect 65 31 70 32
rect 51 30 55 31
rect 13 25 17 26
rect 2 21 3 25
rect 7 21 8 25
rect 2 18 8 21
rect 2 14 3 18
rect 7 14 8 18
rect 2 13 8 14
rect 30 22 70 26
rect 13 18 17 21
rect 17 14 44 17
rect 13 13 44 14
rect 48 13 49 17
rect 53 14 54 18
rect 58 14 59 18
rect 53 11 59 14
rect 66 13 70 22
rect 53 8 54 11
rect -2 4 24 8
rect 28 4 33 8
rect 37 7 54 8
rect 58 8 59 11
rect 58 7 64 8
rect 37 4 64 7
rect 68 4 74 8
rect -2 0 74 4
<< ntransistor >>
rect 9 10 11 26
rect 19 10 21 26
rect 40 6 42 22
rect 50 6 52 22
<< ptransistor >>
rect 9 38 11 57
rect 22 40 24 66
rect 29 40 31 66
rect 36 40 38 66
rect 46 40 48 66
rect 53 40 55 66
rect 60 40 62 66
<< polycontact >>
rect 10 30 14 34
rect 20 32 24 36
rect 41 32 45 36
rect 65 32 69 36
rect 30 26 34 30
rect 51 26 55 30
<< ndcontact >>
rect 3 21 7 25
rect 3 14 7 18
rect 13 21 17 25
rect 13 14 17 18
rect 24 4 28 8
rect 33 4 37 8
rect 44 13 48 17
rect 54 14 58 18
rect 54 7 58 11
<< pdcontact >>
rect 15 61 19 65
rect 3 52 7 56
rect 3 45 7 49
rect 40 54 44 58
rect 64 61 68 65
rect 64 54 68 58
<< psubstratepcontact >>
rect 64 4 68 8
<< nsubstratencontact >>
rect 4 64 8 68
<< psubstratepdiff >>
rect 63 8 69 24
rect 63 4 64 8
rect 68 4 69 8
rect 63 3 69 4
<< nsubstratendiff >>
rect 3 68 9 69
rect 3 64 4 68
rect 8 64 9 68
rect 3 63 9 64
<< labels >>
rlabel metal1 4 32 4 32 6 z
rlabel metal1 15 19 15 19 6 n3
rlabel metal1 20 32 20 32 6 a1
rlabel metal1 12 36 12 36 6 b
rlabel metal1 20 48 20 48 6 b
rlabel metal1 20 56 20 56 6 z
rlabel metal1 12 56 12 56 6 z
rlabel metal1 36 4 36 4 6 vss
rlabel metal1 36 24 36 24 6 a2
rlabel metal1 28 40 28 40 6 a1
rlabel metal1 36 48 36 48 6 a1
rlabel metal1 36 56 36 56 6 z
rlabel metal1 28 56 28 56 6 z
rlabel metal1 36 68 36 68 6 vdd
rlabel metal1 31 15 31 15 6 n3
rlabel metal1 44 24 44 24 6 a2
rlabel metal1 52 24 52 24 6 a2
rlabel metal1 44 36 44 36 6 a3
rlabel metal1 52 40 52 40 6 a3
rlabel metal1 44 48 44 48 6 a1
rlabel metal1 52 48 52 48 6 a1
rlabel metal1 44 56 44 56 6 z
rlabel metal1 68 16 68 16 6 a2
rlabel metal1 60 24 60 24 6 a2
rlabel metal1 68 40 68 40 6 a1
rlabel metal1 60 48 60 48 6 a1
<< end >>
