magic
tech scmos
timestamp 1179385308
<< checkpaint >>
rect -22 -25 118 105
<< ab >>
rect 0 0 96 80
<< pwell >>
rect -4 -7 100 36
<< nwell >>
rect -4 36 100 87
<< polysilicon >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 39 70 41 74
rect 49 70 51 74
rect 59 70 61 74
rect 69 70 71 74
rect 81 70 83 74
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 39 39 41 42
rect 49 39 51 42
rect 59 39 61 42
rect 69 39 71 42
rect 9 38 15 39
rect 9 34 10 38
rect 14 34 15 38
rect 9 33 15 34
rect 19 38 31 39
rect 19 34 23 38
rect 27 34 31 38
rect 19 33 31 34
rect 12 25 14 33
rect 19 25 21 33
rect 29 30 31 33
rect 36 38 42 39
rect 36 34 37 38
rect 41 34 42 38
rect 36 33 42 34
rect 49 38 55 39
rect 49 34 50 38
rect 54 34 55 38
rect 49 33 55 34
rect 59 38 71 39
rect 59 34 65 38
rect 69 34 71 38
rect 81 39 83 42
rect 81 38 87 39
rect 81 35 82 38
rect 59 33 71 34
rect 36 30 38 33
rect 52 30 54 33
rect 59 30 61 33
rect 69 30 71 33
rect 76 34 82 35
rect 86 34 87 38
rect 76 33 87 34
rect 76 30 78 33
rect 69 15 71 20
rect 76 15 78 20
rect 12 10 14 15
rect 19 10 21 15
rect 29 10 31 15
rect 36 10 38 15
rect 52 10 54 15
rect 59 10 61 15
<< ndiffusion >>
rect 24 25 29 30
rect 4 15 12 25
rect 14 15 19 25
rect 21 21 29 25
rect 21 17 23 21
rect 27 17 29 21
rect 21 15 29 17
rect 31 15 36 30
rect 38 20 52 30
rect 38 16 43 20
rect 47 16 52 20
rect 38 15 52 16
rect 54 15 59 30
rect 61 27 69 30
rect 61 23 63 27
rect 67 23 69 27
rect 61 20 69 23
rect 71 20 76 30
rect 78 25 88 30
rect 78 21 82 25
rect 86 21 88 25
rect 78 20 88 21
rect 61 15 66 20
rect 4 12 10 15
rect 4 8 5 12
rect 9 8 10 12
rect 4 7 10 8
<< pdiffusion >>
rect 73 71 79 72
rect 73 70 74 71
rect 4 64 9 70
rect 2 63 9 64
rect 2 59 3 63
rect 7 59 9 63
rect 2 58 9 59
rect 4 42 9 58
rect 11 54 19 70
rect 11 50 13 54
rect 17 50 19 54
rect 11 42 19 50
rect 21 63 29 70
rect 21 59 23 63
rect 27 59 29 63
rect 21 42 29 59
rect 31 54 39 70
rect 31 50 33 54
rect 37 50 39 54
rect 31 42 39 50
rect 41 62 49 70
rect 41 58 43 62
rect 47 58 49 62
rect 41 55 49 58
rect 41 51 43 55
rect 47 51 49 55
rect 41 42 49 51
rect 51 69 59 70
rect 51 65 53 69
rect 57 65 59 69
rect 51 62 59 65
rect 51 58 53 62
rect 57 58 59 62
rect 51 42 59 58
rect 61 62 69 70
rect 61 58 63 62
rect 67 58 69 62
rect 61 55 69 58
rect 61 51 63 55
rect 67 51 69 55
rect 61 42 69 51
rect 71 67 74 70
rect 78 70 79 71
rect 78 67 81 70
rect 71 42 81 67
rect 83 63 88 70
rect 83 62 90 63
rect 83 58 85 62
rect 89 58 90 62
rect 83 55 90 58
rect 83 51 85 55
rect 89 51 90 55
rect 83 50 90 51
rect 83 42 88 50
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect -2 71 98 78
rect -2 69 74 71
rect -2 68 53 69
rect 52 65 53 68
rect 57 68 74 69
rect 57 65 58 68
rect 73 67 74 68
rect 78 68 98 71
rect 78 67 79 68
rect 2 59 3 63
rect 7 59 23 63
rect 27 62 47 63
rect 27 59 43 62
rect 52 62 58 65
rect 52 58 53 62
rect 57 58 58 62
rect 63 62 89 63
rect 67 59 85 62
rect 43 55 47 58
rect 2 54 39 55
rect 2 50 13 54
rect 17 50 33 54
rect 37 50 39 54
rect 63 55 67 58
rect 85 55 89 58
rect 47 51 63 54
rect 43 50 67 51
rect 2 21 6 50
rect 74 46 78 55
rect 85 50 89 51
rect 10 42 42 46
rect 10 38 14 42
rect 36 38 42 42
rect 10 25 14 34
rect 18 34 23 38
rect 27 34 31 38
rect 36 34 37 38
rect 41 34 42 38
rect 49 42 86 46
rect 49 38 55 42
rect 82 38 86 42
rect 49 34 50 38
rect 54 34 55 38
rect 64 34 65 38
rect 69 34 78 38
rect 18 25 22 34
rect 33 27 67 30
rect 33 26 63 27
rect 33 21 39 26
rect 63 22 67 23
rect 2 17 23 21
rect 27 17 39 21
rect 43 20 47 21
rect 74 17 78 34
rect 82 33 86 34
rect 82 25 86 26
rect 43 12 47 16
rect 82 12 86 21
rect -2 8 5 12
rect 9 8 98 12
rect -2 2 98 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
<< ntransistor >>
rect 12 15 14 25
rect 19 15 21 25
rect 29 15 31 30
rect 36 15 38 30
rect 52 15 54 30
rect 59 15 61 30
rect 69 20 71 30
rect 76 20 78 30
<< ptransistor >>
rect 9 42 11 70
rect 19 42 21 70
rect 29 42 31 70
rect 39 42 41 70
rect 49 42 51 70
rect 59 42 61 70
rect 69 42 71 70
rect 81 42 83 70
<< polycontact >>
rect 10 34 14 38
rect 23 34 27 38
rect 37 34 41 38
rect 50 34 54 38
rect 65 34 69 38
rect 82 34 86 38
<< ndcontact >>
rect 23 17 27 21
rect 43 16 47 20
rect 63 23 67 27
rect 82 21 86 25
rect 5 8 9 12
<< pdcontact >>
rect 3 59 7 63
rect 13 50 17 54
rect 23 59 27 63
rect 33 50 37 54
rect 43 58 47 62
rect 43 51 47 55
rect 53 65 57 69
rect 53 58 57 62
rect 63 58 67 62
rect 63 51 67 55
rect 74 67 78 71
rect 85 58 89 62
rect 85 51 89 55
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
rect 90 -2 94 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
rect 90 78 94 82
<< psubstratepdiff >>
rect 0 2 96 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 96 2
rect 0 -3 96 -2
<< nsubstratendiff >>
rect 0 82 96 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 96 82
rect 0 77 96 78
<< labels >>
rlabel metal1 12 32 12 32 6 b1
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 52 12 52 6 z
rlabel metal1 20 28 20 28 6 b2
rlabel metal1 20 44 20 44 6 b1
rlabel metal1 28 36 28 36 6 b2
rlabel metal1 28 44 28 44 6 b1
rlabel metal1 28 52 28 52 6 z
rlabel metal1 20 52 20 52 6 z
rlabel metal1 48 6 48 6 6 vss
rlabel metal1 36 24 36 24 6 z
rlabel metal1 44 28 44 28 6 z
rlabel metal1 52 28 52 28 6 z
rlabel metal1 36 44 36 44 6 b1
rlabel metal1 52 40 52 40 6 a1
rlabel metal1 45 56 45 56 6 n3
rlabel pdcontact 36 52 36 52 6 z
rlabel pdcontact 24 61 24 61 6 n3
rlabel metal1 48 74 48 74 6 vdd
rlabel metal1 60 28 60 28 6 z
rlabel metal1 76 24 76 24 6 a2
rlabel metal1 60 44 60 44 6 a1
rlabel polycontact 68 36 68 36 6 a2
rlabel metal1 68 44 68 44 6 a1
rlabel metal1 76 48 76 48 6 a1
rlabel metal1 65 56 65 56 6 n3
rlabel polycontact 84 36 84 36 6 a1
rlabel metal1 87 56 87 56 6 n3
<< end >>
