.subckt nd2_x05 a b vdd vss z
*   SPICE3 file   created from nd2_x05.ext -      technology: scmos
m00 z      b      vdd    vdd p w=12u  l=2.3636u ad=60p      pd=22u      as=120p     ps=44u
m01 vdd    a      z      vdd p w=12u  l=2.3636u ad=120p     pd=44u      as=60p      ps=22u
m02 w1     b      z      vss n w=10u  l=2.3636u ad=30p      pd=16u      as=68p      ps=36u
m03 vss    a      w1     vss n w=10u  l=2.3636u ad=80p      pd=36u      as=30p      ps=16u
C0  w1     b      0.003f
C1  z      a      0.080f
C2  a      b      0.204f
C3  z      vdd    0.056f
C4  b      vdd    0.009f
C5  vss    z      0.032f
C6  vss    b      0.020f
C7  z      b      0.096f
C8  a      vdd    0.023f
C9  vss    a      0.003f
C11 z      vss    0.024f
C12 a      vss    0.033f
C13 b      vss    0.035f
.ends
