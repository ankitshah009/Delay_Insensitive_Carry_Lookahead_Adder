magic
tech scmos
timestamp 1180600696
<< checkpaint >>
rect -22 -22 92 122
<< ab >>
rect 0 0 70 100
<< pwell >>
rect -4 -4 74 48
<< nwell >>
rect -4 48 74 104
<< polysilicon >>
rect 11 94 13 98
rect 23 94 25 98
rect 35 94 37 98
rect 47 94 49 98
rect 11 43 13 55
rect 23 43 25 55
rect 7 42 13 43
rect 7 38 8 42
rect 12 38 13 42
rect 7 37 13 38
rect 17 42 25 43
rect 17 38 18 42
rect 22 38 25 42
rect 17 37 25 38
rect 11 25 13 37
rect 23 25 25 37
rect 35 43 37 55
rect 47 43 49 55
rect 35 42 43 43
rect 35 38 38 42
rect 42 38 43 42
rect 35 37 43 38
rect 47 42 53 43
rect 47 38 48 42
rect 52 38 53 42
rect 47 37 53 38
rect 35 25 37 37
rect 47 25 49 37
rect 11 2 13 6
rect 23 2 25 6
rect 35 2 37 6
rect 47 2 49 6
<< ndiffusion >>
rect 15 32 21 33
rect 15 28 16 32
rect 20 28 21 32
rect 15 25 21 28
rect 3 22 11 25
rect 3 18 4 22
rect 8 18 11 22
rect 3 6 11 18
rect 13 6 23 25
rect 25 22 35 25
rect 25 18 28 22
rect 32 18 35 22
rect 25 6 35 18
rect 37 12 47 25
rect 37 8 40 12
rect 44 8 47 12
rect 37 6 47 8
rect 49 22 57 25
rect 49 18 52 22
rect 56 18 57 22
rect 49 6 57 18
<< pdiffusion >>
rect 3 92 11 94
rect 3 88 4 92
rect 8 88 11 92
rect 3 55 11 88
rect 13 55 23 94
rect 25 82 35 94
rect 25 78 28 82
rect 32 78 35 82
rect 25 72 35 78
rect 25 68 28 72
rect 32 68 35 72
rect 25 62 35 68
rect 25 58 28 62
rect 32 58 35 62
rect 25 55 35 58
rect 37 55 47 94
rect 49 92 57 94
rect 49 88 52 92
rect 56 88 57 92
rect 49 73 57 88
rect 49 55 55 73
<< metal1 >>
rect -2 92 72 100
rect -2 88 4 92
rect 8 88 52 92
rect 56 88 72 92
rect 8 42 12 83
rect 8 37 12 38
rect 18 42 22 83
rect 18 37 22 38
rect 28 82 32 83
rect 28 72 32 78
rect 28 62 32 68
rect 28 32 32 58
rect 15 28 16 32
rect 20 28 32 32
rect 28 27 32 28
rect 38 42 42 83
rect 38 27 42 38
rect 48 42 52 83
rect 62 60 66 88
rect 62 55 66 56
rect 48 27 52 38
rect 3 18 4 22
rect 8 18 28 22
rect 32 18 52 22
rect 56 18 57 22
rect -2 8 40 12
rect 44 8 72 12
rect -2 0 72 8
<< ntransistor >>
rect 11 6 13 25
rect 23 6 25 25
rect 35 6 37 25
rect 47 6 49 25
<< ptransistor >>
rect 11 55 13 94
rect 23 55 25 94
rect 35 55 37 94
rect 47 55 49 94
<< polycontact >>
rect 8 38 12 42
rect 18 38 22 42
rect 38 38 42 42
rect 48 38 52 42
<< ndcontact >>
rect 16 28 20 32
rect 4 18 8 22
rect 28 18 32 22
rect 40 8 44 12
rect 52 18 56 22
<< pdcontact >>
rect 4 88 8 92
rect 28 78 32 82
rect 28 68 32 72
rect 28 58 32 62
rect 52 88 56 92
<< nsubstratencontact >>
rect 62 56 66 60
<< nsubstratendiff >>
rect 61 60 67 66
rect 61 56 62 60
rect 66 56 67 60
rect 61 55 67 56
<< labels >>
rlabel metal1 10 60 10 60 6 i0
rlabel metal1 20 30 20 30 6 nq
rlabel metal1 20 60 20 60 6 i1
rlabel metal1 30 55 30 55 6 nq
rlabel metal1 35 6 35 6 6 vss
rlabel metal1 40 55 40 55 6 i3
rlabel metal1 50 55 50 55 6 i2
rlabel metal1 35 94 35 94 6 vdd
<< end >>
