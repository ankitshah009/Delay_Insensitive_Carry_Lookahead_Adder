magic
tech scmos
timestamp 1179386337
<< checkpaint >>
rect -22 -22 118 94
<< ab >>
rect 0 0 96 72
<< pwell >>
rect -4 -4 100 32
<< nwell >>
rect -4 32 100 76
<< polysilicon >>
rect 9 64 11 69
rect 19 64 21 69
rect 29 64 31 69
rect 39 64 41 69
rect 49 64 51 69
rect 59 64 61 69
rect 69 56 71 61
rect 79 56 81 61
rect 9 35 11 38
rect 19 35 21 38
rect 29 35 31 38
rect 39 35 41 38
rect 9 34 15 35
rect 9 30 10 34
rect 14 30 15 34
rect 9 29 15 30
rect 19 34 31 35
rect 19 30 26 34
rect 30 30 31 34
rect 19 29 31 30
rect 35 34 41 35
rect 35 30 36 34
rect 40 31 41 34
rect 49 31 51 38
rect 59 35 61 38
rect 69 35 71 38
rect 79 35 81 38
rect 59 34 71 35
rect 40 30 54 31
rect 35 29 54 30
rect 12 26 14 29
rect 19 26 21 29
rect 29 26 31 29
rect 36 26 38 29
rect 52 26 54 29
rect 59 30 60 34
rect 64 30 71 34
rect 59 29 71 30
rect 75 34 81 35
rect 75 30 76 34
rect 80 30 81 34
rect 75 29 81 30
rect 59 26 61 29
rect 69 26 71 29
rect 76 26 78 29
rect 12 2 14 6
rect 19 2 21 6
rect 29 2 31 6
rect 36 2 38 6
rect 52 2 54 6
rect 59 2 61 6
rect 69 2 71 6
rect 76 2 78 6
<< ndiffusion >>
rect 3 11 12 26
rect 3 7 5 11
rect 9 7 12 11
rect 3 6 12 7
rect 14 6 19 26
rect 21 18 29 26
rect 21 14 23 18
rect 27 14 29 18
rect 21 6 29 14
rect 31 6 36 26
rect 38 11 52 26
rect 38 7 43 11
rect 47 7 52 11
rect 38 6 52 7
rect 54 6 59 26
rect 61 18 69 26
rect 61 14 63 18
rect 67 14 69 18
rect 61 6 69 14
rect 71 6 76 26
rect 78 18 86 26
rect 78 14 80 18
rect 84 14 86 18
rect 78 11 86 14
rect 78 7 80 11
rect 84 7 86 11
rect 78 6 86 7
<< pdiffusion >>
rect 2 63 9 64
rect 2 59 3 63
rect 7 59 9 63
rect 2 38 9 59
rect 11 57 19 64
rect 11 53 13 57
rect 17 53 19 57
rect 11 50 19 53
rect 11 46 13 50
rect 17 46 19 50
rect 11 38 19 46
rect 21 63 29 64
rect 21 59 23 63
rect 27 59 29 63
rect 21 38 29 59
rect 31 58 39 64
rect 31 54 33 58
rect 37 54 39 58
rect 31 50 39 54
rect 31 46 33 50
rect 37 46 39 50
rect 31 38 39 46
rect 41 63 49 64
rect 41 59 43 63
rect 47 59 49 63
rect 41 38 49 59
rect 51 50 59 64
rect 51 46 53 50
rect 57 46 59 50
rect 51 43 59 46
rect 51 39 53 43
rect 57 39 59 43
rect 51 38 59 39
rect 61 56 67 64
rect 61 55 69 56
rect 61 51 63 55
rect 67 51 69 55
rect 61 38 69 51
rect 71 50 79 56
rect 71 46 73 50
rect 77 46 79 50
rect 71 43 79 46
rect 71 39 73 43
rect 77 39 79 43
rect 71 38 79 39
rect 81 55 88 56
rect 81 51 83 55
rect 87 51 88 55
rect 81 38 88 51
<< metal1 >>
rect -2 68 98 72
rect -2 64 74 68
rect 78 64 82 68
rect 86 64 98 68
rect 3 63 7 64
rect 3 58 7 59
rect 23 63 27 64
rect 43 63 47 64
rect 23 58 27 59
rect 33 58 38 59
rect 43 58 47 59
rect 13 57 17 58
rect 13 51 17 53
rect 2 50 17 51
rect 37 54 38 58
rect 33 50 38 54
rect 63 55 67 64
rect 83 55 87 64
rect 63 50 67 51
rect 73 50 79 51
rect 83 50 87 51
rect 2 46 13 50
rect 17 46 33 50
rect 37 46 53 50
rect 57 46 58 50
rect 2 18 6 46
rect 53 43 58 46
rect 25 38 49 42
rect 57 42 58 43
rect 77 46 79 50
rect 73 43 79 46
rect 57 39 73 42
rect 77 39 79 43
rect 53 38 79 39
rect 10 34 14 35
rect 25 34 31 38
rect 45 34 49 38
rect 25 30 26 34
rect 30 30 31 34
rect 35 30 36 34
rect 40 30 41 34
rect 45 30 60 34
rect 64 30 65 34
rect 75 30 76 34
rect 80 30 81 34
rect 10 26 14 30
rect 35 26 41 30
rect 75 26 81 30
rect 10 22 87 26
rect 2 14 23 18
rect 27 14 63 18
rect 67 14 71 18
rect 79 14 80 18
rect 84 14 85 18
rect 79 11 85 14
rect 4 8 5 11
rect -2 7 5 8
rect 9 8 10 11
rect 42 8 43 11
rect 9 7 43 8
rect 47 8 48 11
rect 79 8 80 11
rect 47 7 80 8
rect 84 8 85 11
rect 84 7 98 8
rect -2 0 98 7
<< ntransistor >>
rect 12 6 14 26
rect 19 6 21 26
rect 29 6 31 26
rect 36 6 38 26
rect 52 6 54 26
rect 59 6 61 26
rect 69 6 71 26
rect 76 6 78 26
<< ptransistor >>
rect 9 38 11 64
rect 19 38 21 64
rect 29 38 31 64
rect 39 38 41 64
rect 49 38 51 64
rect 59 38 61 64
rect 69 38 71 56
rect 79 38 81 56
<< polycontact >>
rect 10 30 14 34
rect 26 30 30 34
rect 36 30 40 34
rect 60 30 64 34
rect 76 30 80 34
<< ndcontact >>
rect 5 7 9 11
rect 23 14 27 18
rect 43 7 47 11
rect 63 14 67 18
rect 80 14 84 18
rect 80 7 84 11
<< pdcontact >>
rect 3 59 7 63
rect 13 53 17 57
rect 13 46 17 50
rect 23 59 27 63
rect 33 54 37 58
rect 33 46 37 50
rect 43 59 47 63
rect 53 46 57 50
rect 53 39 57 43
rect 63 51 67 55
rect 73 46 77 50
rect 73 39 77 43
rect 83 51 87 55
<< nsubstratencontact >>
rect 74 64 78 68
rect 82 64 86 68
<< nsubstratendiff >>
rect 73 68 87 69
rect 73 64 74 68
rect 78 64 82 68
rect 86 64 87 68
rect 73 63 87 64
<< labels >>
rlabel metal1 12 16 12 16 6 z
rlabel polycontact 12 32 12 32 6 a
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 48 12 48 6 z
rlabel metal1 28 16 28 16 6 z
rlabel metal1 20 16 20 16 6 z
rlabel metal1 20 24 20 24 6 a
rlabel metal1 28 24 28 24 6 a
rlabel polycontact 28 32 28 32 6 b
rlabel metal1 28 36 28 36 6 b
rlabel metal1 20 48 20 48 6 z
rlabel metal1 28 48 28 48 6 z
rlabel metal1 48 4 48 4 6 vss
rlabel metal1 44 16 44 16 6 z
rlabel metal1 52 16 52 16 6 z
rlabel metal1 36 16 36 16 6 z
rlabel metal1 36 24 36 24 6 a
rlabel metal1 44 24 44 24 6 a
rlabel metal1 52 24 52 24 6 a
rlabel metal1 52 32 52 32 6 b
rlabel metal1 36 40 36 40 6 b
rlabel metal1 44 40 44 40 6 b
rlabel metal1 36 52 36 52 6 z
rlabel metal1 44 48 44 48 6 z
rlabel metal1 52 48 52 48 6 z
rlabel metal1 48 68 48 68 6 vdd
rlabel metal1 68 16 68 16 6 z
rlabel metal1 60 16 60 16 6 z
rlabel metal1 60 24 60 24 6 a
rlabel metal1 68 24 68 24 6 a
rlabel metal1 76 24 76 24 6 a
rlabel metal1 60 32 60 32 6 b
rlabel metal1 60 40 60 40 6 z
rlabel metal1 68 40 68 40 6 z
rlabel metal1 76 44 76 44 6 z
rlabel metal1 84 24 84 24 6 a
<< end >>
