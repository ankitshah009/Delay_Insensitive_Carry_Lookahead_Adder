magic
tech scmos
timestamp 1179386159
<< checkpaint >>
rect -22 -25 118 105
<< ab >>
rect 0 0 96 80
<< pwell >>
rect -4 -7 100 36
<< nwell >>
rect -4 36 100 87
<< polysilicon >>
rect 30 72 87 74
rect 20 64 22 69
rect 30 64 32 72
rect 40 64 42 68
rect 54 64 56 68
rect 9 55 11 60
rect 72 55 74 60
rect 85 60 87 72
rect 9 39 11 42
rect 20 39 22 42
rect 7 38 13 39
rect 7 34 8 38
rect 12 34 13 38
rect 7 33 13 34
rect 18 38 24 39
rect 30 38 32 42
rect 40 39 42 42
rect 54 39 56 42
rect 40 38 46 39
rect 18 34 19 38
rect 23 34 24 38
rect 40 34 41 38
rect 45 34 46 38
rect 18 33 24 34
rect 11 29 13 33
rect 22 29 24 33
rect 32 32 46 34
rect 52 38 61 39
rect 72 38 74 42
rect 52 34 56 38
rect 60 34 61 38
rect 52 33 61 34
rect 71 37 77 38
rect 71 33 72 37
rect 76 33 77 37
rect 85 36 87 50
rect 32 29 34 32
rect 11 15 13 19
rect 42 24 44 28
rect 52 27 54 33
rect 71 32 77 33
rect 81 35 87 36
rect 72 27 74 32
rect 81 31 82 35
rect 86 31 87 35
rect 81 30 87 31
rect 85 27 87 30
rect 22 13 24 18
rect 32 13 34 18
rect 42 8 44 13
rect 52 12 54 16
rect 72 12 74 17
rect 85 8 87 20
rect 42 6 87 8
<< ndiffusion >>
rect 4 28 11 29
rect 4 24 5 28
rect 9 24 11 28
rect 4 23 11 24
rect 6 19 11 23
rect 13 23 22 29
rect 13 19 16 23
rect 20 19 22 23
rect 15 18 22 19
rect 24 28 32 29
rect 24 24 26 28
rect 30 24 32 28
rect 24 18 32 24
rect 34 24 39 29
rect 47 24 52 27
rect 34 23 42 24
rect 34 19 36 23
rect 40 19 42 23
rect 34 18 42 19
rect 37 13 42 18
rect 44 23 52 24
rect 44 19 46 23
rect 50 19 52 23
rect 44 16 52 19
rect 54 21 61 27
rect 65 26 72 27
rect 65 22 66 26
rect 70 22 72 26
rect 65 21 72 22
rect 54 17 56 21
rect 60 17 61 21
rect 67 17 72 21
rect 74 20 85 27
rect 87 26 94 27
rect 87 22 89 26
rect 93 22 94 26
rect 87 20 94 22
rect 74 17 83 20
rect 54 16 61 17
rect 44 13 49 16
rect 77 15 83 17
rect 77 11 78 15
rect 82 11 83 15
rect 77 10 83 11
<< pdiffusion >>
rect 13 62 20 64
rect 13 58 14 62
rect 18 58 20 62
rect 13 55 20 58
rect 2 54 9 55
rect 2 50 3 54
rect 7 50 9 54
rect 2 49 9 50
rect 4 42 9 49
rect 11 42 20 55
rect 22 54 30 64
rect 22 50 24 54
rect 28 50 30 54
rect 22 42 30 50
rect 32 61 40 64
rect 32 57 34 61
rect 38 57 40 61
rect 32 54 40 57
rect 32 50 34 54
rect 38 50 40 54
rect 32 47 40 50
rect 32 43 34 47
rect 38 43 40 47
rect 32 42 40 43
rect 42 47 54 64
rect 42 43 48 47
rect 52 43 54 47
rect 42 42 54 43
rect 56 63 63 64
rect 56 59 58 63
rect 62 59 63 63
rect 76 63 83 64
rect 56 52 63 59
rect 76 59 77 63
rect 81 60 83 63
rect 81 59 85 60
rect 76 55 85 59
rect 56 42 61 52
rect 67 48 72 55
rect 65 47 72 48
rect 65 43 66 47
rect 70 43 72 47
rect 65 42 72 43
rect 74 50 85 55
rect 87 56 92 60
rect 87 55 94 56
rect 87 51 89 55
rect 93 51 94 55
rect 87 50 94 51
rect 74 42 83 50
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect -2 68 98 78
rect 13 62 19 68
rect 57 63 63 68
rect 13 58 14 62
rect 18 58 19 62
rect 25 61 38 62
rect 25 58 34 61
rect 57 59 58 63
rect 62 59 63 63
rect 76 63 82 68
rect 76 59 77 63
rect 81 59 82 63
rect 34 54 38 57
rect 2 50 3 54
rect 7 50 19 54
rect 23 50 24 54
rect 28 50 30 54
rect 2 39 6 47
rect 15 46 19 50
rect 15 42 23 46
rect 2 38 14 39
rect 2 34 8 38
rect 12 34 14 38
rect 2 33 14 34
rect 19 38 23 42
rect 19 30 23 34
rect 5 28 23 30
rect 9 26 23 28
rect 26 28 30 50
rect 5 23 9 24
rect 26 23 30 24
rect 34 47 38 50
rect 34 23 38 43
rect 41 51 89 55
rect 93 51 94 55
rect 41 38 45 51
rect 41 33 45 34
rect 48 47 52 48
rect 48 23 52 43
rect 64 47 70 48
rect 64 43 66 47
rect 64 42 70 43
rect 64 38 68 42
rect 55 34 56 38
rect 60 34 68 38
rect 74 41 86 47
rect 74 37 78 41
rect 15 19 16 23
rect 20 19 21 23
rect 34 19 36 23
rect 40 19 41 23
rect 45 19 46 23
rect 50 19 52 23
rect 64 27 68 34
rect 71 33 72 37
rect 76 33 78 37
rect 82 35 86 36
rect 64 26 70 27
rect 64 22 66 26
rect 82 22 86 31
rect 90 27 94 51
rect 56 21 60 22
rect 64 21 70 22
rect 15 12 21 19
rect 73 18 86 22
rect 89 26 94 27
rect 93 22 94 26
rect 89 21 94 22
rect 56 12 60 17
rect 77 12 78 15
rect -2 11 78 12
rect 82 12 83 15
rect 82 11 98 12
rect -2 2 98 11
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
<< ntransistor >>
rect 11 19 13 29
rect 22 18 24 29
rect 32 18 34 29
rect 42 13 44 24
rect 52 16 54 27
rect 72 17 74 27
rect 85 20 87 27
<< ptransistor >>
rect 9 42 11 55
rect 20 42 22 64
rect 30 42 32 64
rect 40 42 42 64
rect 54 42 56 64
rect 72 42 74 55
rect 85 50 87 60
<< polycontact >>
rect 8 34 12 38
rect 19 34 23 38
rect 41 34 45 38
rect 56 34 60 38
rect 72 33 76 37
rect 82 31 86 35
<< ndcontact >>
rect 5 24 9 28
rect 16 19 20 23
rect 26 24 30 28
rect 36 19 40 23
rect 46 19 50 23
rect 66 22 70 26
rect 56 17 60 21
rect 89 22 93 26
rect 78 11 82 15
<< pdcontact >>
rect 14 58 18 62
rect 3 50 7 54
rect 24 50 28 54
rect 34 57 38 61
rect 34 50 38 54
rect 34 43 38 47
rect 48 43 52 47
rect 58 59 62 63
rect 77 59 81 63
rect 66 43 70 47
rect 89 51 93 55
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
rect 90 -2 94 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
rect 90 78 94 82
<< psubstratepdiff >>
rect 0 2 96 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 96 2
rect 0 -3 96 -2
<< nsubstratendiff >>
rect 0 82 96 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 96 82
rect 0 77 96 78
<< labels >>
rlabel polycontact 21 36 21 36 6 a0n
rlabel polycontact 43 35 43 35 6 sn
rlabel polysilicon 56 36 56 36 6 a1n
rlabel metal1 4 40 4 40 6 a0
rlabel metal1 12 36 12 36 6 a0
rlabel metal1 14 28 14 28 6 a0n
rlabel polycontact 21 36 21 36 6 a0n
rlabel metal1 10 52 10 52 6 a0n
rlabel metal1 28 38 28 38 6 a0i
rlabel metal1 28 60 28 60 6 z
rlabel metal1 48 6 48 6 6 vss
rlabel metal1 36 40 36 40 6 z
rlabel metal1 43 44 43 44 6 sn
rlabel metal1 50 33 50 33 6 a1i
rlabel metal1 48 74 48 74 6 vdd
rlabel metal1 76 20 76 20 6 s
rlabel metal1 61 36 61 36 6 a1n
rlabel metal1 76 40 76 40 6 a1
rlabel metal1 66 34 66 34 6 a1n
rlabel metal1 84 28 84 28 6 s
rlabel metal1 84 44 84 44 6 a1
rlabel metal1 92 38 92 38 6 sn
rlabel metal1 67 53 67 53 6 sn
<< end >>
