magic
tech scmos
timestamp 1170759770
<< checkpaint >>
rect -22 -26 86 114
<< ab >>
rect 0 0 64 88
<< pwell >>
rect -4 -8 68 40
<< nwell >>
rect -4 40 68 96
<< polysilicon >>
rect 2 82 11 83
rect 2 78 6 82
rect 10 78 11 82
rect 2 77 11 78
rect 9 74 11 77
rect 21 77 30 83
rect 34 82 43 83
rect 34 78 38 82
rect 42 78 43 82
rect 34 77 43 78
rect 21 74 23 77
rect 41 74 43 77
rect 53 82 62 83
rect 53 78 54 82
rect 58 78 62 82
rect 53 77 62 78
rect 53 74 55 77
rect 9 43 11 46
rect 21 43 23 46
rect 41 43 43 46
rect 53 43 55 46
rect 2 37 14 43
rect 18 42 30 43
rect 18 38 22 42
rect 26 38 30 42
rect 18 37 30 38
rect 34 42 46 43
rect 34 38 35 42
rect 39 38 46 42
rect 34 37 46 38
rect 50 37 62 43
rect 9 34 11 37
rect 21 34 23 37
rect 41 34 43 37
rect 53 34 55 37
rect 9 11 11 14
rect 2 5 11 11
rect 21 11 23 14
rect 41 11 43 14
rect 21 5 30 11
rect 34 5 43 11
rect 53 11 55 14
rect 53 5 62 11
<< ndiffusion >>
rect 2 14 9 34
rect 11 26 21 34
rect 11 22 14 26
rect 18 22 21 26
rect 11 19 21 22
rect 11 15 14 19
rect 18 15 21 19
rect 11 14 21 15
rect 23 29 30 34
rect 23 25 25 29
rect 29 25 30 29
rect 23 22 30 25
rect 23 18 25 22
rect 29 18 30 22
rect 23 14 30 18
rect 34 19 41 34
rect 34 15 35 19
rect 39 15 41 19
rect 34 14 41 15
rect 43 30 53 34
rect 43 26 46 30
rect 50 26 53 30
rect 43 22 53 26
rect 43 18 46 22
rect 50 18 53 22
rect 43 14 53 18
rect 55 26 62 34
rect 55 22 57 26
rect 61 22 62 26
rect 55 19 62 22
rect 55 15 57 19
rect 61 15 62 19
rect 55 14 62 15
rect 13 2 19 14
rect 45 2 51 14
<< pdiffusion >>
rect 13 74 19 86
rect 45 74 51 86
rect 2 46 9 74
rect 11 73 21 74
rect 11 69 14 73
rect 18 69 21 73
rect 11 66 21 69
rect 11 62 14 66
rect 18 62 21 66
rect 11 46 21 62
rect 23 62 30 74
rect 23 58 25 62
rect 29 58 30 62
rect 23 55 30 58
rect 23 51 25 55
rect 29 51 30 55
rect 23 46 30 51
rect 34 73 41 74
rect 34 69 35 73
rect 39 69 41 73
rect 34 66 41 69
rect 34 62 35 66
rect 39 62 41 66
rect 34 46 41 62
rect 43 62 53 74
rect 43 58 46 62
rect 50 58 53 62
rect 43 54 53 58
rect 43 50 46 54
rect 50 50 53 54
rect 43 46 53 50
rect 55 72 62 74
rect 55 68 57 72
rect 61 68 62 72
rect 55 65 62 68
rect 55 61 57 65
rect 61 61 62 65
rect 55 46 62 61
<< metal1 >>
rect -2 86 2 90
rect 10 86 22 90
rect 30 86 34 90
rect 42 86 54 90
rect 62 86 66 90
rect 6 82 10 86
rect 6 77 10 78
rect 14 82 18 86
rect 37 78 38 82
rect 42 78 54 82
rect 58 78 59 82
rect 14 73 18 78
rect 18 69 35 73
rect 39 72 61 73
rect 39 69 57 72
rect 14 66 18 69
rect 35 66 39 69
rect 14 61 18 62
rect 22 62 29 63
rect 22 58 25 62
rect 57 65 61 68
rect 35 61 39 62
rect 46 62 50 63
rect 22 57 29 58
rect 25 55 29 57
rect 14 38 18 55
rect 57 60 61 61
rect 46 54 50 58
rect 29 51 46 54
rect 25 50 46 51
rect 22 42 26 43
rect 35 42 39 43
rect 14 34 39 38
rect 14 33 18 34
rect 46 30 50 50
rect 25 29 46 30
rect 14 26 18 27
rect 29 26 46 29
rect 25 23 29 25
rect 14 19 18 22
rect 22 22 29 23
rect 22 18 25 22
rect 46 22 50 26
rect 22 17 29 18
rect 35 19 39 20
rect 14 10 18 15
rect 14 2 18 6
rect 46 17 50 18
rect 57 26 61 27
rect 57 19 61 22
rect 35 10 39 15
rect 35 2 39 6
rect 57 10 61 15
rect 57 2 61 6
rect -2 -2 2 2
rect 10 -2 22 2
rect 30 -2 34 2
rect 42 -2 54 2
rect 62 -2 66 2
<< metal2 >>
rect -2 86 6 90
rect 10 86 22 90
rect 26 86 38 90
rect 42 86 54 90
rect 58 86 66 90
rect -2 82 66 86
rect -2 78 14 82
rect 18 78 66 82
rect -2 76 66 78
rect -2 10 66 12
rect -2 6 14 10
rect 18 6 35 10
rect 39 6 57 10
rect 61 6 66 10
rect -2 2 66 6
rect -2 -2 6 2
rect 10 -2 22 2
rect 26 -2 38 2
rect 42 -2 54 2
rect 58 -2 66 2
<< ntransistor >>
rect 9 14 11 34
rect 21 14 23 34
rect 41 14 43 34
rect 53 14 55 34
<< ptransistor >>
rect 9 46 11 74
rect 21 46 23 74
rect 41 46 43 74
rect 53 46 55 74
<< polycontact >>
rect 6 78 10 82
rect 38 78 42 82
rect 54 78 58 82
rect 22 38 26 42
rect 35 38 39 42
<< ndcontact >>
rect 14 22 18 26
rect 14 15 18 19
rect 25 25 29 29
rect 25 18 29 22
rect 35 15 39 19
rect 46 26 50 30
rect 46 18 50 22
rect 57 22 61 26
rect 57 15 61 19
<< pdcontact >>
rect 14 69 18 73
rect 14 62 18 66
rect 25 58 29 62
rect 25 51 29 55
rect 35 69 39 73
rect 35 62 39 66
rect 46 58 50 62
rect 46 50 50 54
rect 57 68 61 72
rect 57 61 61 65
<< m2contact >>
rect 6 86 10 90
rect 22 86 26 90
rect 38 86 42 90
rect 54 86 58 90
rect 14 78 18 82
rect 14 6 18 10
rect 35 6 39 10
rect 57 6 61 10
rect 6 -2 10 2
rect 22 -2 26 2
rect 38 -2 42 2
rect 54 -2 58 2
<< psubstratepcontact >>
rect 2 -2 6 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 58 -2 62 2
<< nsubstratencontact >>
rect 2 86 6 90
rect 26 86 30 90
rect 34 86 38 90
rect 58 86 62 90
<< psubstratepdiff >>
rect 0 2 7 3
rect 25 2 39 3
rect 57 2 64 3
rect 0 -2 2 2
rect 6 -2 7 2
rect 0 -3 7 -2
rect 25 -2 26 2
rect 30 -2 34 2
rect 38 -2 39 2
rect 25 -3 39 -2
rect 57 -2 58 2
rect 62 -2 64 2
rect 57 -3 64 -2
<< nsubstratendiff >>
rect 0 90 7 91
rect 0 86 2 90
rect 6 86 7 90
rect 25 90 39 91
rect 25 86 26 90
rect 30 86 34 90
rect 38 86 39 90
rect 57 90 64 91
rect 57 86 58 90
rect 62 86 64 90
rect 0 85 7 86
rect 25 85 39 86
rect 57 85 64 86
<< labels >>
rlabel metal1 16 44 16 44 6 a
rlabel metal1 24 20 24 20 6 z
rlabel metal1 32 28 32 28 6 z
rlabel metal1 32 36 32 36 6 a
rlabel metal1 24 36 24 36 6 a
rlabel metal1 32 52 32 52 6 z
rlabel metal1 24 60 24 60 6 z
rlabel metal1 40 28 40 28 6 z
rlabel metal1 48 40 48 40 6 z
rlabel metal1 40 52 40 52 6 z
rlabel metal2 32 6 32 6 6 vss
rlabel metal2 32 82 32 82 6 vdd
<< end >>
