magic
tech scmos
timestamp 1179385708
<< checkpaint >>
rect -22 -25 150 105
<< ab >>
rect 0 0 128 80
<< pwell >>
rect -4 -7 132 36
<< nwell >>
rect -4 36 132 87
<< polysilicon >>
rect 19 70 21 74
rect 29 70 31 74
rect 39 70 41 74
rect 49 70 51 74
rect 59 70 61 74
rect 71 70 73 74
rect 78 70 80 74
rect 88 70 90 74
rect 95 70 97 74
rect 107 70 109 74
rect 117 70 119 74
rect 9 58 11 63
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 9 38 21 39
rect 9 34 10 38
rect 14 34 21 38
rect 9 33 21 34
rect 25 38 31 39
rect 25 34 26 38
rect 30 34 31 38
rect 25 33 31 34
rect 9 30 11 33
rect 19 27 21 33
rect 29 30 31 33
rect 39 39 41 42
rect 49 39 51 42
rect 39 38 51 39
rect 39 34 40 38
rect 44 34 51 38
rect 39 33 51 34
rect 39 30 41 33
rect 49 30 51 33
rect 59 39 61 42
rect 71 39 73 42
rect 59 38 73 39
rect 59 34 62 38
rect 66 34 73 38
rect 59 33 73 34
rect 59 30 61 33
rect 71 30 73 33
rect 78 39 80 42
rect 88 39 90 42
rect 78 38 90 39
rect 78 34 85 38
rect 89 34 90 38
rect 78 33 90 34
rect 78 30 80 33
rect 88 30 90 33
rect 95 39 97 42
rect 107 39 109 42
rect 117 39 119 42
rect 95 38 103 39
rect 95 34 98 38
rect 102 34 103 38
rect 95 33 103 34
rect 107 38 119 39
rect 107 34 114 38
rect 118 34 119 38
rect 107 33 119 34
rect 95 30 97 33
rect 107 30 109 33
rect 117 30 119 33
rect 9 15 11 19
rect 19 11 21 16
rect 29 11 31 16
rect 39 11 41 16
rect 49 11 51 16
rect 59 11 61 16
rect 88 15 90 19
rect 95 15 97 19
rect 71 8 73 13
rect 78 8 80 13
rect 107 11 109 16
rect 117 11 119 16
<< ndiffusion >>
rect 2 24 9 30
rect 2 20 3 24
rect 7 20 9 24
rect 2 19 9 20
rect 11 27 16 30
rect 23 27 29 30
rect 11 26 19 27
rect 11 22 13 26
rect 17 22 19 26
rect 11 19 19 22
rect 14 16 19 19
rect 21 21 29 27
rect 21 17 23 21
rect 27 17 29 21
rect 21 16 29 17
rect 31 21 39 30
rect 31 17 33 21
rect 37 17 39 21
rect 31 16 39 17
rect 41 29 49 30
rect 41 25 43 29
rect 47 25 49 29
rect 41 16 49 25
rect 51 21 59 30
rect 51 17 53 21
rect 57 17 59 21
rect 51 16 59 17
rect 61 16 71 30
rect 63 13 71 16
rect 73 13 78 30
rect 80 29 88 30
rect 80 25 82 29
rect 86 25 88 29
rect 80 19 88 25
rect 90 19 95 30
rect 97 19 107 30
rect 80 13 85 19
rect 99 16 107 19
rect 109 21 117 30
rect 109 17 111 21
rect 115 17 117 21
rect 109 16 117 17
rect 119 28 126 30
rect 119 24 121 28
rect 125 24 126 28
rect 119 21 126 24
rect 119 17 121 21
rect 125 17 126 21
rect 119 16 126 17
rect 63 12 69 13
rect 63 8 64 12
rect 68 8 69 12
rect 99 12 105 16
rect 99 8 100 12
rect 104 8 105 12
rect 63 7 69 8
rect 99 7 105 8
<< pdiffusion >>
rect 14 58 19 70
rect 2 57 9 58
rect 2 53 3 57
rect 7 53 9 57
rect 2 42 9 53
rect 11 54 19 58
rect 11 50 13 54
rect 17 50 19 54
rect 11 47 19 50
rect 11 43 13 47
rect 17 43 19 47
rect 11 42 19 43
rect 21 69 29 70
rect 21 65 23 69
rect 27 65 29 69
rect 21 62 29 65
rect 21 58 23 62
rect 27 58 29 62
rect 21 42 29 58
rect 31 62 39 70
rect 31 58 33 62
rect 37 58 39 62
rect 31 42 39 58
rect 41 47 49 70
rect 41 43 43 47
rect 47 43 49 47
rect 41 42 49 43
rect 51 62 59 70
rect 51 58 53 62
rect 57 58 59 62
rect 51 42 59 58
rect 61 69 71 70
rect 61 65 64 69
rect 68 65 71 69
rect 61 42 71 65
rect 73 42 78 70
rect 80 47 88 70
rect 80 43 82 47
rect 86 43 88 47
rect 80 42 88 43
rect 90 42 95 70
rect 97 69 107 70
rect 97 65 100 69
rect 104 65 107 69
rect 97 42 107 65
rect 109 62 117 70
rect 109 58 111 62
rect 115 58 117 62
rect 109 55 117 58
rect 109 51 111 55
rect 115 51 117 55
rect 109 42 117 51
rect 119 69 126 70
rect 119 65 121 69
rect 125 65 126 69
rect 119 61 126 65
rect 119 57 121 61
rect 125 57 126 61
rect 119 42 126 57
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect 118 78 122 82
rect 126 78 130 82
rect -2 69 130 78
rect -2 68 23 69
rect 3 57 7 68
rect 27 68 64 69
rect 63 65 64 68
rect 68 68 100 69
rect 68 65 69 68
rect 99 65 100 68
rect 104 68 121 69
rect 104 65 105 68
rect 125 68 130 69
rect 23 62 27 65
rect 32 58 33 62
rect 37 58 53 62
rect 57 58 111 62
rect 115 58 116 62
rect 23 57 27 58
rect 111 55 116 58
rect 121 61 125 65
rect 121 56 125 57
rect 3 52 7 53
rect 13 54 17 55
rect 13 47 17 50
rect 2 39 6 47
rect 26 50 103 54
rect 115 51 116 55
rect 111 50 116 51
rect 17 43 22 46
rect 13 42 22 43
rect 2 38 14 39
rect 2 34 10 38
rect 2 33 14 34
rect 18 29 22 42
rect 26 38 30 50
rect 42 46 43 47
rect 41 43 43 46
rect 47 46 48 47
rect 47 43 55 46
rect 41 42 55 43
rect 26 33 30 34
rect 34 34 40 38
rect 44 34 45 38
rect 34 29 38 34
rect 50 30 55 42
rect 62 38 66 50
rect 81 46 82 47
rect 62 33 66 34
rect 73 43 82 46
rect 86 43 87 47
rect 73 42 87 43
rect 97 42 103 50
rect 73 30 78 42
rect 98 38 102 42
rect 84 34 85 38
rect 89 30 95 38
rect 98 33 102 34
rect 114 38 118 39
rect 114 30 118 34
rect 13 26 38 29
rect 41 29 86 30
rect 41 26 43 29
rect 3 24 7 25
rect 17 25 38 26
rect 42 25 43 26
rect 47 26 82 29
rect 47 25 48 26
rect 73 25 82 26
rect 89 26 118 30
rect 121 28 125 29
rect 73 24 86 25
rect 13 21 17 22
rect 23 21 27 22
rect 121 21 125 24
rect 3 12 7 20
rect 32 17 33 21
rect 37 17 53 21
rect 57 17 111 21
rect 115 17 116 21
rect 23 12 27 17
rect 121 12 125 17
rect -2 8 64 12
rect 68 8 100 12
rect 104 8 130 12
rect -2 2 130 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 122 2
rect 126 -2 130 2
<< ntransistor >>
rect 9 19 11 30
rect 19 16 21 27
rect 29 16 31 30
rect 39 16 41 30
rect 49 16 51 30
rect 59 16 61 30
rect 71 13 73 30
rect 78 13 80 30
rect 88 19 90 30
rect 95 19 97 30
rect 107 16 109 30
rect 117 16 119 30
<< ptransistor >>
rect 9 42 11 58
rect 19 42 21 70
rect 29 42 31 70
rect 39 42 41 70
rect 49 42 51 70
rect 59 42 61 70
rect 71 42 73 70
rect 78 42 80 70
rect 88 42 90 70
rect 95 42 97 70
rect 107 42 109 70
rect 117 42 119 70
<< polycontact >>
rect 10 34 14 38
rect 26 34 30 38
rect 40 34 44 38
rect 62 34 66 38
rect 85 34 89 38
rect 98 34 102 38
rect 114 34 118 38
<< ndcontact >>
rect 3 20 7 24
rect 13 22 17 26
rect 23 17 27 21
rect 33 17 37 21
rect 43 25 47 29
rect 53 17 57 21
rect 82 25 86 29
rect 111 17 115 21
rect 121 24 125 28
rect 121 17 125 21
rect 64 8 68 12
rect 100 8 104 12
<< pdcontact >>
rect 3 53 7 57
rect 13 50 17 54
rect 13 43 17 47
rect 23 65 27 69
rect 23 58 27 62
rect 33 58 37 62
rect 43 43 47 47
rect 53 58 57 62
rect 64 65 68 69
rect 82 43 86 47
rect 100 65 104 69
rect 111 58 115 62
rect 111 51 115 55
rect 121 65 125 69
rect 121 57 125 61
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
rect 90 -2 94 2
rect 98 -2 102 2
rect 106 -2 110 2
rect 114 -2 118 2
rect 122 -2 126 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
rect 90 78 94 82
rect 98 78 102 82
rect 106 78 110 82
rect 114 78 118 82
rect 122 78 126 82
<< psubstratepdiff >>
rect 0 2 128 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 122 2
rect 126 -2 128 2
rect 0 -3 128 -2
<< nsubstratendiff >>
rect 0 82 128 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect 118 78 122 82
rect 126 78 128 82
rect 0 77 128 78
<< labels >>
rlabel polysilicon 45 36 45 36 6 cn
rlabel metal1 4 40 4 40 6 c
rlabel polycontact 12 36 12 36 6 c
rlabel metal1 15 48 15 48 6 cn
rlabel metal1 25 27 25 27 6 cn
rlabel ndcontact 44 28 44 28 6 z
rlabel metal1 39 36 39 36 6 cn
rlabel metal1 28 40 28 40 6 a
rlabel pdcontact 44 44 44 44 6 z
rlabel metal1 36 52 36 52 6 a
rlabel metal1 44 52 44 52 6 a
rlabel metal1 64 6 64 6 6 vss
rlabel metal1 60 28 60 28 6 z
rlabel metal1 68 28 68 28 6 z
rlabel metal1 52 36 52 36 6 z
rlabel metal1 60 52 60 52 6 a
rlabel metal1 68 52 68 52 6 a
rlabel metal1 52 52 52 52 6 a
rlabel metal1 64 74 64 74 6 vdd
rlabel metal1 100 28 100 28 6 b
rlabel metal1 92 32 92 32 6 b
rlabel metal1 76 36 76 36 6 z
rlabel pdcontact 84 44 84 44 6 z
rlabel metal1 100 48 100 48 6 a
rlabel metal1 84 52 84 52 6 a
rlabel metal1 92 52 92 52 6 a
rlabel metal1 76 52 76 52 6 a
rlabel metal1 74 19 74 19 6 n3
rlabel metal1 108 28 108 28 6 b
rlabel polycontact 116 36 116 36 6 b
rlabel metal1 113 56 113 56 6 n1
rlabel metal1 74 60 74 60 6 n1
<< end >>
