magic
tech scmos
timestamp 1180600719
<< checkpaint >>
rect -22 -22 102 122
<< ab >>
rect 0 0 80 100
<< pwell >>
rect -4 -4 84 48
<< nwell >>
rect -4 48 84 104
<< polysilicon >>
rect 11 94 13 98
rect 19 94 21 98
rect 27 94 29 98
rect 43 94 45 98
rect 55 94 57 98
rect 11 33 13 56
rect 19 43 21 56
rect 27 53 29 56
rect 67 76 69 80
rect 27 52 33 53
rect 27 48 28 52
rect 32 49 33 52
rect 32 48 37 49
rect 27 47 37 48
rect 17 42 23 43
rect 17 38 18 42
rect 22 38 23 42
rect 17 37 23 38
rect 7 32 13 33
rect 7 28 8 32
rect 12 28 13 32
rect 7 27 13 28
rect 19 29 21 37
rect 19 27 25 29
rect 11 24 13 27
rect 23 24 25 27
rect 35 25 37 47
rect 43 43 45 55
rect 55 43 57 55
rect 67 53 69 56
rect 61 52 69 53
rect 61 48 62 52
rect 66 48 69 52
rect 61 47 69 48
rect 43 42 63 43
rect 43 38 58 42
rect 62 38 63 42
rect 43 37 63 38
rect 45 25 47 37
rect 57 25 59 37
rect 67 25 69 47
rect 11 10 13 14
rect 23 10 25 14
rect 35 11 37 15
rect 67 11 69 15
rect 45 2 47 6
rect 57 2 59 6
<< ndiffusion >>
rect 30 24 35 25
rect 3 22 11 24
rect 3 18 4 22
rect 8 18 11 22
rect 3 14 11 18
rect 13 14 23 24
rect 25 22 35 24
rect 25 18 28 22
rect 32 18 35 22
rect 25 15 35 18
rect 37 15 45 25
rect 25 14 33 15
rect 15 12 21 14
rect 15 8 16 12
rect 20 8 21 12
rect 39 9 45 15
rect 15 7 21 8
rect 37 8 45 9
rect 37 4 38 8
rect 42 6 45 8
rect 47 22 57 25
rect 47 18 50 22
rect 54 18 57 22
rect 47 6 57 18
rect 59 15 67 25
rect 69 22 77 25
rect 69 18 72 22
rect 76 18 77 22
rect 69 15 77 18
rect 59 9 65 15
rect 59 8 67 9
rect 59 6 62 8
rect 42 4 43 6
rect 37 3 43 4
rect 61 4 62 6
rect 66 4 67 8
rect 61 3 67 4
<< pdiffusion >>
rect 3 82 11 94
rect 3 78 4 82
rect 8 78 11 82
rect 3 56 11 78
rect 13 56 19 94
rect 21 56 27 94
rect 29 92 43 94
rect 29 88 36 92
rect 40 88 43 92
rect 29 56 43 88
rect 35 55 43 56
rect 45 72 55 94
rect 45 68 48 72
rect 52 68 55 72
rect 45 62 55 68
rect 45 58 48 62
rect 52 58 55 62
rect 45 55 55 58
rect 57 92 65 94
rect 57 88 60 92
rect 64 88 65 92
rect 57 76 65 88
rect 57 56 67 76
rect 69 62 77 76
rect 69 58 72 62
rect 76 58 77 62
rect 69 56 77 58
rect 57 55 62 56
<< metal1 >>
rect -2 96 82 100
rect -2 92 72 96
rect 76 92 82 96
rect -2 88 36 92
rect 40 88 60 92
rect 64 88 82 92
rect 3 78 4 82
rect 8 78 66 82
rect 8 32 12 73
rect 8 27 12 28
rect 18 42 22 73
rect 18 27 22 38
rect 28 52 32 73
rect 28 27 32 48
rect 38 22 42 78
rect 3 18 4 22
rect 8 18 28 22
rect 32 18 42 22
rect 48 72 52 73
rect 48 62 52 68
rect 48 22 52 58
rect 62 52 66 78
rect 62 47 66 48
rect 72 62 76 63
rect 72 42 76 58
rect 57 38 58 42
rect 62 38 76 42
rect 72 22 76 38
rect 48 18 50 22
rect 54 18 55 22
rect 48 17 52 18
rect 72 17 76 18
rect -2 8 16 12
rect 20 8 82 12
rect -2 4 38 8
rect 42 4 62 8
rect 66 4 82 8
rect -2 0 82 4
<< ntransistor >>
rect 11 14 13 24
rect 23 14 25 24
rect 35 15 37 25
rect 45 6 47 25
rect 57 6 59 25
rect 67 15 69 25
<< ptransistor >>
rect 11 56 13 94
rect 19 56 21 94
rect 27 56 29 94
rect 43 55 45 94
rect 55 55 57 94
rect 67 56 69 76
<< polycontact >>
rect 28 48 32 52
rect 18 38 22 42
rect 8 28 12 32
rect 62 48 66 52
rect 58 38 62 42
<< ndcontact >>
rect 4 18 8 22
rect 28 18 32 22
rect 16 8 20 12
rect 38 4 42 8
rect 50 18 54 22
rect 72 18 76 22
rect 62 4 66 8
<< pdcontact >>
rect 4 78 8 82
rect 36 88 40 92
rect 48 68 52 72
rect 48 58 52 62
rect 60 88 64 92
rect 72 58 76 62
<< nsubstratencontact >>
rect 72 92 76 96
<< nsubstratendiff >>
rect 71 96 77 97
rect 71 92 72 96
rect 76 92 77 96
rect 71 86 77 92
<< labels >>
rlabel metal1 10 50 10 50 6 i2
rlabel polycontact 30 50 30 50 6 i0
rlabel metal1 20 50 20 50 6 i1
rlabel ndcontact 40 6 40 6 6 vss
rlabel metal1 50 45 50 45 6 nq
rlabel metal1 40 94 40 94 6 vdd
<< end >>
