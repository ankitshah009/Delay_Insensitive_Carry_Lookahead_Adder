magic
tech scmos
timestamp 1179387127
<< checkpaint >>
rect -22 -25 158 105
<< ab >>
rect 0 0 136 80
<< pwell >>
rect -4 -7 140 36
<< nwell >>
rect -4 36 140 87
<< polysilicon >>
rect 31 70 33 74
rect 39 70 41 74
rect 47 70 49 74
rect 57 70 59 74
rect 65 70 67 74
rect 73 70 75 74
rect 83 70 85 74
rect 91 70 93 74
rect 99 70 101 74
rect 109 70 111 74
rect 116 70 118 74
rect 123 70 125 74
rect 9 61 11 65
rect 19 63 21 68
rect 9 39 11 42
rect 19 39 21 42
rect 31 39 33 42
rect 39 39 41 42
rect 47 39 49 42
rect 57 39 59 42
rect 65 39 67 42
rect 73 39 75 42
rect 83 39 85 42
rect 91 39 93 42
rect 99 39 101 42
rect 109 39 111 42
rect 9 38 21 39
rect 9 34 13 38
rect 17 34 21 38
rect 9 33 21 34
rect 26 38 33 39
rect 26 34 27 38
rect 31 34 33 38
rect 26 33 33 34
rect 37 38 43 39
rect 37 34 38 38
rect 42 34 43 38
rect 47 38 59 39
rect 47 37 50 38
rect 37 33 43 34
rect 49 34 50 37
rect 54 37 59 38
rect 63 38 69 39
rect 54 34 55 37
rect 49 33 55 34
rect 63 34 64 38
rect 68 34 69 38
rect 63 33 69 34
rect 73 38 85 39
rect 73 34 74 38
rect 78 37 85 38
rect 89 38 95 39
rect 78 34 79 37
rect 73 33 79 34
rect 89 34 90 38
rect 94 34 95 38
rect 89 33 95 34
rect 99 37 111 39
rect 99 33 100 37
rect 104 33 105 37
rect 116 33 118 42
rect 123 39 125 42
rect 123 38 134 39
rect 123 34 129 38
rect 133 34 134 38
rect 123 33 134 34
rect 9 30 11 33
rect 19 30 21 33
rect 29 29 33 33
rect 51 30 53 33
rect 29 27 43 29
rect 29 24 31 27
rect 41 24 43 27
rect 9 7 11 12
rect 19 7 21 12
rect 29 7 31 12
rect 67 28 69 33
rect 89 28 91 33
rect 67 26 91 28
rect 67 23 69 26
rect 77 23 79 26
rect 89 23 91 26
rect 99 32 105 33
rect 113 32 119 33
rect 99 23 101 32
rect 113 28 114 32
rect 118 28 119 32
rect 113 27 119 28
rect 125 23 127 33
rect 41 6 43 10
rect 51 6 53 10
rect 67 8 69 13
rect 77 8 79 13
rect 125 12 127 17
rect 89 6 91 11
rect 99 6 101 11
<< ndiffusion >>
rect 4 23 9 30
rect 2 22 9 23
rect 2 18 3 22
rect 7 18 9 22
rect 2 17 9 18
rect 4 12 9 17
rect 11 29 19 30
rect 11 25 13 29
rect 17 25 19 29
rect 11 12 19 25
rect 21 24 26 30
rect 46 24 51 30
rect 21 22 29 24
rect 21 18 23 22
rect 27 18 29 22
rect 21 12 29 18
rect 31 15 41 24
rect 31 12 34 15
rect 33 11 34 12
rect 38 11 41 15
rect 33 10 41 11
rect 43 22 51 24
rect 43 18 45 22
rect 49 18 51 22
rect 43 10 51 18
rect 53 23 65 30
rect 53 15 67 23
rect 53 11 58 15
rect 62 13 67 15
rect 69 22 77 23
rect 69 18 71 22
rect 75 18 77 22
rect 69 13 77 18
rect 79 13 89 23
rect 62 11 65 13
rect 53 10 65 11
rect 81 12 89 13
rect 81 8 82 12
rect 86 11 89 12
rect 91 22 99 23
rect 91 18 93 22
rect 97 18 99 22
rect 91 11 99 18
rect 101 12 109 23
rect 118 22 125 23
rect 118 18 119 22
rect 123 18 125 22
rect 118 17 125 18
rect 127 22 134 23
rect 127 18 129 22
rect 133 18 134 22
rect 127 17 134 18
rect 101 11 104 12
rect 86 8 87 11
rect 81 7 87 8
rect 103 8 104 11
rect 108 8 109 12
rect 103 7 109 8
<< pdiffusion >>
rect 23 69 31 70
rect 23 65 24 69
rect 28 65 31 69
rect 23 63 31 65
rect 14 61 19 63
rect 2 60 9 61
rect 2 56 3 60
rect 7 56 9 60
rect 2 42 9 56
rect 11 60 19 61
rect 11 56 13 60
rect 17 56 19 60
rect 11 53 19 56
rect 11 49 13 53
rect 17 49 19 53
rect 11 42 19 49
rect 21 42 31 63
rect 33 42 39 70
rect 41 42 47 70
rect 49 62 57 70
rect 49 58 51 62
rect 55 58 57 62
rect 49 42 57 58
rect 59 42 65 70
rect 67 42 73 70
rect 75 69 83 70
rect 75 65 77 69
rect 81 65 83 69
rect 75 42 83 65
rect 85 42 91 70
rect 93 42 99 70
rect 101 62 109 70
rect 101 58 103 62
rect 107 58 109 62
rect 101 42 109 58
rect 111 42 116 70
rect 118 42 123 70
rect 125 69 134 70
rect 125 65 129 69
rect 133 65 134 69
rect 125 62 134 65
rect 125 58 129 62
rect 133 58 134 62
rect 125 42 134 58
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect 118 78 122 82
rect 126 78 130 82
rect 134 78 138 82
rect -2 69 138 78
rect -2 68 24 69
rect 2 60 8 68
rect 23 65 24 68
rect 28 68 77 69
rect 28 65 29 68
rect 76 65 77 68
rect 81 68 129 69
rect 81 65 82 68
rect 128 65 129 68
rect 133 68 138 69
rect 133 65 134 68
rect 128 62 134 65
rect 2 56 3 60
rect 7 56 8 60
rect 13 60 51 62
rect 17 58 51 60
rect 55 58 103 62
rect 107 58 108 62
rect 128 58 129 62
rect 133 58 134 62
rect 17 56 18 58
rect 13 53 18 56
rect 2 49 13 53
rect 17 49 18 53
rect 25 50 134 54
rect 2 29 6 49
rect 17 39 23 46
rect 10 38 23 39
rect 10 34 13 38
rect 17 34 23 38
rect 10 33 23 34
rect 27 38 31 50
rect 41 42 69 46
rect 41 39 45 42
rect 27 33 31 34
rect 34 38 45 39
rect 63 38 69 42
rect 2 25 13 29
rect 17 25 18 29
rect 34 25 38 38
rect 42 34 45 38
rect 49 34 50 38
rect 54 34 55 38
rect 63 34 64 38
rect 68 34 69 38
rect 73 38 79 50
rect 73 34 74 38
rect 78 34 79 38
rect 89 42 119 46
rect 89 38 95 42
rect 89 34 90 38
rect 94 34 95 38
rect 100 37 106 38
rect 49 30 55 34
rect 104 33 106 37
rect 100 30 106 33
rect 49 26 106 30
rect 113 32 119 42
rect 129 38 134 50
rect 133 34 134 38
rect 129 33 134 34
rect 113 28 114 32
rect 118 28 119 32
rect 113 26 119 28
rect 129 22 133 23
rect 2 18 3 22
rect 7 18 23 22
rect 27 18 45 22
rect 49 18 71 22
rect 75 18 93 22
rect 97 18 119 22
rect 123 18 124 22
rect 33 12 34 15
rect -2 11 34 12
rect 38 12 39 15
rect 57 12 58 15
rect 38 11 58 12
rect 62 12 63 15
rect 129 12 133 18
rect 62 11 82 12
rect -2 8 82 11
rect 86 8 104 12
rect 108 8 138 12
rect -2 2 138 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 122 2
rect 126 -2 130 2
rect 134 -2 138 2
<< ntransistor >>
rect 9 12 11 30
rect 19 12 21 30
rect 29 12 31 24
rect 41 10 43 24
rect 51 10 53 30
rect 67 13 69 23
rect 77 13 79 23
rect 89 11 91 23
rect 99 11 101 23
rect 125 17 127 23
<< ptransistor >>
rect 9 42 11 61
rect 19 42 21 63
rect 31 42 33 70
rect 39 42 41 70
rect 47 42 49 70
rect 57 42 59 70
rect 65 42 67 70
rect 73 42 75 70
rect 83 42 85 70
rect 91 42 93 70
rect 99 42 101 70
rect 109 42 111 70
rect 116 42 118 70
rect 123 42 125 70
<< polycontact >>
rect 13 34 17 38
rect 27 34 31 38
rect 38 34 42 38
rect 50 34 54 38
rect 64 34 68 38
rect 74 34 78 38
rect 90 34 94 38
rect 100 33 104 37
rect 129 34 133 38
rect 114 28 118 32
<< ndcontact >>
rect 3 18 7 22
rect 13 25 17 29
rect 23 18 27 22
rect 34 11 38 15
rect 45 18 49 22
rect 58 11 62 15
rect 71 18 75 22
rect 82 8 86 12
rect 93 18 97 22
rect 119 18 123 22
rect 129 18 133 22
rect 104 8 108 12
<< pdcontact >>
rect 24 65 28 69
rect 3 56 7 60
rect 13 56 17 60
rect 13 49 17 53
rect 51 58 55 62
rect 77 65 81 69
rect 103 58 107 62
rect 129 65 133 69
rect 129 58 133 62
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
rect 90 -2 94 2
rect 98 -2 102 2
rect 106 -2 110 2
rect 114 -2 118 2
rect 122 -2 126 2
rect 130 -2 134 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
rect 90 78 94 82
rect 98 78 102 82
rect 106 78 110 82
rect 114 78 118 82
rect 122 78 126 82
rect 130 78 134 82
<< psubstratepdiff >>
rect 0 2 136 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 122 2
rect 126 -2 130 2
rect 134 -2 136 2
rect 0 -3 136 -2
<< nsubstratendiff >>
rect 0 82 136 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect 118 78 122 82
rect 126 78 130 82
rect 134 78 136 82
rect 0 77 136 78
<< labels >>
rlabel metal1 12 36 12 36 6 b
rlabel metal1 4 36 4 36 6 z
rlabel metal1 36 32 36 32 6 a2
rlabel metal1 20 40 20 40 6 b
rlabel metal1 28 52 28 52 6 a1
rlabel metal1 36 52 36 52 6 a1
rlabel metal1 20 60 20 60 6 z
rlabel metal1 36 60 36 60 6 z
rlabel metal1 28 60 28 60 6 z
rlabel metal1 60 28 60 28 6 a3
rlabel metal1 52 32 52 32 6 a3
rlabel metal1 52 44 52 44 6 a2
rlabel metal1 60 44 60 44 6 a2
rlabel metal1 44 44 44 44 6 a2
rlabel metal1 44 52 44 52 6 a1
rlabel metal1 52 52 52 52 6 a1
rlabel metal1 60 52 60 52 6 a1
rlabel metal1 44 60 44 60 6 z
rlabel metal1 60 60 60 60 6 z
rlabel pdcontact 52 60 52 60 6 z
rlabel metal1 68 6 68 6 6 vss
rlabel metal1 76 28 76 28 6 a3
rlabel metal1 84 28 84 28 6 a3
rlabel metal1 68 28 68 28 6 a3
rlabel metal1 76 44 76 44 6 a1
rlabel metal1 68 52 68 52 6 a1
rlabel metal1 84 52 84 52 6 a1
rlabel metal1 68 60 68 60 6 z
rlabel metal1 84 60 84 60 6 z
rlabel metal1 76 60 76 60 6 z
rlabel metal1 68 74 68 74 6 vdd
rlabel metal1 100 28 100 28 6 a3
rlabel metal1 92 28 92 28 6 a3
rlabel metal1 108 44 108 44 6 a2
rlabel metal1 100 44 100 44 6 a2
rlabel metal1 92 40 92 40 6 a2
rlabel metal1 92 52 92 52 6 a1
rlabel metal1 108 52 108 52 6 a1
rlabel metal1 100 52 100 52 6 a1
rlabel metal1 92 60 92 60 6 z
rlabel metal1 100 60 100 60 6 z
rlabel metal1 63 20 63 20 6 n3
rlabel metal1 116 36 116 36 6 a2
rlabel metal1 132 40 132 40 6 a1
rlabel metal1 116 52 116 52 6 a1
rlabel metal1 124 52 124 52 6 a1
<< end >>
