magic
tech scmos
timestamp 1179386072
<< checkpaint >>
rect -22 -25 78 105
<< ab >>
rect 0 0 56 80
<< pwell >>
rect -4 -7 60 36
<< nwell >>
rect -4 36 60 87
<< polysilicon >>
rect 10 70 12 74
rect 18 70 20 74
rect 28 70 30 74
rect 36 70 38 74
rect 48 63 54 64
rect 48 60 49 63
rect 45 59 49 60
rect 53 59 54 63
rect 45 58 54 59
rect 45 55 47 58
rect 10 42 12 45
rect 18 42 20 45
rect 28 42 30 45
rect 36 42 38 45
rect 45 43 47 46
rect 9 39 12 42
rect 16 41 22 42
rect 9 31 11 39
rect 16 37 17 41
rect 21 37 22 41
rect 16 36 22 37
rect 26 41 32 42
rect 26 37 27 41
rect 31 37 32 41
rect 36 40 40 42
rect 45 41 50 43
rect 26 36 32 37
rect 38 37 40 40
rect 38 36 44 37
rect 26 32 28 36
rect 38 32 39 36
rect 43 32 44 36
rect 2 30 11 31
rect 2 26 3 30
rect 7 26 11 30
rect 2 25 11 26
rect 9 22 11 25
rect 16 30 28 32
rect 35 31 44 32
rect 35 30 41 31
rect 16 22 18 30
rect 35 27 37 30
rect 48 27 50 41
rect 26 22 28 26
rect 45 25 50 27
rect 45 22 47 25
rect 35 12 37 16
rect 9 6 11 10
rect 16 6 18 10
rect 26 8 28 11
rect 45 8 47 16
rect 26 6 47 8
<< ndiffusion >>
rect 30 22 35 27
rect 2 15 9 22
rect 2 11 3 15
rect 7 11 9 15
rect 2 10 9 11
rect 11 10 16 22
rect 18 21 26 22
rect 18 17 20 21
rect 24 17 26 21
rect 18 11 26 17
rect 28 16 35 22
rect 37 22 42 27
rect 37 21 45 22
rect 37 17 39 21
rect 43 17 45 21
rect 37 16 45 17
rect 47 21 54 22
rect 47 17 49 21
rect 53 17 54 21
rect 47 16 54 17
rect 28 11 33 16
rect 18 10 23 11
<< pdiffusion >>
rect 2 69 10 70
rect 2 65 3 69
rect 7 65 10 69
rect 2 62 10 65
rect 2 58 3 62
rect 7 58 10 62
rect 2 45 10 58
rect 12 45 18 70
rect 20 62 28 70
rect 20 58 22 62
rect 26 58 28 62
rect 20 45 28 58
rect 30 45 36 70
rect 38 69 45 70
rect 38 65 40 69
rect 44 65 45 69
rect 38 63 45 65
rect 38 55 43 63
rect 38 46 45 55
rect 47 54 54 55
rect 47 50 49 54
rect 53 50 54 54
rect 47 49 54 50
rect 47 46 52 49
rect 38 45 43 46
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect -2 69 58 78
rect -2 68 3 69
rect 7 68 40 69
rect 39 65 40 68
rect 44 68 58 69
rect 44 65 45 68
rect 3 62 7 65
rect 3 57 7 58
rect 10 62 27 63
rect 48 62 49 63
rect 10 58 22 62
rect 26 58 27 62
rect 32 59 49 62
rect 53 59 54 63
rect 32 58 54 59
rect 10 32 14 58
rect 32 54 36 58
rect 18 50 36 54
rect 42 50 49 54
rect 53 50 54 54
rect 18 42 22 50
rect 42 46 46 50
rect 17 41 22 42
rect 30 42 46 46
rect 30 41 34 42
rect 21 37 22 41
rect 26 37 27 41
rect 31 37 34 41
rect 50 38 54 47
rect 17 36 22 37
rect 2 30 7 31
rect 2 26 3 30
rect 10 28 23 32
rect 2 22 7 26
rect 2 18 15 22
rect 19 21 23 28
rect 30 28 34 37
rect 38 36 54 38
rect 38 32 39 36
rect 43 32 54 36
rect 30 24 54 28
rect 48 21 54 24
rect 19 17 20 21
rect 24 17 25 21
rect 38 17 39 21
rect 43 17 44 21
rect 48 17 49 21
rect 53 17 54 21
rect 2 12 3 15
rect -2 11 3 12
rect 7 12 8 15
rect 38 12 44 17
rect 7 11 58 12
rect -2 2 58 11
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
<< ntransistor >>
rect 9 10 11 22
rect 16 10 18 22
rect 26 11 28 22
rect 35 16 37 27
rect 45 16 47 22
<< ptransistor >>
rect 10 45 12 70
rect 18 45 20 70
rect 28 45 30 70
rect 36 45 38 70
rect 45 46 47 55
<< polycontact >>
rect 49 59 53 63
rect 17 37 21 41
rect 27 37 31 41
rect 39 32 43 36
rect 3 26 7 30
<< ndcontact >>
rect 3 11 7 15
rect 20 17 24 21
rect 39 17 43 21
rect 49 17 53 21
<< pdcontact >>
rect 3 65 7 69
rect 3 58 7 62
rect 22 58 26 62
rect 40 65 44 69
rect 49 50 53 54
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
<< psubstratepdiff >>
rect 0 2 56 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 56 2
rect 0 -3 56 -2
<< nsubstratendiff >>
rect 0 82 56 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 56 82
rect 0 77 56 78
<< labels >>
rlabel ptransistor 29 55 29 55 6 sn
rlabel polycontact 4 28 4 28 6 a0
rlabel metal1 12 20 12 20 6 a0
rlabel metal1 12 48 12 48 6 z
rlabel metal1 28 6 28 6 6 vss
rlabel metal1 32 35 32 35 6 sn
rlabel metal1 20 44 20 44 6 s
rlabel metal1 28 52 28 52 6 s
rlabel metal1 20 60 20 60 6 z
rlabel metal1 28 74 28 74 6 vdd
rlabel metal1 44 36 44 36 6 a1
rlabel metal1 36 60 36 60 6 s
rlabel metal1 44 60 44 60 6 s
rlabel metal1 51 22 51 22 6 sn
rlabel metal1 52 40 52 40 6 a1
rlabel metal1 48 52 48 52 6 sn
<< end >>
