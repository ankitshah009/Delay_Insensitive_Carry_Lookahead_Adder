magic
tech scmos
timestamp 1183911760
<< checkpaint >>
rect -22 -25 166 105
<< ab >>
rect 0 0 144 80
<< pwell >>
rect -4 -7 148 36
<< nwell >>
rect -4 36 148 87
<< polysilicon >>
rect 9 70 11 74
rect 55 72 111 74
rect 55 64 57 72
rect 65 64 67 68
rect 75 64 77 68
rect 82 64 84 72
rect 92 64 94 68
rect 99 64 101 68
rect 19 56 21 61
rect 38 58 40 63
rect 45 58 47 63
rect 9 38 11 42
rect 19 39 21 42
rect 19 38 34 39
rect 9 37 15 38
rect 19 37 29 38
rect 9 33 10 37
rect 14 33 15 37
rect 9 32 15 33
rect 27 34 29 37
rect 33 34 34 38
rect 27 33 34 34
rect 9 28 11 32
rect 27 30 29 33
rect 38 23 40 52
rect 45 48 47 52
rect 45 47 51 48
rect 45 43 46 47
rect 50 43 51 47
rect 45 42 51 43
rect 55 38 57 52
rect 45 36 57 38
rect 45 23 47 36
rect 65 33 67 52
rect 75 48 77 58
rect 71 47 77 48
rect 71 43 72 47
rect 76 43 77 47
rect 71 42 77 43
rect 65 32 71 33
rect 51 31 57 32
rect 51 27 52 31
rect 56 27 57 31
rect 51 26 57 27
rect 55 23 57 26
rect 65 28 66 32
rect 70 28 71 32
rect 65 27 71 28
rect 65 23 67 27
rect 75 23 77 42
rect 82 38 84 58
rect 109 62 111 72
rect 129 63 131 68
rect 92 48 94 51
rect 88 47 94 48
rect 88 43 89 47
rect 93 43 94 47
rect 88 42 94 43
rect 99 39 101 51
rect 109 48 111 51
rect 129 49 131 53
rect 122 48 131 49
rect 109 46 117 48
rect 115 39 117 46
rect 122 44 123 48
rect 127 44 131 48
rect 122 43 131 44
rect 99 38 105 39
rect 82 36 94 38
rect 82 31 88 32
rect 82 27 83 31
rect 87 27 88 31
rect 82 26 88 27
rect 82 23 84 26
rect 92 23 94 36
rect 99 34 100 38
rect 104 34 105 38
rect 99 33 105 34
rect 115 38 121 39
rect 115 34 116 38
rect 120 34 121 38
rect 115 33 121 34
rect 99 23 101 33
rect 119 30 121 33
rect 129 30 131 43
rect 27 18 29 23
rect 119 19 121 24
rect 129 18 131 23
rect 9 11 11 14
rect 38 11 40 17
rect 45 12 47 17
rect 9 9 40 11
rect 55 8 57 17
rect 65 12 67 17
rect 75 12 77 17
rect 82 8 84 17
rect 92 12 94 17
rect 99 12 101 17
rect 55 6 84 8
<< ndiffusion >>
rect 20 29 27 30
rect 2 27 9 28
rect 2 23 3 27
rect 7 23 9 27
rect 2 22 9 23
rect 4 14 9 22
rect 11 20 16 28
rect 20 25 21 29
rect 25 25 27 29
rect 20 24 27 25
rect 22 23 27 24
rect 29 23 36 30
rect 112 29 119 30
rect 112 25 113 29
rect 117 25 119 29
rect 112 24 119 25
rect 121 29 129 30
rect 121 25 123 29
rect 127 25 129 29
rect 121 24 129 25
rect 11 19 18 20
rect 11 15 13 19
rect 17 15 18 19
rect 31 22 38 23
rect 31 18 32 22
rect 36 18 38 22
rect 31 17 38 18
rect 40 17 45 23
rect 47 22 55 23
rect 47 18 49 22
rect 53 18 55 22
rect 47 17 55 18
rect 57 22 65 23
rect 57 18 59 22
rect 63 18 65 22
rect 57 17 65 18
rect 67 22 75 23
rect 67 18 69 22
rect 73 18 75 22
rect 67 17 75 18
rect 77 17 82 23
rect 84 22 92 23
rect 84 18 86 22
rect 90 18 92 22
rect 84 17 92 18
rect 94 17 99 23
rect 101 22 108 23
rect 101 18 103 22
rect 107 18 108 22
rect 123 23 129 24
rect 131 29 138 30
rect 131 25 133 29
rect 137 25 138 29
rect 131 23 138 25
rect 101 17 108 18
rect 11 14 18 15
<< pdiffusion >>
rect 4 56 9 70
rect 2 54 9 56
rect 2 50 3 54
rect 7 50 9 54
rect 2 47 9 50
rect 2 43 3 47
rect 7 43 9 47
rect 2 42 9 43
rect 11 69 18 70
rect 11 65 13 69
rect 17 65 18 69
rect 11 64 18 65
rect 11 56 17 64
rect 50 58 55 64
rect 30 57 38 58
rect 11 55 19 56
rect 11 51 13 55
rect 17 51 19 55
rect 11 42 19 51
rect 21 48 26 56
rect 30 53 31 57
rect 35 53 38 57
rect 30 52 38 53
rect 40 52 45 58
rect 47 57 55 58
rect 47 53 49 57
rect 53 53 55 57
rect 47 52 55 53
rect 57 57 65 64
rect 57 53 59 57
rect 63 53 65 57
rect 57 52 65 53
rect 67 63 75 64
rect 67 59 69 63
rect 73 59 75 63
rect 67 58 75 59
rect 77 58 82 64
rect 84 63 92 64
rect 84 59 86 63
rect 90 59 92 63
rect 84 58 92 59
rect 67 52 73 58
rect 21 47 28 48
rect 21 43 23 47
rect 27 43 28 47
rect 21 42 28 43
rect 87 51 92 58
rect 94 51 99 64
rect 101 62 106 64
rect 122 62 129 63
rect 101 61 109 62
rect 101 57 103 61
rect 107 57 109 61
rect 101 51 109 57
rect 111 57 116 62
rect 122 58 123 62
rect 127 58 129 62
rect 111 56 118 57
rect 111 52 113 56
rect 117 52 118 56
rect 122 53 129 58
rect 131 59 136 63
rect 131 58 138 59
rect 131 54 133 58
rect 137 54 138 58
rect 131 53 138 54
rect 111 51 118 52
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect 118 78 122 82
rect 126 78 130 82
rect 134 78 138 82
rect 142 78 146 82
rect -2 69 146 78
rect -2 68 13 69
rect 17 68 146 69
rect 13 55 17 65
rect 2 54 7 55
rect 2 50 3 54
rect 31 57 35 68
rect 69 63 73 68
rect 69 58 73 59
rect 81 59 86 63
rect 90 59 91 63
rect 102 61 108 68
rect 59 57 63 58
rect 31 52 35 53
rect 38 53 49 57
rect 53 53 54 57
rect 13 50 17 51
rect 2 47 7 50
rect 2 43 3 47
rect 7 43 15 46
rect 2 42 15 43
rect 21 43 23 47
rect 27 43 28 47
rect 2 28 6 42
rect 21 37 25 43
rect 38 38 42 53
rect 59 47 63 53
rect 45 43 46 47
rect 9 33 10 37
rect 14 33 25 37
rect 28 34 29 38
rect 33 34 44 38
rect 21 29 25 33
rect 2 27 7 28
rect 2 23 3 27
rect 21 24 25 25
rect 2 22 7 23
rect 32 22 36 23
rect 13 19 17 20
rect 13 12 17 15
rect 40 22 44 34
rect 50 32 54 47
rect 59 43 72 47
rect 76 43 77 47
rect 50 31 56 32
rect 50 27 52 31
rect 50 26 56 27
rect 59 22 63 43
rect 81 40 85 59
rect 102 57 103 61
rect 107 57 108 61
rect 122 62 128 68
rect 122 58 123 62
rect 127 58 128 62
rect 133 58 137 59
rect 113 56 117 57
rect 76 36 85 40
rect 89 52 113 54
rect 89 50 117 52
rect 89 47 93 50
rect 121 48 127 54
rect 121 46 123 48
rect 76 33 80 36
rect 66 32 80 33
rect 89 32 93 43
rect 97 38 103 46
rect 113 44 123 46
rect 113 42 127 44
rect 133 38 137 54
rect 97 34 100 38
rect 104 34 111 38
rect 115 34 116 38
rect 120 34 137 38
rect 70 28 80 32
rect 66 27 80 28
rect 40 18 49 22
rect 53 18 54 22
rect 32 12 36 18
rect 59 17 63 18
rect 69 22 73 23
rect 76 22 80 27
rect 83 31 93 32
rect 87 30 93 31
rect 87 29 118 30
rect 87 27 113 29
rect 83 26 113 27
rect 112 25 113 26
rect 117 25 118 29
rect 123 29 127 30
rect 76 18 86 22
rect 90 18 91 22
rect 102 18 103 22
rect 107 18 108 22
rect 69 12 73 18
rect 102 12 108 18
rect 123 12 127 25
rect 133 29 137 34
rect 133 24 137 25
rect -2 2 146 12
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 122 2
rect 126 -2 130 2
rect 134 -2 138 2
rect 142 -2 146 2
<< ntransistor >>
rect 9 14 11 28
rect 27 23 29 30
rect 119 24 121 30
rect 38 17 40 23
rect 45 17 47 23
rect 55 17 57 23
rect 65 17 67 23
rect 75 17 77 23
rect 82 17 84 23
rect 92 17 94 23
rect 99 17 101 23
rect 129 23 131 30
<< ptransistor >>
rect 9 42 11 70
rect 19 42 21 56
rect 38 52 40 58
rect 45 52 47 58
rect 55 52 57 64
rect 65 52 67 64
rect 75 58 77 64
rect 82 58 84 64
rect 92 51 94 64
rect 99 51 101 64
rect 109 51 111 62
rect 129 53 131 63
<< polycontact >>
rect 10 33 14 37
rect 29 34 33 38
rect 46 43 50 47
rect 72 43 76 47
rect 52 27 56 31
rect 66 28 70 32
rect 89 43 93 47
rect 123 44 127 48
rect 83 27 87 31
rect 100 34 104 38
rect 116 34 120 38
<< ndcontact >>
rect 3 23 7 27
rect 21 25 25 29
rect 113 25 117 29
rect 123 25 127 29
rect 13 15 17 19
rect 32 18 36 22
rect 49 18 53 22
rect 59 18 63 22
rect 69 18 73 22
rect 86 18 90 22
rect 103 18 107 22
rect 133 25 137 29
<< pdcontact >>
rect 3 50 7 54
rect 3 43 7 47
rect 13 65 17 69
rect 13 51 17 55
rect 31 53 35 57
rect 49 53 53 57
rect 59 53 63 57
rect 69 59 73 63
rect 86 59 90 63
rect 23 43 27 47
rect 103 57 107 61
rect 123 58 127 62
rect 113 52 117 56
rect 133 54 137 58
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
rect 90 -2 94 2
rect 98 -2 102 2
rect 106 -2 110 2
rect 114 -2 118 2
rect 122 -2 126 2
rect 130 -2 134 2
rect 138 -2 142 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
rect 90 78 94 82
rect 98 78 102 82
rect 106 78 110 82
rect 114 78 118 82
rect 122 78 126 82
rect 130 78 134 82
rect 138 78 142 82
<< psubstratepdiff >>
rect 0 2 144 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 122 2
rect 126 -2 130 2
rect 134 -2 138 2
rect 142 -2 144 2
rect 0 -3 144 -2
<< nsubstratendiff >>
rect 0 82 144 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect 118 78 122 82
rect 126 78 130 82
rect 134 78 138 82
rect 142 78 144 82
rect 0 77 144 78
<< labels >>
rlabel polycontact 12 35 12 35 6 zn
rlabel polycontact 30 36 30 36 6 n4
rlabel polycontact 54 29 54 29 6 ci
rlabel polycontact 48 45 48 45 6 ci
rlabel polycontact 68 30 68 30 6 n1
rlabel polycontact 85 29 85 29 6 ci
rlabel polycontact 91 45 91 45 6 ci
rlabel polycontact 74 45 74 45 6 n2
rlabel polycontact 118 36 118 36 6 cn
rlabel metal1 23 35 23 35 6 zn
rlabel metal1 17 35 17 35 6 zn
rlabel metal1 4 40 4 40 6 z
rlabel metal1 12 44 12 44 6 z
rlabel metal1 47 20 47 20 6 n4
rlabel polycontact 53 29 53 29 6 ci
rlabel metal1 36 36 36 36 6 n4
rlabel pdcontact 24 45 24 45 6 zn
rlabel polycontact 49 45 49 45 6 ci
rlabel metal1 46 55 46 55 6 n4
rlabel metal1 72 6 72 6 6 vss
rlabel metal1 73 30 73 30 6 n1
rlabel metal1 68 45 68 45 6 n2
rlabel metal1 61 37 61 37 6 n2
rlabel metal1 72 74 72 74 6 vdd
rlabel metal1 83 20 83 20 6 n1
rlabel metal1 108 36 108 36 6 d
rlabel metal1 100 40 100 40 6 d
rlabel metal1 91 40 91 40 6 ci
rlabel metal1 86 61 86 61 6 n1
rlabel metal1 100 28 100 28 6 ci
rlabel metal1 116 44 116 44 6 cp
rlabel metal1 126 36 126 36 6 cn
rlabel metal1 124 48 124 48 6 cp
rlabel metal1 103 52 103 52 6 ci
rlabel metal1 135 41 135 41 6 cn
<< end >>
