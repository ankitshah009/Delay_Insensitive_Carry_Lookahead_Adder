magic
tech scmos
timestamp 1179386742
<< checkpaint >>
rect -22 -22 70 94
<< ab >>
rect 0 0 48 72
<< pwell >>
rect -4 -4 52 32
<< nwell >>
rect -4 32 52 76
<< polysilicon >>
rect 9 66 11 70
rect 16 66 18 70
rect 26 66 28 70
rect 33 66 35 70
rect 9 30 11 39
rect 16 36 18 39
rect 26 36 28 39
rect 16 34 28 36
rect 21 30 23 34
rect 27 30 28 34
rect 9 29 17 30
rect 9 27 12 29
rect 11 25 12 27
rect 16 25 17 29
rect 11 24 17 25
rect 21 29 28 30
rect 11 21 13 24
rect 21 21 23 29
rect 33 27 35 39
rect 33 26 39 27
rect 33 22 34 26
rect 38 22 39 26
rect 33 21 39 22
rect 11 2 13 6
rect 21 2 23 6
<< ndiffusion >>
rect 3 11 11 21
rect 3 7 5 11
rect 9 7 11 11
rect 3 6 11 7
rect 13 18 21 21
rect 13 14 15 18
rect 19 14 21 18
rect 13 6 21 14
rect 23 18 31 21
rect 23 14 25 18
rect 29 14 31 18
rect 23 11 31 14
rect 23 7 25 11
rect 29 7 31 11
rect 23 6 31 7
<< pdiffusion >>
rect 2 65 9 66
rect 2 61 3 65
rect 7 61 9 65
rect 2 58 9 61
rect 2 54 3 58
rect 7 54 9 58
rect 2 39 9 54
rect 11 39 16 66
rect 18 51 26 66
rect 18 47 20 51
rect 24 47 26 51
rect 18 44 26 47
rect 18 40 20 44
rect 24 40 26 44
rect 18 39 26 40
rect 28 39 33 66
rect 35 65 42 66
rect 35 61 37 65
rect 41 61 42 65
rect 35 58 42 61
rect 35 54 37 58
rect 41 54 42 58
rect 35 39 42 54
<< metal1 >>
rect -2 65 50 72
rect -2 64 3 65
rect 2 61 3 64
rect 7 64 37 65
rect 7 61 8 64
rect 2 58 8 61
rect 2 54 3 58
rect 7 54 8 58
rect 36 61 37 64
rect 41 64 50 65
rect 41 61 42 64
rect 36 58 42 61
rect 36 54 37 58
rect 41 54 42 58
rect 18 51 24 52
rect 18 47 20 51
rect 18 44 24 47
rect 18 42 20 44
rect 2 40 20 42
rect 2 38 24 40
rect 2 18 6 38
rect 34 34 39 43
rect 22 30 23 34
rect 27 30 39 34
rect 12 29 16 30
rect 16 25 34 26
rect 12 22 34 25
rect 38 22 39 26
rect 2 14 15 18
rect 19 14 20 18
rect 24 14 25 18
rect 29 14 30 18
rect 24 11 30 14
rect 34 13 39 22
rect 4 8 5 11
rect -2 7 5 8
rect 9 8 10 11
rect 24 8 25 11
rect 9 7 25 8
rect 29 8 30 11
rect 29 7 40 8
rect -2 4 40 7
rect 44 4 50 8
rect -2 0 50 4
<< ntransistor >>
rect 11 6 13 21
rect 21 6 23 21
<< ptransistor >>
rect 9 39 11 66
rect 16 39 18 66
rect 26 39 28 66
rect 33 39 35 66
<< polycontact >>
rect 23 30 27 34
rect 12 25 16 29
rect 34 22 38 26
<< ndcontact >>
rect 5 7 9 11
rect 15 14 19 18
rect 25 14 29 18
rect 25 7 29 11
<< pdcontact >>
rect 3 61 7 65
rect 3 54 7 58
rect 20 47 24 51
rect 20 40 24 44
rect 37 61 41 65
rect 37 54 41 58
<< psubstratepcontact >>
rect 40 4 44 8
<< psubstratepdiff >>
rect 39 8 45 18
rect 39 4 40 8
rect 44 4 45 8
rect 39 3 45 4
<< labels >>
rlabel metal1 4 28 4 28 6 z
rlabel metal1 12 16 12 16 6 z
rlabel metal1 20 24 20 24 6 a
rlabel metal1 12 40 12 40 6 z
rlabel metal1 20 44 20 44 6 z
rlabel metal1 24 4 24 4 6 vss
rlabel metal1 28 24 28 24 6 a
rlabel metal1 28 32 28 32 6 b
rlabel metal1 24 68 24 68 6 vdd
rlabel metal1 36 20 36 20 6 a
rlabel metal1 36 36 36 36 6 b
<< end >>
