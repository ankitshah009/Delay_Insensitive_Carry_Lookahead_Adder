.subckt nd2v5x2 a b vdd vss z
*   SPICE3 file   created from nd2v5x2.ext -      technology: scmos
m00 z      b      vdd    vdd p w=28u  l=2.3636u ad=112p     pd=36u      as=210p     ps=71u
m01 vdd    a      z      vdd p w=28u  l=2.3636u ad=210p     pd=71u      as=112p     ps=36u
m02 w1     b      z      vss n w=18u  l=2.3636u ad=45p      pd=23u      as=102p     ps=50u
m03 vss    a      w1     vss n w=18u  l=2.3636u ad=162p     pd=54u      as=45p      ps=23u
C0  b      vdd    0.014f
C1  vss    z      0.081f
C2  vss    b      0.036f
C3  z      b      0.142f
C4  a      vdd    0.042f
C5  vss    w1     0.003f
C6  vss    a      0.027f
C7  w1     b      0.008f
C8  z      a      0.033f
C9  vss    vdd    0.003f
C10 a      b      0.102f
C11 z      vdd    0.192f
C13 z      vss    0.012f
C14 a      vss    0.023f
C15 b      vss    0.015f
.ends
