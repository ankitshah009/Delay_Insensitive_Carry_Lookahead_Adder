.subckt nd3v0x05 a b c vdd vss z
*   SPICE3 file   created from nd3v0x05.ext -      technology: scmos
m00 vdd    c      z      vdd p w=10u  l=2.3636u ad=50p      pd=23.3333u as=47.3333p ps=23.3333u
m01 z      b      vdd    vdd p w=10u  l=2.3636u ad=47.3333p pd=23.3333u as=50p      ps=23.3333u
m02 vdd    a      z      vdd p w=10u  l=2.3636u ad=50p      pd=23.3333u as=47.3333p ps=23.3333u
m03 w1     c      z      vss n w=10u  l=2.3636u ad=25p      pd=15u      as=62p      ps=34u
m04 w2     b      w1     vss n w=10u  l=2.3636u ad=25p      pd=15u      as=25p      ps=15u
m05 vss    a      w2     vss n w=10u  l=2.3636u ad=70p      pd=34u      as=25p      ps=15u
C0  z      c      0.197f
C1  a      b      0.215f
C2  b      c      0.122f
C3  a      vdd    0.018f
C4  c      vdd    0.015f
C5  vss    a      0.062f
C6  vss    c      0.068f
C7  z      b      0.119f
C8  w1     c      0.014f
C9  a      c      0.065f
C10 z      vdd    0.167f
C11 b      vdd    0.074f
C12 vss    z      0.089f
C13 vss    b      0.026f
C14 vss    vdd    0.005f
C15 z      a      0.021f
C17 z      vss    0.026f
C18 a      vss    0.027f
C19 b      vss    0.030f
C20 c      vss    0.026f
.ends
