magic
tech scmos
timestamp 1185039079
<< checkpaint >>
rect -22 -24 82 124
<< ab >>
rect 0 0 60 100
<< pwell >>
rect -2 -4 62 49
<< nwell >>
rect -2 49 62 104
<< polysilicon >>
rect 11 95 13 98
rect 23 95 25 98
rect 47 75 49 78
rect 11 43 13 55
rect 23 53 25 55
rect 23 52 43 53
rect 23 51 38 52
rect 37 48 38 51
rect 42 48 43 52
rect 37 47 43 48
rect 7 42 13 43
rect 7 38 8 42
rect 12 38 13 42
rect 7 37 13 38
rect 17 42 23 43
rect 17 38 18 42
rect 22 41 23 42
rect 47 41 49 55
rect 22 39 49 41
rect 22 38 25 39
rect 17 37 25 38
rect 11 25 13 37
rect 23 25 25 37
rect 47 25 49 39
rect 47 12 49 15
rect 11 2 13 5
rect 23 2 25 5
<< ndiffusion >>
rect 3 12 11 25
rect 3 8 4 12
rect 8 8 11 12
rect 3 5 11 8
rect 13 5 23 25
rect 25 22 33 25
rect 25 18 28 22
rect 32 18 33 22
rect 25 5 33 18
rect 39 22 47 25
rect 39 18 40 22
rect 44 18 47 22
rect 39 15 47 18
rect 49 22 57 25
rect 49 18 52 22
rect 56 18 57 22
rect 49 15 57 18
<< pdiffusion >>
rect 3 92 11 95
rect 3 88 4 92
rect 8 88 11 92
rect 3 55 11 88
rect 13 55 23 95
rect 25 82 33 95
rect 25 78 28 82
rect 32 78 33 82
rect 25 72 33 78
rect 25 68 28 72
rect 32 68 33 72
rect 25 62 33 68
rect 25 58 28 62
rect 32 58 33 62
rect 25 55 33 58
rect 39 72 47 75
rect 39 68 40 72
rect 44 68 47 72
rect 39 62 47 68
rect 39 58 40 62
rect 44 58 47 62
rect 39 55 47 58
rect 49 72 57 75
rect 49 68 52 72
rect 56 68 57 72
rect 49 62 57 68
rect 49 58 52 62
rect 56 58 57 62
rect 49 55 57 58
<< metal1 >>
rect -2 96 62 101
rect -2 92 40 96
rect 44 92 52 96
rect 56 92 62 96
rect -2 88 4 92
rect 8 88 62 92
rect -2 87 62 88
rect 27 82 33 83
rect 7 42 13 82
rect 7 38 8 42
rect 12 38 13 42
rect 7 18 13 38
rect 17 42 23 82
rect 17 38 18 42
rect 22 38 23 42
rect 17 18 23 38
rect 27 78 28 82
rect 32 78 33 82
rect 27 72 33 78
rect 27 68 28 72
rect 32 68 33 72
rect 27 62 33 68
rect 39 72 45 73
rect 39 68 40 72
rect 44 68 45 72
rect 39 67 45 68
rect 51 72 57 87
rect 51 68 52 72
rect 56 68 57 72
rect 40 63 44 67
rect 27 58 28 62
rect 32 58 33 62
rect 27 22 33 58
rect 39 62 45 63
rect 39 58 40 62
rect 44 58 45 62
rect 39 57 45 58
rect 51 62 57 68
rect 51 58 52 62
rect 56 58 57 62
rect 51 57 57 58
rect 40 53 44 57
rect 37 52 44 53
rect 37 48 38 52
rect 42 48 44 52
rect 37 47 44 48
rect 40 23 44 47
rect 27 18 28 22
rect 32 18 33 22
rect 27 17 33 18
rect 39 22 45 23
rect 39 18 40 22
rect 44 18 45 22
rect 39 17 45 18
rect 51 22 57 23
rect 51 18 52 22
rect 56 18 57 22
rect 51 13 57 18
rect -2 12 62 13
rect -2 8 4 12
rect 8 8 62 12
rect -2 4 40 8
rect 44 4 52 8
rect 56 4 62 8
rect -2 -1 62 4
<< ntransistor >>
rect 11 5 13 25
rect 23 5 25 25
rect 47 15 49 25
<< ptransistor >>
rect 11 55 13 95
rect 23 55 25 95
rect 47 55 49 75
<< polycontact >>
rect 38 48 42 52
rect 8 38 12 42
rect 18 38 22 42
<< ndcontact >>
rect 4 8 8 12
rect 28 18 32 22
rect 40 18 44 22
rect 52 18 56 22
<< pdcontact >>
rect 4 88 8 92
rect 28 78 32 82
rect 28 68 32 72
rect 28 58 32 62
rect 40 68 44 72
rect 40 58 44 62
rect 52 68 56 72
rect 52 58 56 62
<< psubstratepcontact >>
rect 40 4 44 8
rect 52 4 56 8
<< nsubstratencontact >>
rect 40 92 44 96
rect 52 92 56 96
<< psubstratepdiff >>
rect 39 8 57 9
rect 39 4 40 8
rect 44 4 52 8
rect 56 4 57 8
rect 39 3 57 4
<< nsubstratendiff >>
rect 39 96 57 97
rect 39 92 40 96
rect 44 92 52 96
rect 56 92 57 96
rect 39 91 57 92
<< labels >>
rlabel metal1 10 50 10 50 6 i
rlabel metal1 10 50 10 50 6 i
rlabel metal1 20 50 20 50 6 cmd
rlabel metal1 20 50 20 50 6 cmd
rlabel metal1 30 6 30 6 6 vss
rlabel metal1 30 6 30 6 6 vss
rlabel metal1 30 50 30 50 6 nq
rlabel metal1 30 50 30 50 6 nq
rlabel metal1 30 94 30 94 6 vdd
rlabel metal1 30 94 30 94 6 vdd
<< end >>
