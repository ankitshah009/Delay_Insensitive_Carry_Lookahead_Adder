magic
tech scmos
timestamp 1179386736
<< checkpaint >>
rect -22 -25 54 105
<< ab >>
rect 0 0 32 80
<< pwell >>
rect -4 -7 36 36
<< nwell >>
rect -4 36 36 87
<< polysilicon >>
rect 12 70 14 74
rect 19 70 21 74
rect 12 39 14 42
rect 9 38 15 39
rect 9 34 10 38
rect 14 34 15 38
rect 9 33 15 34
rect 19 36 21 42
rect 19 35 25 36
rect 10 24 12 33
rect 19 31 20 35
rect 24 31 25 35
rect 19 30 25 31
rect 21 27 23 30
rect 10 11 12 16
rect 21 15 23 19
<< ndiffusion >>
rect 16 24 21 27
rect 2 16 10 24
rect 12 21 21 24
rect 12 17 14 21
rect 18 19 21 21
rect 23 24 30 27
rect 23 20 25 24
rect 29 20 30 24
rect 23 19 30 20
rect 18 17 19 19
rect 12 16 19 17
rect 2 12 8 16
rect 2 8 3 12
rect 7 8 8 12
rect 2 7 8 8
<< pdiffusion >>
rect 7 63 12 70
rect 5 62 12 63
rect 5 58 6 62
rect 10 58 12 62
rect 5 55 12 58
rect 5 51 6 55
rect 10 51 12 55
rect 5 50 12 51
rect 7 42 12 50
rect 14 42 19 70
rect 21 69 30 70
rect 21 65 25 69
rect 29 65 30 69
rect 21 62 30 65
rect 21 58 25 62
rect 29 58 30 62
rect 21 42 30 58
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect -2 69 34 78
rect -2 68 25 69
rect 29 68 34 69
rect 25 62 29 65
rect 5 58 6 62
rect 10 58 11 62
rect 5 55 11 58
rect 25 57 29 58
rect 2 23 6 55
rect 10 51 11 55
rect 18 43 22 47
rect 10 39 22 43
rect 10 38 14 39
rect 26 35 30 39
rect 10 33 14 34
rect 18 31 20 35
rect 24 31 30 35
rect 18 25 22 31
rect 25 24 29 25
rect 2 17 14 23
rect 18 17 19 21
rect 25 12 29 20
rect -2 8 3 12
rect 7 8 34 12
rect -2 2 34 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
<< ntransistor >>
rect 10 16 12 24
rect 21 19 23 27
<< ptransistor >>
rect 12 42 14 70
rect 19 42 21 70
<< polycontact >>
rect 10 34 14 38
rect 20 31 24 35
<< ndcontact >>
rect 14 17 18 21
rect 25 20 29 24
rect 3 8 7 12
<< pdcontact >>
rect 6 58 10 62
rect 6 51 10 55
rect 25 65 29 69
rect 25 58 29 62
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
<< psubstratepdiff >>
rect 0 2 32 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 32 2
rect 0 -3 32 -2
<< nsubstratendiff >>
rect 0 82 32 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 32 82
rect 0 77 32 78
<< labels >>
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 20 12 20 6 z
rlabel polycontact 12 36 12 36 6 b
rlabel metal1 16 6 16 6 6 vss
rlabel metal1 20 28 20 28 6 a
rlabel metal1 20 44 20 44 6 b
rlabel metal1 16 74 16 74 6 vdd
rlabel metal1 28 36 28 36 6 a
<< end >>
