magic
tech scmos
timestamp 1180600776
<< checkpaint >>
rect -22 -22 92 122
<< ab >>
rect 0 0 70 100
<< pwell >>
rect -4 -4 74 48
<< nwell >>
rect -4 48 74 104
<< polysilicon >>
rect 45 94 47 98
rect 57 94 59 98
rect 11 85 13 89
rect 19 85 21 89
rect 27 85 29 89
rect 11 33 13 56
rect 19 43 21 56
rect 27 53 29 56
rect 27 52 33 53
rect 27 48 28 52
rect 32 48 33 52
rect 27 47 33 48
rect 17 42 23 43
rect 17 38 18 42
rect 22 38 23 42
rect 17 37 23 38
rect 7 32 13 33
rect 7 28 8 32
rect 12 28 13 32
rect 7 27 13 28
rect 19 29 21 37
rect 31 29 33 47
rect 45 43 47 55
rect 57 43 59 55
rect 37 42 59 43
rect 37 38 38 42
rect 42 38 59 42
rect 37 37 59 38
rect 19 27 25 29
rect 31 27 37 29
rect 11 24 13 27
rect 23 24 25 27
rect 35 24 37 27
rect 45 25 47 37
rect 57 25 59 37
rect 11 10 13 14
rect 23 10 25 14
rect 35 11 37 15
rect 45 2 47 6
rect 57 2 59 6
<< ndiffusion >>
rect 40 24 45 25
rect 3 22 11 24
rect 3 18 4 22
rect 8 18 11 22
rect 3 14 11 18
rect 13 14 23 24
rect 25 22 35 24
rect 25 18 28 22
rect 32 18 35 22
rect 25 15 35 18
rect 37 15 45 24
rect 25 14 33 15
rect 15 12 21 14
rect 15 8 16 12
rect 20 8 21 12
rect 39 9 45 15
rect 15 7 21 8
rect 37 8 45 9
rect 37 4 38 8
rect 42 6 45 8
rect 47 22 57 25
rect 47 18 50 22
rect 54 18 57 22
rect 47 6 57 18
rect 59 22 67 25
rect 59 18 62 22
rect 66 18 67 22
rect 59 12 67 18
rect 59 8 62 12
rect 66 8 67 12
rect 59 6 67 8
rect 42 4 43 6
rect 37 3 43 4
<< pdiffusion >>
rect 31 92 45 94
rect 31 88 38 92
rect 42 88 45 92
rect 31 85 45 88
rect 3 82 11 85
rect 3 78 4 82
rect 8 78 11 82
rect 3 56 11 78
rect 13 56 19 85
rect 21 56 27 85
rect 29 56 45 85
rect 39 55 45 56
rect 47 82 57 94
rect 47 78 50 82
rect 54 78 57 82
rect 47 72 57 78
rect 47 68 50 72
rect 54 68 57 72
rect 47 62 57 68
rect 47 58 50 62
rect 54 58 57 62
rect 47 55 57 58
rect 59 92 67 94
rect 59 88 62 92
rect 66 88 67 92
rect 59 82 67 88
rect 59 78 62 82
rect 66 78 67 82
rect 59 72 67 78
rect 59 68 62 72
rect 66 68 67 72
rect 59 62 67 68
rect 59 58 62 62
rect 66 58 67 62
rect 59 55 67 58
<< metal1 >>
rect -2 96 72 100
rect -2 92 4 96
rect 8 92 20 96
rect 24 92 72 96
rect -2 88 38 92
rect 42 88 62 92
rect 66 88 72 92
rect 48 82 52 83
rect 62 82 66 88
rect 3 78 4 82
rect 8 78 42 82
rect 8 32 12 73
rect 8 27 12 28
rect 18 42 22 73
rect 18 27 22 38
rect 28 52 32 73
rect 28 27 32 48
rect 38 42 42 78
rect 38 22 42 38
rect 3 18 4 22
rect 8 18 28 22
rect 32 18 42 22
rect 48 78 50 82
rect 54 78 55 82
rect 48 72 52 78
rect 62 72 66 78
rect 48 68 50 72
rect 54 68 55 72
rect 48 62 52 68
rect 62 62 66 68
rect 48 58 50 62
rect 54 58 55 62
rect 48 22 52 58
rect 62 57 66 58
rect 62 22 66 23
rect 48 18 50 22
rect 54 18 55 22
rect 48 17 52 18
rect 62 12 66 18
rect -2 8 16 12
rect 20 8 62 12
rect 66 8 72 12
rect -2 4 38 8
rect 42 4 72 8
rect -2 0 72 4
<< ntransistor >>
rect 11 14 13 24
rect 23 14 25 24
rect 35 15 37 24
rect 45 6 47 25
rect 57 6 59 25
<< ptransistor >>
rect 11 56 13 85
rect 19 56 21 85
rect 27 56 29 85
rect 45 55 47 94
rect 57 55 59 94
<< polycontact >>
rect 28 48 32 52
rect 18 38 22 42
rect 8 28 12 32
rect 38 38 42 42
<< ndcontact >>
rect 4 18 8 22
rect 28 18 32 22
rect 16 8 20 12
rect 38 4 42 8
rect 50 18 54 22
rect 62 18 66 22
rect 62 8 66 12
<< pdcontact >>
rect 38 88 42 92
rect 4 78 8 82
rect 50 78 54 82
rect 50 68 54 72
rect 50 58 54 62
rect 62 88 66 92
rect 62 78 66 82
rect 62 68 66 72
rect 62 58 66 62
<< nsubstratencontact >>
rect 4 92 8 96
rect 20 92 24 96
<< nsubstratendiff >>
rect 3 96 25 97
rect 3 92 4 96
rect 8 92 20 96
rect 24 92 25 96
rect 3 91 25 92
<< labels >>
rlabel metal1 10 50 10 50 6 i2
rlabel polycontact 30 50 30 50 6 i0
rlabel metal1 20 50 20 50 6 i1
rlabel metal1 35 6 35 6 6 vss
rlabel metal1 50 50 50 50 6 q
rlabel metal1 35 94 35 94 6 vdd
<< end >>
