.subckt xaon21v0x1 a1 a2 b vdd vss z
*   SPICE3 file   created from xaon21v0x1.ext -      technology: scmos
m00 z      an     bn     vdd p w=28u  l=2.3636u ad=112p     pd=36u      as=132p     ps=57u
m01 an     bn     z      vdd p w=28u  l=2.3636u ad=125.831p pd=47.9036u as=112p     ps=36u
m02 vdd    a2     an     vdd p w=27u  l=2.3636u ad=193.554p pd=71.5663u as=121.337p ps=46.1928u
m03 vdd    a1     an     vdd p w=28u  l=2.3636u ad=200.723p pd=74.2169u as=125.831p ps=47.9036u
m04 bn     b      vdd    vdd p w=14u  l=2.3636u ad=66p      pd=28.5u    as=100.361p ps=37.1084u
m05 vdd    b      bn     vdd p w=14u  l=2.3636u ad=100.361p pd=37.1084u as=66p      ps=28.5u
m06 w1     an     vss    vss n w=13u  l=2.3636u ad=32.5p    pd=18u      as=123.825p ps=39u
m07 z      bn     w1     vss n w=13u  l=2.3636u ad=54.4375p pd=21.9375u as=32.5p    ps=18u
m08 an     b      z      vss n w=19u  l=2.3636u ad=78.8788p pd=31.0909u as=79.5625p ps=32.0625u
m09 w2     a2     an     vss n w=14u  l=2.3636u ad=35p      pd=19u      as=58.1212p ps=22.9091u
m10 vss    a1     w2     vss n w=14u  l=2.3636u ad=133.35p  pd=42u      as=35p      ps=19u
m11 bn     b      vss    vss n w=13u  l=2.3636u ad=77p      pd=40u      as=123.825p ps=39u
C0  a1     a2     0.233f
C1  b      an     0.015f
C2  z      bn     0.270f
C3  a1     an     0.038f
C4  z      vdd    0.043f
C5  a2     bn     0.227f
C6  a2     vdd    0.017f
C7  bn     an     0.860f
C8  vss    z      0.188f
C9  w2     a2     0.021f
C10 an     vdd    0.119f
C11 b      a1     0.054f
C12 vss    a2     0.055f
C13 z      a2     0.027f
C14 b      bn     0.185f
C15 vss    an     0.106f
C16 b      vdd    0.128f
C17 z      an     0.505f
C18 a1     bn     0.149f
C19 a1     vdd    0.017f
C20 a2     an     0.168f
C21 w1     z      0.010f
C22 vss    b      0.020f
C23 bn     vdd    0.464f
C24 b      z      0.007f
C25 vss    a1     0.178f
C26 b      a2     0.049f
C27 z      a1     0.011f
C28 vss    bn     0.066f
C29 w1     an     0.007f
C31 b      vss    0.047f
C32 z      vss    0.012f
C33 a1     vss    0.016f
C34 a2     vss    0.023f
C35 bn     vss    0.028f
C36 an     vss    0.018f
.ends
