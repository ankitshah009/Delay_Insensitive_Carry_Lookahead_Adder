magic
tech scmos
timestamp 1179386004
<< checkpaint >>
rect -22 -22 54 94
<< ab >>
rect 0 0 32 72
<< pwell >>
rect -4 -4 36 32
<< nwell >>
rect -4 32 36 76
<< polysilicon >>
rect 10 62 12 67
rect 20 54 22 59
rect 10 35 12 38
rect 20 35 22 38
rect 9 34 23 35
rect 9 30 18 34
rect 22 30 23 34
rect 9 29 23 30
rect 9 26 11 29
rect 9 6 11 11
<< ndiffusion >>
rect 2 25 9 26
rect 2 21 3 25
rect 7 21 9 25
rect 2 18 9 21
rect 2 14 3 18
rect 7 14 9 18
rect 2 13 9 14
rect 4 11 9 13
rect 11 24 19 26
rect 11 20 13 24
rect 17 20 19 24
rect 11 16 19 20
rect 11 12 13 16
rect 17 12 19 16
rect 11 11 19 12
<< pdiffusion >>
rect 2 61 10 62
rect 2 57 4 61
rect 8 57 10 61
rect 2 53 10 57
rect 2 49 4 53
rect 8 49 10 53
rect 2 38 10 49
rect 12 54 17 62
rect 12 50 20 54
rect 12 46 14 50
rect 18 46 20 50
rect 12 43 20 46
rect 12 39 14 43
rect 18 39 20 43
rect 12 38 20 39
rect 22 53 30 54
rect 22 49 24 53
rect 28 49 30 53
rect 22 38 30 49
<< metal1 >>
rect -2 68 34 72
rect -2 64 23 68
rect 27 64 34 68
rect 4 61 8 64
rect 4 53 8 57
rect 24 53 28 64
rect 4 48 8 49
rect 13 46 14 50
rect 18 46 19 50
rect 24 48 28 49
rect 13 43 19 46
rect 2 37 14 43
rect 18 39 19 43
rect 2 26 6 37
rect 26 35 30 43
rect 18 34 30 35
rect 22 30 30 34
rect 18 29 30 30
rect 2 25 7 26
rect 2 21 3 25
rect 2 18 7 21
rect 2 14 3 18
rect 2 13 7 14
rect 13 24 17 25
rect 13 16 17 20
rect 13 8 17 12
rect -2 4 24 8
rect 28 4 34 8
rect -2 0 34 4
<< ntransistor >>
rect 9 11 11 26
<< ptransistor >>
rect 10 38 12 62
rect 20 38 22 54
<< polycontact >>
rect 18 30 22 34
<< ndcontact >>
rect 3 21 7 25
rect 3 14 7 18
rect 13 20 17 24
rect 13 12 17 16
<< pdcontact >>
rect 4 57 8 61
rect 4 49 8 53
rect 14 46 18 50
rect 14 39 18 43
rect 24 49 28 53
<< psubstratepcontact >>
rect 24 4 28 8
<< nsubstratencontact >>
rect 23 64 27 68
<< psubstratepdiff >>
rect 23 8 29 24
rect 23 4 24 8
rect 28 4 29 8
rect 23 3 29 4
<< nsubstratendiff >>
rect 22 68 28 69
rect 22 64 23 68
rect 27 64 28 68
rect 22 62 28 64
<< labels >>
rlabel metal1 4 28 4 28 6 z
rlabel metal1 12 40 12 40 6 z
rlabel metal1 16 4 16 4 6 vss
rlabel polycontact 20 32 20 32 6 a
rlabel metal1 16 68 16 68 6 vdd
rlabel metal1 28 36 28 36 6 a
<< end >>
