magic
tech scmos
timestamp 1180600728
<< checkpaint >>
rect -22 -22 122 122
<< ab >>
rect 0 0 100 100
<< pwell >>
rect -4 -4 104 48
<< nwell >>
rect -4 48 104 104
<< polysilicon >>
rect 73 94 75 98
rect 85 94 87 98
rect 13 85 15 89
rect 25 85 27 89
rect 37 85 39 89
rect 61 76 63 80
rect 13 43 15 65
rect 7 42 15 43
rect 7 38 8 42
rect 12 38 15 42
rect 7 37 15 38
rect 13 25 15 37
rect 25 43 27 65
rect 37 43 39 65
rect 61 53 63 56
rect 61 52 69 53
rect 61 48 64 52
rect 68 48 69 52
rect 61 47 69 48
rect 25 42 33 43
rect 25 38 28 42
rect 32 38 33 42
rect 25 37 33 38
rect 37 42 43 43
rect 37 38 38 42
rect 42 38 43 42
rect 37 37 43 38
rect 25 25 27 37
rect 37 25 39 37
rect 61 25 63 47
rect 73 43 75 55
rect 85 43 87 55
rect 67 42 87 43
rect 67 38 68 42
rect 72 38 87 42
rect 67 37 87 38
rect 73 25 75 37
rect 85 25 87 37
rect 13 11 15 15
rect 25 11 27 15
rect 37 11 39 15
rect 61 11 63 15
rect 73 2 75 6
rect 85 2 87 6
<< ndiffusion >>
rect 5 15 13 25
rect 15 22 25 25
rect 15 18 18 22
rect 22 18 25 22
rect 15 15 25 18
rect 27 15 37 25
rect 39 15 47 25
rect 53 22 61 25
rect 53 18 54 22
rect 58 18 61 22
rect 53 15 61 18
rect 63 22 73 25
rect 63 18 66 22
rect 70 18 73 22
rect 63 15 73 18
rect 5 12 11 15
rect 5 8 6 12
rect 10 8 11 12
rect 41 12 47 15
rect 5 7 11 8
rect 41 8 42 12
rect 46 8 47 12
rect 65 12 73 15
rect 41 7 47 8
rect 65 8 66 12
rect 70 8 73 12
rect 65 6 73 8
rect 75 22 85 25
rect 75 18 78 22
rect 82 18 85 22
rect 75 6 85 18
rect 87 22 95 25
rect 87 18 90 22
rect 94 18 95 22
rect 87 12 95 18
rect 87 8 90 12
rect 94 8 95 12
rect 87 6 95 8
<< pdiffusion >>
rect 5 92 11 93
rect 5 88 6 92
rect 10 88 11 92
rect 65 92 73 94
rect 5 85 11 88
rect 65 88 66 92
rect 70 88 73 92
rect 5 65 13 85
rect 15 82 25 85
rect 15 78 18 82
rect 22 78 25 82
rect 15 65 25 78
rect 27 72 37 85
rect 27 68 30 72
rect 34 68 37 72
rect 27 65 37 68
rect 39 82 47 85
rect 39 78 42 82
rect 46 78 47 82
rect 65 82 73 88
rect 39 65 47 78
rect 65 78 66 82
rect 70 78 73 82
rect 65 76 73 78
rect 53 62 61 76
rect 53 58 54 62
rect 58 58 61 62
rect 53 56 61 58
rect 63 56 73 76
rect 68 55 73 56
rect 75 82 85 94
rect 75 78 78 82
rect 82 78 85 82
rect 75 72 85 78
rect 75 68 78 72
rect 82 68 85 72
rect 75 62 85 68
rect 75 58 78 62
rect 82 58 85 62
rect 75 55 85 58
rect 87 92 95 94
rect 87 88 90 92
rect 94 88 95 92
rect 87 82 95 88
rect 87 78 90 82
rect 94 78 95 82
rect 87 72 95 78
rect 87 68 90 72
rect 94 68 95 72
rect 87 62 95 68
rect 87 58 90 62
rect 94 58 95 62
rect 87 55 95 58
<< metal1 >>
rect -2 96 102 100
rect -2 92 18 96
rect 22 92 30 96
rect 34 92 42 96
rect 46 92 54 96
rect 58 92 102 96
rect -2 88 6 92
rect 10 88 66 92
rect 70 88 90 92
rect 94 88 102 92
rect 8 42 12 83
rect 66 82 70 88
rect 17 78 18 82
rect 22 78 42 82
rect 46 78 47 82
rect 66 77 70 78
rect 78 82 82 83
rect 78 72 82 78
rect 8 17 12 38
rect 18 68 30 72
rect 34 68 68 72
rect 18 22 22 68
rect 18 17 22 18
rect 28 42 32 63
rect 28 17 32 38
rect 38 42 42 63
rect 38 17 42 38
rect 54 62 58 63
rect 54 42 58 58
rect 64 52 68 68
rect 64 47 68 48
rect 78 62 82 68
rect 54 38 68 42
rect 72 38 73 42
rect 54 22 58 38
rect 54 17 58 18
rect 66 22 70 23
rect 66 12 70 18
rect 78 22 82 58
rect 90 82 94 88
rect 90 72 94 78
rect 90 62 94 68
rect 90 57 94 58
rect 78 17 82 18
rect 90 22 94 23
rect 90 12 94 18
rect -2 8 6 12
rect 10 8 42 12
rect 46 8 66 12
rect 70 8 90 12
rect 94 8 102 12
rect -2 4 18 8
rect 22 4 30 8
rect 34 4 102 8
rect -2 0 102 4
<< ntransistor >>
rect 13 15 15 25
rect 25 15 27 25
rect 37 15 39 25
rect 61 15 63 25
rect 73 6 75 25
rect 85 6 87 25
<< ptransistor >>
rect 13 65 15 85
rect 25 65 27 85
rect 37 65 39 85
rect 61 56 63 76
rect 73 55 75 94
rect 85 55 87 94
<< polycontact >>
rect 8 38 12 42
rect 64 48 68 52
rect 28 38 32 42
rect 38 38 42 42
rect 68 38 72 42
<< ndcontact >>
rect 18 18 22 22
rect 54 18 58 22
rect 66 18 70 22
rect 6 8 10 12
rect 42 8 46 12
rect 66 8 70 12
rect 78 18 82 22
rect 90 18 94 22
rect 90 8 94 12
<< pdcontact >>
rect 6 88 10 92
rect 66 88 70 92
rect 18 78 22 82
rect 30 68 34 72
rect 42 78 46 82
rect 66 78 70 82
rect 54 58 58 62
rect 78 78 82 82
rect 78 68 82 72
rect 78 58 82 62
rect 90 88 94 92
rect 90 78 94 82
rect 90 68 94 72
rect 90 58 94 62
<< psubstratepcontact >>
rect 18 4 22 8
rect 30 4 34 8
<< nsubstratencontact >>
rect 18 92 22 96
rect 30 92 34 96
rect 42 92 46 96
rect 54 92 58 96
<< psubstratepdiff >>
rect 17 8 35 9
rect 17 4 18 8
rect 22 4 30 8
rect 34 4 35 8
rect 17 3 35 4
<< nsubstratendiff >>
rect 17 96 59 97
rect 17 92 18 96
rect 22 92 30 96
rect 34 92 42 96
rect 46 92 54 96
rect 58 92 59 96
rect 17 91 59 92
<< labels >>
rlabel metal1 10 50 10 50 6 i2
rlabel polycontact 40 40 40 40 6 i0
rlabel polycontact 30 40 30 40 6 i1
rlabel metal1 50 6 50 6 6 vss
rlabel metal1 50 94 50 94 6 vdd
rlabel metal1 80 50 80 50 6 nq
<< end >>
