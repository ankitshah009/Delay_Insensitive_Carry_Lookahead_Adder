magic
tech scmos
timestamp 1179385395
<< checkpaint >>
rect -22 -25 78 105
<< ab >>
rect 0 0 56 80
<< pwell >>
rect -4 -7 60 36
<< nwell >>
rect -4 36 60 87
<< polysilicon >>
rect 9 58 11 63
rect 19 58 21 63
rect 30 59 32 64
rect 40 59 42 64
rect 9 33 11 50
rect 19 47 21 50
rect 19 46 25 47
rect 19 42 20 46
rect 24 42 25 46
rect 19 41 25 42
rect 9 32 15 33
rect 9 28 10 32
rect 14 28 15 32
rect 9 27 15 28
rect 12 24 14 27
rect 19 24 21 41
rect 30 33 32 50
rect 40 47 42 50
rect 39 46 47 47
rect 39 42 42 46
rect 46 42 47 46
rect 39 41 47 42
rect 25 32 34 33
rect 25 28 26 32
rect 30 28 34 32
rect 25 27 34 28
rect 32 24 34 27
rect 39 24 41 41
rect 12 12 14 17
rect 19 12 21 17
rect 32 12 34 17
rect 39 12 41 17
<< ndiffusion >>
rect 5 23 12 24
rect 5 19 6 23
rect 10 19 12 23
rect 5 17 12 19
rect 14 17 19 24
rect 21 22 32 24
rect 21 18 26 22
rect 30 18 32 22
rect 21 17 32 18
rect 34 17 39 24
rect 41 23 48 24
rect 41 19 43 23
rect 47 19 48 23
rect 41 17 48 19
<< pdiffusion >>
rect 23 58 30 59
rect 2 57 9 58
rect 2 53 3 57
rect 7 53 9 57
rect 2 50 9 53
rect 11 55 19 58
rect 11 51 13 55
rect 17 51 19 55
rect 11 50 19 51
rect 21 57 30 58
rect 21 53 24 57
rect 28 53 30 57
rect 21 50 30 53
rect 32 55 40 59
rect 32 51 34 55
rect 38 51 40 55
rect 32 50 40 51
rect 42 57 50 59
rect 42 53 45 57
rect 49 53 50 57
rect 42 50 50 53
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect -2 68 58 78
rect 3 57 7 68
rect 24 57 28 68
rect 3 52 7 53
rect 10 55 17 56
rect 10 51 13 55
rect 45 57 49 68
rect 24 52 28 53
rect 34 55 38 56
rect 10 50 17 51
rect 45 52 49 53
rect 10 47 14 50
rect 2 43 14 47
rect 34 46 38 51
rect 2 19 6 43
rect 19 42 20 46
rect 24 42 38 46
rect 41 46 54 47
rect 41 42 42 46
rect 46 42 54 46
rect 10 32 14 39
rect 26 32 30 39
rect 34 38 38 42
rect 34 34 47 38
rect 14 28 22 31
rect 10 27 22 28
rect 10 19 14 23
rect 2 17 14 19
rect 18 17 22 27
rect 30 28 38 31
rect 26 25 38 28
rect 43 23 47 34
rect 50 25 54 42
rect 25 18 26 22
rect 30 18 31 22
rect 43 18 47 19
rect 25 12 31 18
rect -2 2 58 12
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
<< ntransistor >>
rect 12 17 14 24
rect 19 17 21 24
rect 32 17 34 24
rect 39 17 41 24
<< ptransistor >>
rect 9 50 11 58
rect 19 50 21 58
rect 30 50 32 59
rect 40 50 42 59
<< polycontact >>
rect 20 42 24 46
rect 10 28 14 32
rect 42 42 46 46
rect 26 28 30 32
<< ndcontact >>
rect 6 19 10 23
rect 26 18 30 22
rect 43 19 47 23
<< pdcontact >>
rect 3 53 7 57
rect 13 51 17 55
rect 24 53 28 57
rect 34 51 38 55
rect 45 53 49 57
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
<< psubstratepdiff >>
rect 0 2 56 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 56 2
rect 0 -3 56 -2
<< nsubstratendiff >>
rect 0 82 56 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 56 82
rect 0 77 56 78
<< labels >>
rlabel polycontact 22 44 22 44 6 an
rlabel metal1 4 32 4 32 6 z
rlabel metal1 12 20 12 20 6 z
rlabel metal1 12 36 12 36 6 b
rlabel metal1 20 24 20 24 6 b
rlabel metal1 12 52 12 52 6 z
rlabel metal1 28 6 28 6 6 vss
rlabel metal1 28 32 28 32 6 a1
rlabel metal1 36 28 36 28 6 a1
rlabel metal1 28 44 28 44 6 an
rlabel metal1 28 74 28 74 6 vdd
rlabel metal1 45 28 45 28 6 an
rlabel metal1 52 36 52 36 6 a2
rlabel polycontact 44 44 44 44 6 a2
<< end >>
