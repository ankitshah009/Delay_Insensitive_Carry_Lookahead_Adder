magic
tech scmos
timestamp 1179386924
<< checkpaint >>
rect -22 -25 62 105
<< ab >>
rect 0 0 40 80
<< pwell >>
rect -4 -7 44 36
<< nwell >>
rect -4 36 44 87
<< polysilicon >>
rect 12 70 14 74
rect 19 70 21 74
rect 26 70 28 74
rect 12 39 14 42
rect 9 38 15 39
rect 9 34 10 38
rect 14 34 15 38
rect 9 33 15 34
rect 19 33 21 42
rect 26 39 28 42
rect 26 38 38 39
rect 26 37 33 38
rect 29 34 33 37
rect 37 34 38 38
rect 29 33 38 34
rect 9 29 11 33
rect 19 32 25 33
rect 19 28 20 32
rect 24 28 25 32
rect 19 27 25 28
rect 19 24 21 27
rect 29 24 31 33
rect 9 15 11 19
rect 19 9 21 14
rect 29 9 31 14
<< ndiffusion >>
rect 4 25 9 29
rect 2 24 9 25
rect 2 20 3 24
rect 7 20 9 24
rect 2 19 9 20
rect 11 24 17 29
rect 11 19 19 24
rect 13 14 19 19
rect 21 22 29 24
rect 21 18 23 22
rect 27 18 29 22
rect 21 14 29 18
rect 31 19 38 24
rect 31 15 33 19
rect 37 15 38 19
rect 31 14 38 15
rect 13 13 17 14
rect 11 12 17 13
rect 11 8 12 12
rect 16 8 17 12
rect 11 7 17 8
<< pdiffusion >>
rect 7 63 12 70
rect 5 62 12 63
rect 5 58 6 62
rect 10 58 12 62
rect 5 55 12 58
rect 5 51 6 55
rect 10 51 12 55
rect 5 50 12 51
rect 7 42 12 50
rect 14 42 19 70
rect 21 42 26 70
rect 28 69 38 70
rect 28 65 33 69
rect 37 65 38 69
rect 28 62 38 65
rect 28 58 33 62
rect 37 58 38 62
rect 28 42 38 58
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect -2 69 42 78
rect -2 68 33 69
rect 32 65 33 68
rect 37 68 42 69
rect 37 65 38 68
rect 32 62 38 65
rect 5 58 6 62
rect 10 58 11 62
rect 32 58 33 62
rect 37 58 38 62
rect 5 55 11 58
rect 2 25 6 55
rect 10 51 11 55
rect 18 47 22 55
rect 34 47 38 55
rect 10 43 22 47
rect 10 38 14 43
rect 26 41 38 47
rect 10 33 14 34
rect 18 35 22 39
rect 33 38 37 41
rect 18 32 24 35
rect 33 33 37 34
rect 18 31 20 32
rect 24 28 31 30
rect 20 26 31 28
rect 2 24 7 25
rect 2 20 3 24
rect 7 20 23 22
rect 2 18 23 20
rect 27 18 28 22
rect 33 19 37 20
rect 33 12 37 15
rect -2 8 12 12
rect 16 8 42 12
rect -2 2 42 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
<< ntransistor >>
rect 9 19 11 29
rect 19 14 21 24
rect 29 14 31 24
<< ptransistor >>
rect 12 42 14 70
rect 19 42 21 70
rect 26 42 28 70
<< polycontact >>
rect 10 34 14 38
rect 33 34 37 38
rect 20 28 24 32
<< ndcontact >>
rect 3 20 7 24
rect 23 18 27 22
rect 33 15 37 19
rect 12 8 16 12
<< pdcontact >>
rect 6 58 10 62
rect 6 51 10 55
rect 33 65 37 69
rect 33 58 37 62
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
<< psubstratepdiff >>
rect 0 2 40 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 40 2
rect 0 -3 40 -2
<< nsubstratendiff >>
rect 0 82 40 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 40 82
rect 0 77 40 78
<< labels >>
rlabel metal1 4 40 4 40 6 z
rlabel metal1 12 20 12 20 6 z
rlabel metal1 12 40 12 40 6 c
rlabel metal1 20 6 20 6 6 vss
rlabel metal1 20 6 20 6 6 vss
rlabel metal1 20 20 20 20 6 z
rlabel metal1 20 36 20 36 6 b
rlabel metal1 28 28 28 28 6 b
rlabel metal1 28 44 28 44 6 a
rlabel metal1 20 52 20 52 6 c
rlabel metal1 20 74 20 74 6 vdd
rlabel metal1 20 74 20 74 6 vdd
rlabel metal1 36 48 36 48 6 a
<< end >>
