magic
tech scmos
timestamp 1179386399
<< checkpaint >>
rect -22 -25 78 105
<< ab >>
rect 0 0 56 80
<< pwell >>
rect -4 -7 60 36
<< nwell >>
rect -4 36 60 87
<< polysilicon >>
rect 14 58 16 63
rect 24 58 26 63
rect 35 58 37 63
rect 45 58 47 63
rect 14 39 16 42
rect 24 39 26 42
rect 35 39 37 42
rect 45 39 47 42
rect 9 38 26 39
rect 9 34 10 38
rect 14 34 26 38
rect 9 33 26 34
rect 24 30 26 33
rect 31 38 47 39
rect 31 34 42 38
rect 46 34 47 38
rect 31 33 47 34
rect 31 30 33 33
rect 24 12 26 17
rect 31 12 33 17
<< ndiffusion >>
rect 17 29 24 30
rect 17 25 18 29
rect 22 25 24 29
rect 17 22 24 25
rect 17 18 18 22
rect 22 18 24 22
rect 17 17 24 18
rect 26 17 31 30
rect 33 29 41 30
rect 33 25 35 29
rect 39 25 41 29
rect 33 22 41 25
rect 33 18 35 22
rect 39 18 41 22
rect 33 17 41 18
<< pdiffusion >>
rect 6 57 14 58
rect 6 53 8 57
rect 12 53 14 57
rect 6 42 14 53
rect 16 54 24 58
rect 16 50 18 54
rect 22 50 24 54
rect 16 47 24 50
rect 16 43 18 47
rect 22 43 24 47
rect 16 42 24 43
rect 26 57 35 58
rect 26 53 28 57
rect 32 53 35 57
rect 26 42 35 53
rect 37 54 45 58
rect 37 50 39 54
rect 43 50 45 54
rect 37 47 45 50
rect 37 43 39 47
rect 43 43 45 47
rect 37 42 45 43
rect 47 57 54 58
rect 47 53 49 57
rect 53 53 54 57
rect 47 50 54 53
rect 47 46 49 50
rect 53 46 54 50
rect 47 42 54 46
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect -2 68 58 78
rect 8 57 12 68
rect 28 57 32 68
rect 8 52 12 53
rect 18 54 22 55
rect 49 57 53 68
rect 28 52 32 53
rect 39 54 43 55
rect 18 47 22 50
rect 2 39 6 47
rect 39 47 43 50
rect 22 43 39 46
rect 49 50 53 53
rect 49 45 53 46
rect 18 42 43 43
rect 2 38 14 39
rect 2 34 10 38
rect 2 33 14 34
rect 18 29 22 42
rect 41 34 42 38
rect 46 34 54 38
rect 18 22 22 25
rect 18 17 22 18
rect 35 29 39 30
rect 50 25 54 34
rect 35 22 39 25
rect 35 12 39 18
rect -2 2 58 12
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
<< ntransistor >>
rect 24 17 26 30
rect 31 17 33 30
<< ptransistor >>
rect 14 42 16 58
rect 24 42 26 58
rect 35 42 37 58
rect 45 42 47 58
<< polycontact >>
rect 10 34 14 38
rect 42 34 46 38
<< ndcontact >>
rect 18 25 22 29
rect 18 18 22 22
rect 35 25 39 29
rect 35 18 39 22
<< pdcontact >>
rect 8 53 12 57
rect 18 50 22 54
rect 18 43 22 47
rect 28 53 32 57
rect 39 50 43 54
rect 39 43 43 47
rect 49 53 53 57
rect 49 46 53 50
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
<< psubstratepdiff >>
rect 0 2 56 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 56 2
rect 0 -3 56 -2
<< nsubstratendiff >>
rect 0 82 56 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 56 82
rect 0 77 56 78
<< labels >>
rlabel metal1 4 40 4 40 6 b
rlabel polycontact 12 36 12 36 6 b
rlabel metal1 20 36 20 36 6 z
rlabel metal1 28 6 28 6 6 vss
rlabel metal1 36 44 36 44 6 z
rlabel metal1 28 44 28 44 6 z
rlabel metal1 28 74 28 74 6 vdd
rlabel polycontact 44 36 44 36 6 a
rlabel metal1 52 28 52 28 6 a
<< end >>
