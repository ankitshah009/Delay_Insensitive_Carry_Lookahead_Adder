.subckt oa22_x2 i0 i1 i2 q vdd vss
*   SPICE3 file   created from oa22_x2.ext -      technology: scmos
m00 w1     i0     w2     vdd p w=20u  l=2.3636u ad=100p     pd=30u      as=120p     ps=38.6667u
m01 w2     i1     w1     vdd p w=20u  l=2.3636u ad=120p     pd=38.6667u as=100p     ps=30u
m02 vdd    i2     w2     vdd p w=20u  l=2.3636u ad=120p     pd=33.3333u as=120p     ps=38.6667u
m03 q      w1     vdd    vdd p w=40u  l=2.3636u ad=320p     pd=96u      as=240p     ps=66.6667u
m04 w3     i0     vss    vss n w=10u  l=2.3636u ad=50p      pd=20u      as=77p      ps=28u
m05 w1     i1     w3     vss n w=10u  l=2.3636u ad=50p      pd=20u      as=50p      ps=20u
m06 vss    i2     w1     vss n w=10u  l=2.3636u ad=77p      pd=28u      as=50p      ps=20u
m07 q      w1     vss    vss n w=20u  l=2.3636u ad=160p     pd=56u      as=154p     ps=56u
C0  vss    q      0.099f
C1  i0     vdd    0.010f
C2  q      w2     0.023f
C3  w3     i1     0.016f
C4  vss    i2     0.055f
C5  w2     i2     0.050f
C6  vss    i0     0.051f
C7  q      i1     0.057f
C8  i2     i1     0.134f
C9  w2     i0     0.027f
C10 q      w1     0.139f
C11 i2     w1     0.456f
C12 i1     i0     0.400f
C13 w2     vdd    0.218f
C14 i1     vdd    0.011f
C15 i0     w1     0.111f
C16 w1     vdd    0.045f
C17 vss    i1     0.042f
C18 w3     i0     0.004f
C19 q      i2     0.485f
C20 w2     i1     0.017f
C21 q      i0     0.039f
C22 vss    w1     0.058f
C23 q      vdd    0.123f
C24 i2     i0     0.080f
C25 w2     w1     0.170f
C26 i1     w1     0.343f
C27 i2     vdd    0.088f
C29 q      vss    0.015f
C30 i2     vss    0.043f
C31 i1     vss    0.043f
C32 i0     vss    0.040f
C33 w1     vss    0.045f
.ends
