magic
tech scmos
timestamp 1180600799
<< checkpaint >>
rect -22 -22 172 122
<< ab >>
rect 0 0 150 100
<< pwell >>
rect -4 -4 154 48
<< nwell >>
rect -4 48 154 104
<< polysilicon >>
rect 11 94 13 98
rect 23 94 25 98
rect 47 94 49 98
rect 59 94 61 98
rect 71 94 73 98
rect 83 94 85 98
rect 111 94 113 98
rect 123 94 125 98
rect 135 94 137 98
rect 11 53 13 56
rect 7 52 13 53
rect 7 48 8 52
rect 12 48 13 52
rect 7 47 13 48
rect 11 25 13 47
rect 23 53 25 56
rect 47 53 49 56
rect 59 53 61 56
rect 71 53 73 56
rect 83 53 85 56
rect 111 53 113 56
rect 23 52 33 53
rect 23 48 28 52
rect 32 48 33 52
rect 23 47 33 48
rect 47 52 53 53
rect 47 48 48 52
rect 52 48 53 52
rect 47 47 53 48
rect 57 52 63 53
rect 57 48 58 52
rect 62 48 63 52
rect 57 47 63 48
rect 67 52 73 53
rect 67 48 68 52
rect 72 48 73 52
rect 67 47 73 48
rect 77 52 85 53
rect 77 48 78 52
rect 82 51 85 52
rect 107 52 113 53
rect 82 48 83 51
rect 77 47 83 48
rect 107 48 108 52
rect 112 48 113 52
rect 107 47 113 48
rect 123 53 125 56
rect 123 52 129 53
rect 123 48 124 52
rect 128 48 129 52
rect 123 47 129 48
rect 23 25 25 47
rect 51 25 53 47
rect 59 25 61 47
rect 71 25 73 47
rect 79 25 81 47
rect 93 42 99 43
rect 93 38 94 42
rect 98 41 99 42
rect 135 41 137 55
rect 98 39 137 41
rect 98 38 99 39
rect 93 37 99 38
rect 111 32 117 33
rect 111 28 112 32
rect 116 28 117 32
rect 111 27 117 28
rect 115 24 117 27
rect 123 32 129 33
rect 123 28 124 32
rect 128 28 129 32
rect 123 27 129 28
rect 123 24 125 27
rect 135 25 137 39
rect 11 2 13 6
rect 23 2 25 6
rect 51 2 53 6
rect 59 2 61 6
rect 71 2 73 6
rect 79 2 81 6
rect 115 2 117 6
rect 123 2 125 6
rect 135 2 137 6
<< ndiffusion >>
rect 3 12 11 25
rect 3 8 4 12
rect 8 8 11 12
rect 3 6 11 8
rect 13 6 23 25
rect 25 22 33 25
rect 25 18 28 22
rect 32 18 33 22
rect 25 6 33 18
rect 43 12 51 25
rect 43 8 44 12
rect 48 8 51 12
rect 43 6 51 8
rect 53 6 59 25
rect 61 22 71 25
rect 61 18 64 22
rect 68 18 71 22
rect 61 6 71 18
rect 73 6 79 25
rect 81 12 89 25
rect 130 24 135 25
rect 107 22 115 24
rect 107 18 108 22
rect 112 18 115 22
rect 81 8 84 12
rect 88 8 89 12
rect 81 6 89 8
rect 107 6 115 18
rect 117 6 123 24
rect 125 12 135 24
rect 125 8 128 12
rect 132 8 135 12
rect 125 6 135 8
rect 137 22 145 25
rect 137 18 140 22
rect 144 18 145 22
rect 137 6 145 18
<< pdiffusion >>
rect 3 82 11 94
rect 3 78 4 82
rect 8 78 11 82
rect 3 72 11 78
rect 3 68 4 72
rect 8 68 11 72
rect 3 56 11 68
rect 13 72 23 94
rect 13 68 16 72
rect 20 68 23 72
rect 13 56 23 68
rect 25 82 33 94
rect 25 78 28 82
rect 32 78 33 82
rect 25 72 33 78
rect 25 68 28 72
rect 32 68 33 72
rect 25 56 33 68
rect 39 82 47 94
rect 39 78 40 82
rect 44 78 47 82
rect 39 56 47 78
rect 49 72 59 94
rect 49 68 52 72
rect 56 68 59 72
rect 49 56 59 68
rect 61 82 71 94
rect 61 78 64 82
rect 68 78 71 82
rect 61 72 71 78
rect 61 68 64 72
rect 68 68 71 72
rect 61 56 71 68
rect 73 72 83 94
rect 73 68 76 72
rect 80 68 83 72
rect 73 56 83 68
rect 85 82 93 94
rect 85 78 88 82
rect 92 78 93 82
rect 85 56 93 78
rect 103 92 111 94
rect 103 88 104 92
rect 108 88 111 92
rect 103 82 111 88
rect 103 78 104 82
rect 108 78 111 82
rect 103 56 111 78
rect 113 82 123 94
rect 113 78 116 82
rect 120 78 123 82
rect 113 56 123 78
rect 125 92 135 94
rect 125 88 128 92
rect 132 88 135 92
rect 125 82 135 88
rect 125 78 128 82
rect 132 78 135 82
rect 125 56 135 78
rect 130 55 135 56
rect 137 82 145 94
rect 137 78 140 82
rect 144 78 145 82
rect 137 72 145 78
rect 137 68 140 72
rect 144 68 145 72
rect 137 62 145 68
rect 137 58 140 62
rect 144 58 145 62
rect 137 55 145 58
<< metal1 >>
rect -2 92 152 100
rect -2 88 104 92
rect 108 88 128 92
rect 132 88 152 92
rect 4 82 8 83
rect 28 82 32 83
rect 104 82 108 88
rect 8 78 28 82
rect 39 78 40 82
rect 44 78 64 82
rect 68 78 88 82
rect 92 78 93 82
rect 4 72 8 78
rect 28 72 32 78
rect 64 72 68 78
rect 104 77 108 78
rect 116 82 120 83
rect 116 72 120 78
rect 128 82 132 88
rect 128 77 132 78
rect 138 82 142 83
rect 138 78 140 82
rect 144 78 145 82
rect 15 68 16 72
rect 20 68 22 72
rect 4 67 8 68
rect 8 52 12 63
rect 8 17 12 48
rect 18 22 22 68
rect 32 68 52 72
rect 56 68 57 72
rect 75 68 76 72
rect 80 68 120 72
rect 28 67 32 68
rect 64 67 68 68
rect 28 52 32 63
rect 28 27 32 48
rect 48 52 52 63
rect 48 27 52 48
rect 58 52 62 63
rect 58 27 62 48
rect 68 52 72 63
rect 68 27 72 48
rect 78 52 82 63
rect 78 27 82 48
rect 108 52 112 63
rect 123 48 124 52
rect 94 42 98 43
rect 94 22 98 38
rect 108 27 112 48
rect 116 28 117 32
rect 123 28 124 32
rect 128 27 132 73
rect 138 72 142 78
rect 138 68 140 72
rect 144 68 145 72
rect 138 62 142 68
rect 138 58 140 62
rect 144 58 145 62
rect 138 22 142 58
rect 18 18 28 22
rect 32 18 64 22
rect 68 18 108 22
rect 112 18 113 22
rect 138 18 140 22
rect 144 18 145 22
rect 138 17 142 18
rect -2 8 4 12
rect 8 8 44 12
rect 48 8 84 12
rect 88 10 128 12
rect 88 8 96 10
rect -2 6 96 8
rect 100 8 128 10
rect 132 8 152 12
rect 100 6 152 8
rect -2 0 152 6
<< ntransistor >>
rect 11 6 13 25
rect 23 6 25 25
rect 51 6 53 25
rect 59 6 61 25
rect 71 6 73 25
rect 79 6 81 25
rect 115 6 117 24
rect 123 6 125 24
rect 135 6 137 25
<< ptransistor >>
rect 11 56 13 94
rect 23 56 25 94
rect 47 56 49 94
rect 59 56 61 94
rect 71 56 73 94
rect 83 56 85 94
rect 111 56 113 94
rect 123 56 125 94
rect 135 55 137 94
<< polycontact >>
rect 8 48 12 52
rect 28 48 32 52
rect 48 48 52 52
rect 58 48 62 52
rect 68 48 72 52
rect 78 48 82 52
rect 108 48 112 52
rect 124 48 128 52
rect 94 38 98 42
rect 112 28 116 32
rect 124 28 128 32
<< ndcontact >>
rect 4 8 8 12
rect 28 18 32 22
rect 44 8 48 12
rect 64 18 68 22
rect 108 18 112 22
rect 84 8 88 12
rect 128 8 132 12
rect 140 18 144 22
<< pdcontact >>
rect 4 78 8 82
rect 4 68 8 72
rect 16 68 20 72
rect 28 78 32 82
rect 28 68 32 72
rect 40 78 44 82
rect 52 68 56 72
rect 64 78 68 82
rect 64 68 68 72
rect 76 68 80 72
rect 88 78 92 82
rect 104 88 108 92
rect 104 78 108 82
rect 116 78 120 82
rect 128 88 132 92
rect 128 78 132 82
rect 140 78 144 82
rect 140 68 144 72
rect 140 58 144 62
<< psubstratepcontact >>
rect 96 6 100 10
<< psubstratepdiff >>
rect 95 10 101 16
rect 95 6 96 10
rect 100 6 101 10
rect 95 5 101 6
<< labels >>
rlabel metal1 10 40 10 40 6 i7
rlabel metal1 30 45 30 45 6 i6
rlabel metal1 50 45 50 45 6 i5
rlabel metal1 75 6 75 6 6 vss
rlabel metal1 60 45 60 45 6 i4
rlabel metal1 70 45 70 45 6 i3
rlabel metal1 80 45 80 45 6 i2
rlabel metal1 75 94 75 94 6 vdd
rlabel metal1 110 45 110 45 6 i1
rlabel metal1 140 50 140 50 6 q
rlabel metal1 130 50 130 50 6 i0
<< end >>
