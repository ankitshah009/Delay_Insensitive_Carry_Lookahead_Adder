magic
tech scmos
timestamp 1179387396
<< checkpaint >>
rect -22 -25 46 105
<< ab >>
rect 0 0 24 80
<< pwell >>
rect -4 -7 28 36
<< nwell >>
rect -4 36 28 87
<< polysilicon >>
rect 12 61 14 65
rect 12 40 14 43
rect 4 39 14 40
rect 4 35 5 39
rect 9 35 14 39
rect 4 34 14 35
rect 12 30 14 34
rect 12 6 14 10
<< ndiffusion >>
rect 3 29 12 30
rect 3 25 4 29
rect 8 25 12 29
rect 3 22 12 25
rect 3 18 4 22
rect 8 18 12 22
rect 3 10 12 18
rect 14 22 22 30
rect 14 18 17 22
rect 21 18 22 22
rect 14 15 22 18
rect 14 11 17 15
rect 21 11 22 15
rect 14 10 22 11
<< pdiffusion >>
rect 3 72 10 73
rect 3 68 5 72
rect 9 68 10 72
rect 3 64 10 68
rect 3 60 5 64
rect 9 61 10 64
rect 9 60 12 61
rect 3 56 12 60
rect 3 52 5 56
rect 9 52 12 56
rect 3 48 12 52
rect 3 44 5 48
rect 9 44 12 48
rect 3 43 12 44
rect 14 56 22 61
rect 14 52 17 56
rect 21 52 22 56
rect 14 48 22 52
rect 14 44 17 48
rect 21 44 22 48
rect 14 43 22 44
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect -2 72 26 78
rect -2 68 5 72
rect 9 68 26 72
rect 4 64 10 68
rect 4 60 5 64
rect 9 60 10 64
rect 4 56 10 60
rect 4 52 5 56
rect 9 52 10 56
rect 4 48 10 52
rect 4 44 5 48
rect 9 44 10 48
rect 4 39 10 44
rect 4 35 5 39
rect 9 35 10 39
rect 17 56 22 63
rect 21 52 22 56
rect 17 48 22 52
rect 21 44 22 48
rect 17 31 22 44
rect 2 29 22 31
rect 2 25 4 29
rect 8 25 22 29
rect 2 22 8 25
rect 2 18 4 22
rect 2 17 8 18
rect 16 18 17 22
rect 21 18 22 22
rect 16 15 22 18
rect 16 12 17 15
rect -2 11 17 12
rect 21 12 22 15
rect 21 11 26 12
rect -2 2 26 11
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
<< ntransistor >>
rect 12 10 14 30
<< ptransistor >>
rect 12 43 14 61
<< polycontact >>
rect 5 35 9 39
<< ndcontact >>
rect 4 25 8 29
rect 4 18 8 22
rect 17 18 21 22
rect 17 11 21 15
<< pdcontact >>
rect 5 68 9 72
rect 5 60 9 64
rect 5 52 9 56
rect 5 44 9 48
rect 17 52 21 56
rect 17 44 21 48
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
<< psubstratepdiff >>
rect 0 2 24 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 24 2
rect 0 -3 24 -2
<< nsubstratendiff >>
rect 0 82 24 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 24 82
rect 0 77 24 78
<< labels >>
rlabel metal1 4 24 4 24 6 z
rlabel metal1 12 6 12 6 6 vss
rlabel metal1 12 28 12 28 6 z
rlabel metal1 12 74 12 74 6 vdd
rlabel metal1 20 44 20 44 6 z
<< end >>
