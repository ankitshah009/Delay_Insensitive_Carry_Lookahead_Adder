magic
tech scmos
timestamp 1179386318
<< checkpaint >>
rect -22 -22 78 94
<< ab >>
rect 0 0 56 72
<< pwell >>
rect -4 -4 60 32
<< nwell >>
rect -4 32 60 76
<< polysilicon >>
rect 9 66 11 70
rect 19 66 21 70
rect 29 58 31 63
rect 39 58 41 63
rect 9 35 11 38
rect 19 35 21 38
rect 29 35 31 38
rect 39 35 41 38
rect 9 34 15 35
rect 9 30 10 34
rect 14 30 15 34
rect 9 29 15 30
rect 19 34 31 35
rect 19 30 26 34
rect 30 30 31 34
rect 19 29 31 30
rect 12 26 14 29
rect 19 26 21 29
rect 29 26 31 29
rect 36 34 42 35
rect 36 30 37 34
rect 41 30 42 34
rect 36 29 42 30
rect 36 26 38 29
rect 12 2 14 6
rect 19 2 21 6
rect 29 2 31 6
rect 36 2 38 6
<< ndiffusion >>
rect 3 8 12 26
rect 3 4 5 8
rect 9 6 12 8
rect 14 6 19 26
rect 21 18 29 26
rect 21 14 23 18
rect 27 14 29 18
rect 21 6 29 14
rect 31 6 36 26
rect 38 18 46 26
rect 38 14 41 18
rect 45 14 46 18
rect 38 13 46 14
rect 38 6 43 13
rect 9 4 10 6
rect 3 3 10 4
<< pdiffusion >>
rect 2 65 9 66
rect 2 61 3 65
rect 7 61 9 65
rect 2 58 9 61
rect 2 54 3 58
rect 7 54 9 58
rect 2 38 9 54
rect 11 50 19 66
rect 11 46 13 50
rect 17 46 19 50
rect 11 43 19 46
rect 11 39 13 43
rect 17 39 19 43
rect 11 38 19 39
rect 21 58 27 66
rect 21 57 29 58
rect 21 53 23 57
rect 27 53 29 57
rect 21 38 29 53
rect 31 57 39 58
rect 31 53 33 57
rect 37 53 39 57
rect 31 50 39 53
rect 31 46 33 50
rect 37 46 39 50
rect 31 38 39 46
rect 41 57 49 58
rect 41 53 43 57
rect 47 53 49 57
rect 41 50 49 53
rect 41 46 43 50
rect 47 46 49 50
rect 41 38 49 46
<< metal1 >>
rect -2 68 58 72
rect -2 65 48 68
rect -2 64 3 65
rect 2 61 3 64
rect 7 64 48 65
rect 52 64 58 68
rect 7 61 8 64
rect 2 58 8 61
rect 2 54 3 58
rect 7 54 8 58
rect 22 57 28 64
rect 22 53 23 57
rect 27 53 28 57
rect 33 57 38 59
rect 37 53 38 57
rect 33 50 38 53
rect 12 46 13 50
rect 17 46 33 50
rect 37 46 38 50
rect 42 57 48 64
rect 42 53 43 57
rect 47 53 48 57
rect 42 50 48 53
rect 42 46 43 50
rect 47 46 48 50
rect 12 43 18 46
rect 2 39 13 43
rect 17 39 18 43
rect 2 18 6 39
rect 25 38 39 42
rect 10 34 14 35
rect 25 34 31 38
rect 25 30 26 34
rect 30 30 31 34
rect 36 30 37 34
rect 41 30 42 34
rect 10 26 14 30
rect 36 26 42 30
rect 10 22 47 26
rect 2 14 23 18
rect 27 14 31 18
rect 40 14 41 18
rect 45 14 46 18
rect 40 8 46 14
rect -2 4 5 8
rect 9 4 48 8
rect 52 4 58 8
rect -2 0 58 4
<< ntransistor >>
rect 12 6 14 26
rect 19 6 21 26
rect 29 6 31 26
rect 36 6 38 26
<< ptransistor >>
rect 9 38 11 66
rect 19 38 21 66
rect 29 38 31 58
rect 39 38 41 58
<< polycontact >>
rect 10 30 14 34
rect 26 30 30 34
rect 37 30 41 34
<< ndcontact >>
rect 5 4 9 8
rect 23 14 27 18
rect 41 14 45 18
<< pdcontact >>
rect 3 61 7 65
rect 3 54 7 58
rect 13 46 17 50
rect 13 39 17 43
rect 23 53 27 57
rect 33 53 37 57
rect 33 46 37 50
rect 43 53 47 57
rect 43 46 47 50
<< psubstratepcontact >>
rect 48 4 52 8
<< nsubstratencontact >>
rect 48 64 52 68
<< psubstratepdiff >>
rect 47 8 53 9
rect 47 4 48 8
rect 52 4 53 8
rect 47 3 53 4
<< nsubstratendiff >>
rect 47 68 53 69
rect 47 64 48 68
rect 52 64 53 68
rect 47 63 53 64
<< labels >>
rlabel metal1 4 32 4 32 6 z
rlabel metal1 20 16 20 16 6 z
rlabel metal1 12 16 12 16 6 z
rlabel polycontact 12 32 12 32 6 a
rlabel metal1 20 24 20 24 6 a
rlabel metal1 20 48 20 48 6 z
rlabel metal1 28 4 28 4 6 vss
rlabel metal1 28 16 28 16 6 z
rlabel metal1 28 24 28 24 6 a
rlabel metal1 36 24 36 24 6 a
rlabel metal1 36 40 36 40 6 b
rlabel metal1 28 36 28 36 6 b
rlabel metal1 28 48 28 48 6 z
rlabel pdcontact 36 56 36 56 6 z
rlabel metal1 28 68 28 68 6 vdd
rlabel metal1 44 24 44 24 6 a
<< end >>
