magic
tech scmos
timestamp 1179385305
<< checkpaint >>
rect -22 -22 118 94
<< ab >>
rect 0 0 96 72
<< pwell >>
rect -4 -4 100 32
<< nwell >>
rect -4 32 100 76
<< polysilicon >>
rect 9 66 11 70
rect 19 66 21 70
rect 29 66 31 70
rect 39 66 41 70
rect 49 66 51 70
rect 59 66 61 70
rect 69 66 71 70
rect 81 66 83 70
rect 9 35 11 38
rect 19 35 21 38
rect 29 35 31 38
rect 39 35 41 38
rect 49 35 51 38
rect 59 35 61 38
rect 69 35 71 38
rect 9 34 15 35
rect 9 30 10 34
rect 14 30 15 34
rect 9 29 15 30
rect 19 34 31 35
rect 19 30 23 34
rect 27 30 31 34
rect 19 29 31 30
rect 12 21 14 29
rect 19 21 21 29
rect 29 26 31 29
rect 36 34 42 35
rect 36 30 37 34
rect 41 30 42 34
rect 36 29 42 30
rect 49 34 55 35
rect 49 30 50 34
rect 54 30 55 34
rect 49 29 55 30
rect 59 34 71 35
rect 59 30 65 34
rect 69 30 71 34
rect 81 35 83 38
rect 81 34 87 35
rect 81 31 82 34
rect 59 29 71 30
rect 36 26 38 29
rect 52 26 54 29
rect 59 26 61 29
rect 69 26 71 29
rect 76 30 82 31
rect 86 30 87 34
rect 76 29 87 30
rect 76 26 78 29
rect 69 11 71 16
rect 76 11 78 16
rect 12 6 14 11
rect 19 6 21 11
rect 29 6 31 11
rect 36 6 38 11
rect 52 6 54 11
rect 59 6 61 11
<< ndiffusion >>
rect 24 21 29 26
rect 4 11 12 21
rect 14 11 19 21
rect 21 17 29 21
rect 21 13 23 17
rect 27 13 29 17
rect 21 11 29 13
rect 31 11 36 26
rect 38 16 52 26
rect 38 12 43 16
rect 47 12 52 16
rect 38 11 52 12
rect 54 11 59 26
rect 61 23 69 26
rect 61 19 63 23
rect 67 19 69 23
rect 61 16 69 19
rect 71 16 76 26
rect 78 21 88 26
rect 78 17 82 21
rect 86 17 88 21
rect 78 16 88 17
rect 61 11 66 16
rect 4 8 10 11
rect 4 4 5 8
rect 9 4 10 8
rect 4 3 10 4
<< pdiffusion >>
rect 73 67 79 68
rect 73 66 74 67
rect 4 60 9 66
rect 2 59 9 60
rect 2 55 3 59
rect 7 55 9 59
rect 2 54 9 55
rect 4 38 9 54
rect 11 50 19 66
rect 11 46 13 50
rect 17 46 19 50
rect 11 38 19 46
rect 21 59 29 66
rect 21 55 23 59
rect 27 55 29 59
rect 21 38 29 55
rect 31 50 39 66
rect 31 46 33 50
rect 37 46 39 50
rect 31 38 39 46
rect 41 58 49 66
rect 41 54 43 58
rect 47 54 49 58
rect 41 51 49 54
rect 41 47 43 51
rect 47 47 49 51
rect 41 38 49 47
rect 51 65 59 66
rect 51 61 53 65
rect 57 61 59 65
rect 51 58 59 61
rect 51 54 53 58
rect 57 54 59 58
rect 51 38 59 54
rect 61 58 69 66
rect 61 54 63 58
rect 67 54 69 58
rect 61 51 69 54
rect 61 47 63 51
rect 67 47 69 51
rect 61 38 69 47
rect 71 63 74 66
rect 78 66 79 67
rect 78 63 81 66
rect 71 38 81 63
rect 83 59 88 66
rect 83 58 90 59
rect 83 54 85 58
rect 89 54 90 58
rect 83 51 90 54
rect 83 47 85 51
rect 89 47 90 51
rect 83 46 90 47
rect 83 38 88 46
<< metal1 >>
rect -2 67 98 72
rect -2 65 74 67
rect -2 64 53 65
rect 52 61 53 64
rect 57 64 74 65
rect 57 61 58 64
rect 73 63 74 64
rect 78 64 98 67
rect 78 63 79 64
rect 2 55 3 59
rect 7 55 23 59
rect 27 58 47 59
rect 27 55 43 58
rect 52 58 58 61
rect 52 54 53 58
rect 57 54 58 58
rect 63 58 89 59
rect 67 55 85 58
rect 43 51 47 54
rect 2 50 39 51
rect 2 46 13 50
rect 17 46 33 50
rect 37 46 39 50
rect 63 51 67 54
rect 85 51 89 54
rect 47 47 63 50
rect 43 46 67 47
rect 2 17 6 46
rect 74 42 78 51
rect 85 46 89 47
rect 10 38 42 42
rect 10 34 14 38
rect 36 34 42 38
rect 10 21 14 30
rect 18 30 23 34
rect 27 30 31 34
rect 36 30 37 34
rect 41 30 42 34
rect 49 38 86 42
rect 49 34 55 38
rect 82 34 86 38
rect 49 30 50 34
rect 54 30 55 34
rect 64 30 65 34
rect 69 30 78 34
rect 18 21 22 30
rect 33 23 67 26
rect 33 22 63 23
rect 33 17 39 22
rect 63 18 67 19
rect 2 13 23 17
rect 27 13 39 17
rect 43 16 47 17
rect 74 13 78 30
rect 82 29 86 30
rect 82 21 86 22
rect 43 8 47 12
rect 82 8 86 17
rect -2 4 5 8
rect 9 4 74 8
rect 78 4 82 8
rect 86 4 98 8
rect -2 0 98 4
<< ntransistor >>
rect 12 11 14 21
rect 19 11 21 21
rect 29 11 31 26
rect 36 11 38 26
rect 52 11 54 26
rect 59 11 61 26
rect 69 16 71 26
rect 76 16 78 26
<< ptransistor >>
rect 9 38 11 66
rect 19 38 21 66
rect 29 38 31 66
rect 39 38 41 66
rect 49 38 51 66
rect 59 38 61 66
rect 69 38 71 66
rect 81 38 83 66
<< polycontact >>
rect 10 30 14 34
rect 23 30 27 34
rect 37 30 41 34
rect 50 30 54 34
rect 65 30 69 34
rect 82 30 86 34
<< ndcontact >>
rect 23 13 27 17
rect 43 12 47 16
rect 63 19 67 23
rect 82 17 86 21
rect 5 4 9 8
<< pdcontact >>
rect 3 55 7 59
rect 13 46 17 50
rect 23 55 27 59
rect 33 46 37 50
rect 43 54 47 58
rect 43 47 47 51
rect 53 61 57 65
rect 53 54 57 58
rect 63 54 67 58
rect 63 47 67 51
rect 74 63 78 67
rect 85 54 89 58
rect 85 47 89 51
<< psubstratepcontact >>
rect 74 4 78 8
rect 82 4 86 8
<< psubstratepdiff >>
rect 73 8 87 9
rect 73 4 74 8
rect 78 4 82 8
rect 86 4 87 8
rect 73 3 87 4
<< labels >>
rlabel metal1 12 28 12 28 6 b1
rlabel metal1 4 32 4 32 6 z
rlabel metal1 12 48 12 48 6 z
rlabel metal1 20 24 20 24 6 b2
rlabel metal1 28 32 28 32 6 b2
rlabel metal1 20 40 20 40 6 b1
rlabel metal1 28 40 28 40 6 b1
rlabel metal1 20 48 20 48 6 z
rlabel metal1 28 48 28 48 6 z
rlabel metal1 48 4 48 4 6 vss
rlabel metal1 36 20 36 20 6 z
rlabel metal1 44 24 44 24 6 z
rlabel metal1 52 24 52 24 6 z
rlabel metal1 36 40 36 40 6 b1
rlabel metal1 52 36 52 36 6 a1
rlabel pdcontact 36 48 36 48 6 z
rlabel metal1 45 52 45 52 6 n3
rlabel pdcontact 24 57 24 57 6 n3
rlabel metal1 48 68 48 68 6 vdd
rlabel metal1 60 24 60 24 6 z
rlabel metal1 76 20 76 20 6 a2
rlabel polycontact 68 32 68 32 6 a2
rlabel metal1 60 40 60 40 6 a1
rlabel metal1 68 40 68 40 6 a1
rlabel metal1 76 44 76 44 6 a1
rlabel metal1 65 52 65 52 6 n3
rlabel polycontact 84 32 84 32 6 a1
rlabel metal1 87 52 87 52 6 n3
<< end >>
