magic
tech scmos
timestamp 1179385174
<< checkpaint >>
rect -22 -25 70 105
<< ab >>
rect 0 0 48 80
<< pwell >>
rect -4 -7 52 36
<< nwell >>
rect -4 36 52 87
<< polysilicon >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 37 70 39 74
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 2 38 11 39
rect 2 34 3 38
rect 7 34 11 38
rect 2 33 11 34
rect 9 30 11 33
rect 16 38 23 39
rect 16 34 18 38
rect 22 34 23 38
rect 16 33 23 34
rect 27 38 33 39
rect 27 34 28 38
rect 32 34 33 38
rect 27 33 33 34
rect 16 30 18 33
rect 27 28 29 33
rect 37 31 39 42
rect 37 30 43 31
rect 37 28 38 30
rect 26 25 29 28
rect 36 26 38 28
rect 42 26 43 30
rect 36 25 43 26
rect 26 22 28 25
rect 36 22 38 25
rect 9 16 11 21
rect 16 17 18 21
rect 26 11 28 16
rect 36 11 38 16
<< ndiffusion >>
rect 2 29 9 30
rect 2 25 3 29
rect 7 25 9 29
rect 2 24 9 25
rect 4 21 9 24
rect 11 21 16 30
rect 18 22 24 30
rect 18 21 26 22
rect 20 16 26 21
rect 28 21 36 22
rect 28 17 30 21
rect 34 17 36 21
rect 28 16 36 17
rect 38 16 46 22
rect 20 15 24 16
rect 18 14 24 15
rect 18 10 19 14
rect 23 10 24 14
rect 40 12 46 16
rect 18 9 24 10
rect 40 8 41 12
rect 45 8 46 12
rect 40 7 46 8
<< pdiffusion >>
rect 4 64 9 70
rect 2 63 9 64
rect 2 59 3 63
rect 7 59 9 63
rect 2 58 9 59
rect 4 42 9 58
rect 11 47 19 70
rect 11 43 13 47
rect 17 43 19 47
rect 11 42 19 43
rect 21 63 29 70
rect 21 59 23 63
rect 27 59 29 63
rect 21 42 29 59
rect 31 42 37 70
rect 39 69 46 70
rect 39 65 41 69
rect 45 65 46 69
rect 39 62 46 65
rect 39 58 41 62
rect 45 58 46 62
rect 39 42 46 58
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect -2 69 50 78
rect -2 68 41 69
rect 40 65 41 68
rect 45 68 50 69
rect 45 65 46 68
rect 2 59 3 63
rect 7 59 23 63
rect 27 59 28 63
rect 40 62 46 65
rect 40 58 41 62
rect 45 58 46 62
rect 2 50 15 55
rect 2 39 6 50
rect 11 43 13 47
rect 17 43 18 47
rect 25 46 31 54
rect 11 39 15 43
rect 21 42 31 46
rect 21 39 25 42
rect 42 39 46 55
rect 2 38 7 39
rect 2 34 3 38
rect 2 33 7 34
rect 10 35 15 39
rect 18 38 25 39
rect 10 29 14 35
rect 22 34 25 38
rect 18 33 25 34
rect 28 38 46 39
rect 32 34 46 38
rect 28 33 37 34
rect 2 25 3 29
rect 7 25 14 29
rect 33 26 38 30
rect 10 22 14 25
rect 10 21 36 22
rect 10 17 30 21
rect 34 17 36 21
rect 42 17 46 30
rect 18 12 19 14
rect -2 10 19 12
rect 23 12 24 14
rect 23 10 41 12
rect -2 8 41 10
rect 45 8 50 12
rect -2 2 50 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
<< ntransistor >>
rect 9 21 11 30
rect 16 21 18 30
rect 26 16 28 22
rect 36 16 38 22
<< ptransistor >>
rect 9 42 11 70
rect 19 42 21 70
rect 29 42 31 70
rect 37 42 39 70
<< polycontact >>
rect 3 34 7 38
rect 18 34 22 38
rect 28 34 32 38
rect 38 26 42 30
<< ndcontact >>
rect 3 25 7 29
rect 30 17 34 21
rect 19 10 23 14
rect 41 8 45 12
<< pdcontact >>
rect 3 59 7 63
rect 13 43 17 47
rect 23 59 27 63
rect 41 65 45 69
rect 41 58 45 62
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
<< psubstratepdiff >>
rect 0 2 48 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 48 2
rect 0 -3 48 -2
<< nsubstratendiff >>
rect 0 82 48 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 48 82
rect 0 77 48 78
<< labels >>
rlabel metal1 4 44 4 44 6 c2
rlabel metal1 12 28 12 28 6 z
rlabel metal1 12 52 12 52 6 c2
rlabel metal1 24 6 24 6 6 vss
rlabel metal1 20 20 20 20 6 z
rlabel polycontact 20 36 20 36 6 c1
rlabel metal1 15 61 15 61 6 n2
rlabel metal1 24 74 24 74 6 vdd
rlabel metal1 28 20 28 20 6 z
rlabel metal1 36 28 36 28 6 a
rlabel metal1 36 36 36 36 6 b
rlabel metal1 28 48 28 48 6 c1
rlabel metal1 44 20 44 20 6 a
rlabel metal1 44 48 44 48 6 b
<< end >>
