.subckt nd2v6x2 a b vdd vss z
*   SPICE3 file   created from nd2v6x2.ext -      technology: scmos
m00 z      a      vdd    vdd p w=28u  l=2.3636u ad=176p     pd=50u      as=196p     ps=70u
m01 vdd    b      z      vdd p w=28u  l=2.3636u ad=196p     pd=70u      as=176p     ps=50u
m02 w1     a      vss    vss n w=20u  l=2.3636u ad=136p     pd=42u      as=140p     ps=54u
m03 z      b      w1     vss n w=20u  l=2.3636u ad=140p     pd=54u      as=136p     ps=42u
C0  w1     vss    0.010f
C1  w1     z      0.037f
C2  vss    b      0.011f
C3  vss    a      0.046f
C4  b      z      0.132f
C5  z      a      0.113f
C6  b      vdd    0.042f
C7  a      vdd    0.042f
C8  vss    z      0.049f
C9  b      a      0.100f
C10 z      vdd    0.014f
C12 b      vss    0.045f
C13 z      vss    0.006f
C14 a      vss    0.045f
.ends
