.subckt na3_x4 i0 i1 i2 nq vdd vss
*   SPICE3 file   created from na3_x4.ext -      technology: scmos
m00 vdd    i0     w1     vdd p w=20u  l=2.3636u ad=105.5p   pd=35u      as=120p     ps=38.6667u
m01 w1     i2     vdd    vdd p w=20u  l=2.3636u ad=120p     pd=38.6667u as=105.5p   ps=35u
m02 vdd    i1     w1     vdd p w=20u  l=2.3636u ad=105.5p   pd=35u      as=120p     ps=38.6667u
m03 nq     w2     vdd    vdd p w=40u  l=2.3636u ad=200p     pd=50u      as=211p     ps=70u
m04 vdd    w2     nq     vdd p w=40u  l=2.3636u ad=211p     pd=70u      as=200p     ps=50u
m05 w2     w1     vdd    vdd p w=20u  l=2.3636u ad=160p     pd=56u      as=105.5p   ps=35u
m06 w3     i0     w1     vss n w=20u  l=2.3636u ad=60p      pd=26u      as=160p     ps=56u
m07 w4     i2     w3     vss n w=20u  l=2.3636u ad=60p      pd=26u      as=60p      ps=26u
m08 vss    i1     w4     vss n w=20u  l=2.3636u ad=142.857p pd=41.1429u as=60p      ps=26u
m09 nq     w2     vss    vss n w=20u  l=2.3636u ad=100p     pd=30u      as=142.857p ps=41.1429u
m10 vss    w2     nq     vss n w=20u  l=2.3636u ad=142.857p pd=41.1429u as=100p     ps=30u
m11 w2     w1     vss    vss n w=10u  l=2.3636u ad=80p      pd=36u      as=71.4286p ps=20.5714u
C0  w3     i2     0.012f
C1  nq     i1     0.095f
C2  w1     i2     0.163f
C3  nq     i0     0.039f
C4  nq     w2     0.183f
C5  i1     i0     0.127f
C6  w1     vdd    0.536f
C7  vss    nq     0.069f
C8  i2     vdd    0.032f
C9  i1     w2     0.090f
C10 w4     w1     0.012f
C11 vss    i1     0.022f
C12 i0     w2     0.012f
C13 nq     w1     0.407f
C14 w4     i2     0.004f
C15 vss    i0     0.016f
C16 vss    w2     0.074f
C17 w1     i1     0.381f
C18 nq     i2     0.056f
C19 i1     i2     0.409f
C20 w1     i0     0.162f
C21 nq     vdd    0.043f
C22 i1     vdd    0.012f
C23 i2     i0     0.419f
C24 w1     w2     0.199f
C25 vss    w1     0.288f
C26 i2     w2     0.029f
C27 i0     vdd    0.017f
C28 w3     w1     0.012f
C29 w4     i1     0.008f
C30 vss    i2     0.017f
C31 vdd    w2     0.026f
C33 nq     vss    0.018f
C34 w1     vss    0.035f
C35 i1     vss    0.037f
C36 i2     vss    0.035f
C37 i0     vss    0.033f
C39 w2     vss    0.069f
.ends
