.subckt mxi2v2x3 a0 a1 s vdd vss z
*   SPICE3 file   created from mxi2v2x3.ext -      technology: scmos
m00 a1n    a1     vdd    vdd p w=18u  l=2.3636u ad=73.0909p pd=25.6364u as=88.8462p ps=28.3846u
m01 vdd    a1     a1n    vdd p w=24u  l=2.3636u ad=118.462p pd=37.8462u as=97.4545p ps=34.1818u
m02 a1n    a1     vdd    vdd p w=24u  l=2.3636u ad=97.4545p pd=34.1818u as=118.462p ps=37.8462u
m03 z      sn     a1n    vdd p w=22u  l=2.3636u ad=88p      pd=30u      as=89.3333p ps=31.3333u
m04 a1n    sn     z      vdd p w=22u  l=2.3636u ad=89.3333p pd=31.3333u as=88p      ps=30u
m05 z      sn     a1n    vdd p w=22u  l=2.3636u ad=88p      pd=30u      as=89.3333p ps=31.3333u
m06 a0n    s      z      vdd p w=22u  l=2.3636u ad=88p      pd=30u      as=88p      ps=30u
m07 z      s      a0n    vdd p w=22u  l=2.3636u ad=88p      pd=30u      as=88p      ps=30u
m08 a0n    s      z      vdd p w=22u  l=2.3636u ad=88p      pd=30u      as=88p      ps=30u
m09 vdd    a0     a0n    vdd p w=22u  l=2.3636u ad=108.59p  pd=34.6923u as=88p      ps=30u
m10 a0n    a0     vdd    vdd p w=22u  l=2.3636u ad=88p      pd=30u      as=108.59p  ps=34.6923u
m11 vdd    a0     a0n    vdd p w=22u  l=2.3636u ad=108.59p  pd=34.6923u as=88p      ps=30u
m12 sn     s      vdd    vdd p w=24u  l=2.3636u ad=146p     pd=62u      as=118.462p ps=37.8462u
m13 a1n    a1     vss    vss n w=11u  l=2.3636u ad=49.6667p pd=22.3333u as=62.3333p ps=24.4444u
m14 vss    a1     a1n    vss n w=11u  l=2.3636u ad=62.3333p pd=24.4444u as=49.6667p ps=22.3333u
m15 a1n    a1     vss    vss n w=11u  l=2.3636u ad=49.6667p pd=22.3333u as=62.3333p ps=24.4444u
m16 z      s      a1n    vss n w=15u  l=2.3636u ad=65.9091p pd=28.6364u as=67.7273p ps=30.4545u
m17 a1n    s      z      vss n w=18u  l=2.3636u ad=81.2727p pd=36.5455u as=79.0909p ps=34.3636u
m18 a0n    sn     z      vss n w=11u  l=2.3636u ad=44p      pd=19u      as=48.3333p ps=21u
m19 z      sn     a0n    vss n w=11u  l=2.3636u ad=48.3333p pd=21u      as=44p      ps=19u
m20 a0n    sn     z      vss n w=11u  l=2.3636u ad=44p      pd=19u      as=48.3333p ps=21u
m21 vss    a0     a0n    vss n w=11u  l=2.3636u ad=62.3333p pd=24.4444u as=44p      ps=19u
m22 a0n    a0     vss    vss n w=11u  l=2.3636u ad=44p      pd=19u      as=62.3333p ps=24.4444u
m23 vss    a0     a0n    vss n w=11u  l=2.3636u ad=62.3333p pd=24.4444u as=44p      ps=19u
m24 sn     s      vss    vss n w=15u  l=2.3636u ad=87p      pd=44u      as=85p      ps=33.3333u
C0  a0n    z      0.489f
C1  vss    a0     0.036f
C2  a1     vdd    0.049f
C3  z      a0     0.027f
C4  vss    sn     0.057f
C5  a0n    a1n    0.021f
C6  z      sn     0.431f
C7  vss    s      0.123f
C8  a0n    vdd    0.124f
C9  a1n    sn     0.119f
C10 z      s      0.021f
C11 a1n    s      0.010f
C12 sn     a1     0.047f
C13 a0     vdd    0.023f
C14 vss    z      0.110f
C15 a1     s      0.026f
C16 sn     vdd    0.560f
C17 a0n    a0     0.234f
C18 vss    a1n    0.335f
C19 s      vdd    0.068f
C20 a0n    sn     0.580f
C21 vss    a1     0.041f
C22 z      a1n    0.432f
C23 a0     sn     0.135f
C24 vss    vdd    0.014f
C25 z      a1     0.018f
C26 a0n    s      0.047f
C27 z      vdd    0.058f
C28 a1n    a1     0.239f
C29 a0     s      0.218f
C30 vss    a0n    0.374f
C31 sn     s      0.429f
C32 a1n    vdd    0.315f
C34 a0n    vss    0.009f
C35 z      vss    0.024f
C36 a0     vss    0.056f
C37 a1n    vss    0.008f
C38 sn     vss    0.057f
C39 a1     vss    0.053f
C40 s      vss    0.105f
.ends
