.subckt noa2a2a2a24_x4 i0 i1 i2 i3 i4 i5 i6 i7 nq vdd vss
*   SPICE3 file   created from noa2a2a2a24_x4.ext -      technology: scmos
m00 w1     i7     w2     vdd p w=40u  l=2.3636u ad=200p     pd=50u      as=260p     ps=73u
m01 w2     i6     w1     vdd p w=40u  l=2.3636u ad=260p     pd=73u      as=200p     ps=50u
m02 w2     i5     w3     vdd p w=40u  l=2.3636u ad=260p     pd=73u      as=260p     ps=73u
m03 w3     i4     w2     vdd p w=40u  l=2.3636u ad=260p     pd=73u      as=260p     ps=73u
m04 w4     i3     w3     vdd p w=40u  l=2.3636u ad=200p     pd=50u      as=260p     ps=73u
m05 w3     i2     w4     vdd p w=40u  l=2.3636u ad=260p     pd=73u      as=200p     ps=50u
m06 w4     i1     vdd    vdd p w=40u  l=2.3636u ad=200p     pd=50u      as=240p     ps=65.7778u
m07 vdd    i0     w4     vdd p w=40u  l=2.3636u ad=240p     pd=65.7778u as=200p     ps=50u
m08 nq     w5     vdd    vdd p w=40u  l=2.3636u ad=200p     pd=50u      as=240p     ps=65.7778u
m09 vdd    w5     nq     vdd p w=40u  l=2.3636u ad=240p     pd=65.7778u as=200p     ps=50u
m10 w5     w1     vdd    vdd p w=20u  l=2.3636u ad=160p     pd=56u      as=120p     ps=32.8889u
m11 w6     i7     vss    vss n w=20u  l=2.3636u ad=100p     pd=30u      as=132.308p ps=44.3077u
m12 w1     i6     w6     vss n w=20u  l=2.3636u ad=130p     pd=43u      as=100p     ps=30u
m13 w7     i5     vss    vss n w=20u  l=2.3636u ad=60p      pd=26u      as=132.308p ps=44.3077u
m14 w1     i4     w7     vss n w=20u  l=2.3636u ad=130p     pd=43u      as=60p      ps=26u
m15 w8     i3     w1     vss n w=20u  l=2.3636u ad=60p      pd=26u      as=130p     ps=43u
m16 vss    i2     w8     vss n w=20u  l=2.3636u ad=132.308p pd=44.3077u as=60p      ps=26u
m17 w9     i1     w1     vss n w=20u  l=2.3636u ad=60p      pd=26u      as=130p     ps=43u
m18 vss    i0     w9     vss n w=20u  l=2.3636u ad=132.308p pd=44.3077u as=60p      ps=26u
m19 nq     w5     vss    vss n w=20u  l=2.3636u ad=124p     pd=38u      as=132.308p ps=44.3077u
m20 vss    w5     nq     vss n w=20u  l=2.3636u ad=132.308p pd=44.3077u as=124p     ps=38u
m21 w5     w1     vss    vss n w=10u  l=2.3636u ad=80p      pd=36u      as=66.1538p ps=22.1538u
C0  vss    i1     0.017f
C1  nq     i0     0.334f
C2  w4     w2     0.012f
C3  w3     w1     0.004f
C4  vdd    w5     0.066f
C5  w1     i7     0.273f
C6  w2     i6     0.062f
C7  i1     i3     0.047f
C8  vdd    i1     0.020f
C9  vss    i3     0.017f
C10 w4     i0     0.013f
C11 w1     w2     0.129f
C12 i2     i4     0.108f
C13 w8     w1     0.012f
C14 w1     i0     0.072f
C15 w4     i2     0.056f
C16 vss    i5     0.017f
C17 vdd    i3     0.012f
C18 i3     i5     0.108f
C19 nq     w4     0.024f
C20 w6     w1     0.016f
C21 w5     i0     0.195f
C22 w1     i2     0.036f
C23 vdd    i5     0.012f
C24 w3     i3     0.039f
C25 vss    i7     0.053f
C26 i4     i6     0.062f
C27 nq     w1     0.079f
C28 vdd    w3     0.451f
C29 w1     i4     0.065f
C30 i0     i1     0.153f
C31 w3     i5     0.020f
C32 vdd    i7     0.012f
C33 w8     vss    0.014f
C34 i5     i7     0.047f
C35 vss    i0     0.025f
C36 nq     w5     0.120f
C37 vdd    w2     0.319f
C38 i1     i2     0.065f
C39 w1     i6     0.248f
C40 w2     i5     0.050f
C41 w6     vss    0.023f
C42 w4     w5     0.004f
C43 w3     w2     0.209f
C44 vdd    i0     0.080f
C45 nq     i1     0.043f
C46 vss    i2     0.017f
C47 w2     i7     0.039f
C48 i2     i3     0.360f
C49 vss    nq     0.036f
C50 w9     w1     0.012f
C51 w1     w5     0.263f
C52 vss    i4     0.017f
C53 w4     i1     0.043f
C54 vdd    i2     0.012f
C55 i3     i4     0.332f
C56 i2     i5     0.065f
C57 w7     w1     0.012f
C58 nq     vdd    0.186f
C59 w3     i2     0.017f
C60 w4     i3     0.004f
C61 w6     i7     0.004f
C62 vss    i6     0.017f
C63 vdd    i4     0.012f
C64 w1     i1     0.047f
C65 i3     i6     0.033f
C66 i4     i5     0.360f
C67 vss    w1     1.007f
C68 vdd    w4     0.288f
C69 w5     i1     0.051f
C70 w1     i3     0.038f
C71 vdd    i6     0.012f
C72 w3     i4     0.024f
C73 w9     vss    0.014f
C74 i5     i6     0.100f
C75 vss    w5     0.075f
C76 w4     w3     0.178f
C77 vdd    w1     0.042f
C78 i0     i2     0.020f
C79 w1     i5     0.077f
C80 w2     i4     0.008f
C81 w7     vss    0.014f
C82 i6     i7     0.133f
C84 nq     vss    0.015f
C86 w4     vss    0.004f
C87 w1     vss    0.051f
C88 w2     vss    0.003f
C89 w5     vss    0.060f
C90 i0     vss    0.040f
C91 i1     vss    0.032f
C92 i2     vss    0.032f
C93 i3     vss    0.030f
C94 i4     vss    0.030f
C95 i5     vss    0.030f
C96 i6     vss    0.041f
C97 i7     vss    0.032f
.ends
