magic
tech scmos
timestamp 1179386607
<< checkpaint >>
rect -22 -25 134 105
<< ab >>
rect 0 0 112 80
<< pwell >>
rect -4 -7 116 36
<< nwell >>
rect -4 36 116 87
<< polysilicon >>
rect 10 62 12 67
rect 20 62 22 67
rect 30 62 32 67
rect 40 62 42 67
rect 50 62 52 67
rect 60 62 62 67
rect 70 62 72 67
rect 80 62 82 67
rect 90 62 92 67
rect 10 39 12 42
rect 20 39 22 42
rect 30 39 32 42
rect 10 38 32 39
rect 10 34 11 38
rect 15 34 18 38
rect 22 34 32 38
rect 10 33 32 34
rect 10 30 12 33
rect 20 30 22 33
rect 30 30 32 33
rect 40 39 42 42
rect 50 39 52 42
rect 60 39 62 42
rect 40 38 62 39
rect 40 34 42 38
rect 46 34 50 38
rect 54 34 62 38
rect 40 33 62 34
rect 40 30 42 33
rect 50 30 52 33
rect 60 30 62 33
rect 70 39 72 42
rect 80 39 82 42
rect 90 39 92 42
rect 70 38 103 39
rect 70 34 98 38
rect 102 34 103 38
rect 70 33 103 34
rect 70 30 72 33
rect 80 30 82 33
rect 90 30 92 33
rect 101 30 103 33
rect 90 15 92 20
rect 101 15 103 20
rect 10 6 12 10
rect 20 6 22 10
rect 30 6 32 10
rect 40 6 42 10
rect 50 6 52 10
rect 60 6 62 10
rect 70 6 72 10
rect 80 6 82 10
<< ndiffusion >>
rect 2 22 10 30
rect 2 18 3 22
rect 7 18 10 22
rect 2 15 10 18
rect 2 11 3 15
rect 7 11 10 15
rect 2 10 10 11
rect 12 29 20 30
rect 12 25 14 29
rect 18 25 20 29
rect 12 22 20 25
rect 12 18 14 22
rect 18 18 20 22
rect 12 10 20 18
rect 22 15 30 30
rect 22 11 24 15
rect 28 11 30 15
rect 22 10 30 11
rect 32 22 40 30
rect 32 18 34 22
rect 38 18 40 22
rect 32 10 40 18
rect 42 29 50 30
rect 42 25 44 29
rect 48 25 50 29
rect 42 10 50 25
rect 52 22 60 30
rect 52 18 54 22
rect 58 18 60 22
rect 52 10 60 18
rect 62 29 70 30
rect 62 25 64 29
rect 68 25 70 29
rect 62 22 70 25
rect 62 18 64 22
rect 68 18 70 22
rect 62 10 70 18
rect 72 29 80 30
rect 72 25 74 29
rect 78 25 80 29
rect 72 10 80 25
rect 82 25 90 30
rect 82 21 84 25
rect 88 21 90 25
rect 82 20 90 21
rect 92 29 101 30
rect 92 25 94 29
rect 98 25 101 29
rect 92 20 101 25
rect 103 26 108 30
rect 103 25 110 26
rect 103 21 105 25
rect 109 21 110 25
rect 103 20 110 21
rect 82 10 87 20
<< pdiffusion >>
rect 2 61 10 62
rect 2 57 3 61
rect 7 57 10 61
rect 2 54 10 57
rect 2 50 3 54
rect 7 50 10 54
rect 2 42 10 50
rect 12 54 20 62
rect 12 50 14 54
rect 18 50 20 54
rect 12 47 20 50
rect 12 43 14 47
rect 18 43 20 47
rect 12 42 20 43
rect 22 61 30 62
rect 22 57 24 61
rect 28 57 30 61
rect 22 54 30 57
rect 22 50 24 54
rect 28 50 30 54
rect 22 42 30 50
rect 32 54 40 62
rect 32 50 34 54
rect 38 50 40 54
rect 32 47 40 50
rect 32 43 34 47
rect 38 43 40 47
rect 32 42 40 43
rect 42 61 50 62
rect 42 57 44 61
rect 48 57 50 61
rect 42 54 50 57
rect 42 50 44 54
rect 48 50 50 54
rect 42 42 50 50
rect 52 54 60 62
rect 52 50 54 54
rect 58 50 60 54
rect 52 47 60 50
rect 52 43 54 47
rect 58 43 60 47
rect 52 42 60 43
rect 62 61 70 62
rect 62 57 64 61
rect 68 57 70 61
rect 62 54 70 57
rect 62 50 64 54
rect 68 50 70 54
rect 62 42 70 50
rect 72 54 80 62
rect 72 50 74 54
rect 78 50 80 54
rect 72 47 80 50
rect 72 43 74 47
rect 78 43 80 47
rect 72 42 80 43
rect 82 61 90 62
rect 82 57 84 61
rect 88 57 90 61
rect 82 54 90 57
rect 82 50 84 54
rect 88 50 90 54
rect 82 42 90 50
rect 92 55 97 62
rect 92 54 99 55
rect 92 50 94 54
rect 98 50 99 54
rect 92 47 99 50
rect 92 43 94 47
rect 98 43 99 47
rect 92 42 99 43
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect -2 68 114 78
rect 2 61 8 68
rect 2 57 3 61
rect 7 57 8 61
rect 2 54 8 57
rect 23 61 29 68
rect 23 57 24 61
rect 28 57 29 61
rect 2 50 3 54
rect 7 50 8 54
rect 14 54 18 55
rect 23 54 29 57
rect 43 61 49 68
rect 43 57 44 61
rect 48 57 49 61
rect 23 50 24 54
rect 28 50 29 54
rect 34 54 38 55
rect 43 54 49 57
rect 63 61 69 68
rect 63 57 64 61
rect 68 57 69 61
rect 43 50 44 54
rect 48 50 49 54
rect 54 54 58 55
rect 63 54 69 57
rect 63 50 64 54
rect 68 50 69 54
rect 74 54 78 63
rect 83 61 89 68
rect 83 57 84 61
rect 88 57 89 61
rect 83 54 89 57
rect 83 50 84 54
rect 88 50 89 54
rect 94 54 98 55
rect 14 47 18 50
rect 2 38 6 47
rect 34 47 38 50
rect 18 43 34 46
rect 54 47 58 50
rect 38 43 54 46
rect 74 47 78 50
rect 94 47 98 50
rect 58 43 74 46
rect 90 46 94 47
rect 78 43 94 46
rect 14 42 98 43
rect 74 41 95 42
rect 2 34 11 38
rect 15 34 18 38
rect 22 34 23 38
rect 33 34 42 38
rect 46 34 50 38
rect 54 34 55 38
rect 2 25 6 34
rect 13 29 18 30
rect 13 25 14 29
rect 33 26 39 34
rect 74 29 78 41
rect 43 25 44 29
rect 48 25 64 29
rect 68 25 69 29
rect 13 22 18 25
rect 64 22 69 25
rect 91 29 95 41
rect 106 39 110 55
rect 98 38 110 39
rect 102 34 110 38
rect 98 33 110 34
rect 74 24 78 25
rect 84 25 88 26
rect 91 25 94 29
rect 98 25 99 29
rect 105 25 109 26
rect 2 18 3 22
rect 7 18 8 22
rect 13 18 14 22
rect 18 18 34 22
rect 38 18 54 22
rect 58 18 59 22
rect 68 21 69 22
rect 68 18 109 21
rect 2 15 8 18
rect 64 17 109 18
rect 2 12 3 15
rect -2 11 3 12
rect 7 12 8 15
rect 23 12 24 15
rect 7 11 24 12
rect 28 12 29 15
rect 28 11 114 12
rect -2 2 114 11
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
<< ntransistor >>
rect 10 10 12 30
rect 20 10 22 30
rect 30 10 32 30
rect 40 10 42 30
rect 50 10 52 30
rect 60 10 62 30
rect 70 10 72 30
rect 80 10 82 30
rect 90 20 92 30
rect 101 20 103 30
<< ptransistor >>
rect 10 42 12 62
rect 20 42 22 62
rect 30 42 32 62
rect 40 42 42 62
rect 50 42 52 62
rect 60 42 62 62
rect 70 42 72 62
rect 80 42 82 62
rect 90 42 92 62
<< polycontact >>
rect 11 34 15 38
rect 18 34 22 38
rect 42 34 46 38
rect 50 34 54 38
rect 98 34 102 38
<< ndcontact >>
rect 3 18 7 22
rect 3 11 7 15
rect 14 25 18 29
rect 14 18 18 22
rect 24 11 28 15
rect 34 18 38 22
rect 44 25 48 29
rect 54 18 58 22
rect 64 25 68 29
rect 64 18 68 22
rect 74 25 78 29
rect 84 21 88 25
rect 94 25 98 29
rect 105 21 109 25
<< pdcontact >>
rect 3 57 7 61
rect 3 50 7 54
rect 14 50 18 54
rect 14 43 18 47
rect 24 57 28 61
rect 24 50 28 54
rect 34 50 38 54
rect 34 43 38 47
rect 44 57 48 61
rect 44 50 48 54
rect 54 50 58 54
rect 54 43 58 47
rect 64 57 68 61
rect 64 50 68 54
rect 74 50 78 54
rect 74 43 78 47
rect 84 57 88 61
rect 84 50 88 54
rect 94 50 98 54
rect 94 43 98 47
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
rect 90 -2 94 2
rect 98 -2 102 2
rect 106 -2 110 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
rect 90 78 94 82
rect 98 78 102 82
rect 106 78 110 82
<< psubstratepdiff >>
rect 0 2 112 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 112 2
rect 0 -3 112 -2
<< nsubstratendiff >>
rect 0 82 112 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 112 82
rect 0 77 112 78
<< labels >>
rlabel metal1 15 24 15 24 6 n1
rlabel polycontact 12 36 12 36 6 a
rlabel metal1 4 36 4 36 6 a
rlabel metal1 36 32 36 32 6 b
rlabel metal1 20 44 20 44 6 z
rlabel polycontact 20 36 20 36 6 a
rlabel metal1 28 44 28 44 6 z
rlabel metal1 36 48 36 48 6 z
rlabel metal1 56 6 56 6 6 vss
rlabel ndcontact 36 20 36 20 6 n1
rlabel metal1 44 44 44 44 6 z
rlabel polycontact 44 36 44 36 6 b
rlabel metal1 52 44 52 44 6 z
rlabel metal1 60 44 60 44 6 z
rlabel polycontact 52 36 52 36 6 b
rlabel metal1 56 74 56 74 6 vdd
rlabel metal1 66 23 66 23 6 n2
rlabel metal1 56 27 56 27 6 n2
rlabel metal1 86 21 86 21 6 n2
rlabel metal1 68 44 68 44 6 z
rlabel pdcontact 76 44 76 44 6 z
rlabel metal1 84 44 84 44 6 z
rlabel metal1 107 21 107 21 6 n2
rlabel metal1 92 44 92 44 6 z
rlabel metal1 108 44 108 44 6 c
rlabel polycontact 100 36 100 36 6 c
<< end >>
