magic
tech scmos
timestamp 1179387008
<< checkpaint >>
rect -22 -22 62 94
<< ab >>
rect 0 0 40 72
<< pwell >>
rect -4 -4 44 32
<< nwell >>
rect -4 32 44 76
<< polysilicon >>
rect 12 62 14 67
rect 22 62 24 67
rect 29 62 31 67
rect 12 45 14 54
rect 9 44 15 45
rect 9 40 10 44
rect 14 40 15 44
rect 9 39 15 40
rect 9 26 11 39
rect 22 35 24 46
rect 18 34 24 35
rect 18 30 19 34
rect 23 30 24 34
rect 18 29 24 30
rect 29 43 31 46
rect 29 42 35 43
rect 29 38 30 42
rect 34 38 35 42
rect 29 37 35 38
rect 19 26 21 29
rect 9 14 11 19
rect 19 14 21 19
rect 29 18 31 37
rect 29 6 31 11
<< ndiffusion >>
rect 2 24 9 26
rect 2 20 3 24
rect 7 20 9 24
rect 2 19 9 20
rect 11 24 19 26
rect 11 20 13 24
rect 17 20 19 24
rect 11 19 19 20
rect 21 19 27 26
rect 23 18 27 19
rect 23 12 29 18
rect 21 11 29 12
rect 31 17 38 18
rect 31 13 33 17
rect 37 13 38 17
rect 31 11 38 13
rect 21 8 27 11
rect 21 4 22 8
rect 26 4 27 8
rect 21 3 27 4
<< pdiffusion >>
rect 3 68 10 69
rect 3 64 5 68
rect 9 64 10 68
rect 3 62 10 64
rect 3 54 12 62
rect 14 59 22 62
rect 14 55 16 59
rect 20 55 22 59
rect 14 54 22 55
rect 17 46 22 54
rect 24 46 29 62
rect 31 59 38 62
rect 31 55 33 59
rect 37 55 38 59
rect 31 46 38 55
<< metal1 >>
rect -2 68 42 72
rect -2 64 5 68
rect 9 64 42 68
rect 32 59 38 64
rect 2 55 16 59
rect 20 55 23 59
rect 32 55 33 59
rect 37 55 38 59
rect 2 54 23 55
rect 2 25 6 54
rect 10 46 23 50
rect 10 44 14 46
rect 10 29 14 40
rect 25 38 30 42
rect 34 38 38 51
rect 18 30 19 34
rect 23 30 31 34
rect 25 27 31 30
rect 2 24 7 25
rect 2 20 3 24
rect 2 19 7 20
rect 13 24 17 25
rect 25 21 38 27
rect 2 13 6 19
rect 13 17 17 20
rect 13 13 33 17
rect 37 13 38 17
rect -2 4 4 8
rect 8 4 12 8
rect 16 4 22 8
rect 26 4 42 8
rect -2 0 42 4
<< ntransistor >>
rect 9 19 11 26
rect 19 19 21 26
rect 29 11 31 18
<< ptransistor >>
rect 12 54 14 62
rect 22 46 24 62
rect 29 46 31 62
<< polycontact >>
rect 10 40 14 44
rect 19 30 23 34
rect 30 38 34 42
<< ndcontact >>
rect 3 20 7 24
rect 13 20 17 24
rect 33 13 37 17
rect 22 4 26 8
<< pdcontact >>
rect 5 64 9 68
rect 16 55 20 59
rect 33 55 37 59
<< psubstratepcontact >>
rect 4 4 8 8
rect 12 4 16 8
<< psubstratepdiff >>
rect 3 8 17 9
rect 3 4 4 8
rect 8 4 12 8
rect 16 4 17 8
rect 3 3 17 4
<< labels >>
rlabel metal1 4 36 4 36 6 z
rlabel metal1 15 19 15 19 6 n1
rlabel metal1 12 36 12 36 6 b
rlabel metal1 12 56 12 56 6 z
rlabel metal1 20 4 20 4 6 vss
rlabel metal1 28 28 28 28 6 a2
rlabel metal1 28 40 28 40 6 a1
rlabel metal1 20 48 20 48 6 b
rlabel metal1 20 56 20 56 6 z
rlabel metal1 20 68 20 68 6 vdd
rlabel metal1 25 15 25 15 6 n1
rlabel metal1 36 24 36 24 6 a2
rlabel metal1 36 48 36 48 6 a1
<< end >>
