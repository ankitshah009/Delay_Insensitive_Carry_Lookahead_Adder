magic
tech scmos
timestamp 1180600839
<< checkpaint >>
rect -22 -22 122 122
<< ab >>
rect 0 0 100 100
<< pwell >>
rect -4 -4 104 48
<< nwell >>
rect -4 48 104 104
<< polysilicon >>
rect 11 94 13 98
rect 23 94 25 98
rect 35 94 37 98
rect 63 85 65 89
rect 75 85 77 89
rect 87 86 89 90
rect 35 63 37 75
rect 45 66 51 67
rect 35 62 41 63
rect 35 58 36 62
rect 40 58 41 62
rect 45 62 46 66
rect 50 63 51 66
rect 63 63 65 66
rect 50 62 65 63
rect 45 61 65 62
rect 35 57 41 58
rect 75 57 77 65
rect 87 63 89 66
rect 81 62 89 63
rect 81 58 82 62
rect 86 58 89 62
rect 81 57 89 58
rect 35 56 77 57
rect 35 55 66 56
rect 11 47 13 55
rect 23 47 25 55
rect 65 52 66 55
rect 70 55 77 56
rect 70 52 71 55
rect 65 51 71 52
rect 91 48 97 49
rect 91 47 92 48
rect 11 45 92 47
rect 91 44 92 45
rect 96 44 97 48
rect 91 43 97 44
rect 11 38 61 39
rect 11 37 56 38
rect 11 25 13 37
rect 23 25 25 37
rect 55 34 56 37
rect 60 34 61 38
rect 55 33 61 34
rect 65 38 89 39
rect 65 34 66 38
rect 70 37 89 38
rect 70 34 71 37
rect 65 33 71 34
rect 29 32 37 33
rect 29 28 30 32
rect 34 28 37 32
rect 29 27 37 28
rect 45 32 51 33
rect 45 28 46 32
rect 50 29 51 32
rect 75 32 83 33
rect 50 28 65 29
rect 45 27 65 28
rect 35 24 37 27
rect 63 24 65 27
rect 75 28 78 32
rect 82 28 83 32
rect 75 27 83 28
rect 75 24 77 27
rect 87 25 89 37
rect 35 11 37 15
rect 63 11 65 15
rect 11 2 13 6
rect 23 2 25 6
rect 75 11 77 15
rect 87 11 89 15
<< ndiffusion >>
rect 3 22 11 25
rect 3 18 4 22
rect 8 18 11 22
rect 3 12 11 18
rect 3 8 4 12
rect 8 8 11 12
rect 3 6 11 8
rect 13 22 23 25
rect 13 18 16 22
rect 20 18 23 22
rect 13 6 23 18
rect 25 24 30 25
rect 82 24 87 25
rect 25 15 35 24
rect 37 22 45 24
rect 37 18 40 22
rect 44 18 45 22
rect 37 15 45 18
rect 55 22 63 24
rect 55 18 56 22
rect 60 18 63 22
rect 55 15 63 18
rect 65 15 75 24
rect 77 22 87 24
rect 77 18 80 22
rect 84 18 87 22
rect 77 15 87 18
rect 89 22 97 25
rect 89 18 92 22
rect 96 18 97 22
rect 89 15 97 18
rect 25 12 33 15
rect 25 8 28 12
rect 32 8 33 12
rect 67 12 73 15
rect 25 6 33 8
rect 67 8 68 12
rect 72 8 73 12
rect 67 7 73 8
<< pdiffusion >>
rect 3 92 11 94
rect 3 88 4 92
rect 8 88 11 92
rect 3 82 11 88
rect 3 78 4 82
rect 8 78 11 82
rect 3 72 11 78
rect 3 68 4 72
rect 8 68 11 72
rect 3 62 11 68
rect 3 58 4 62
rect 8 58 11 62
rect 3 55 11 58
rect 13 82 23 94
rect 13 78 16 82
rect 20 78 23 82
rect 13 72 23 78
rect 13 68 16 72
rect 20 68 23 72
rect 13 62 23 68
rect 13 58 16 62
rect 20 58 23 62
rect 13 55 23 58
rect 25 92 35 94
rect 25 88 28 92
rect 32 88 35 92
rect 25 75 35 88
rect 37 82 45 94
rect 79 92 85 94
rect 79 88 80 92
rect 84 88 85 92
rect 79 86 85 88
rect 79 85 87 86
rect 37 78 40 82
rect 44 78 45 82
rect 37 75 45 78
rect 55 82 63 85
rect 55 78 56 82
rect 60 78 63 82
rect 25 55 33 75
rect 55 72 63 78
rect 55 68 56 72
rect 60 68 63 72
rect 55 66 63 68
rect 65 82 75 85
rect 65 78 68 82
rect 72 78 75 82
rect 65 72 75 78
rect 65 68 68 72
rect 72 68 75 72
rect 65 66 75 68
rect 70 65 75 66
rect 77 66 87 85
rect 89 82 97 86
rect 89 78 92 82
rect 96 78 97 82
rect 89 72 97 78
rect 89 68 92 72
rect 96 68 97 72
rect 89 66 97 68
rect 77 65 82 66
<< metal1 >>
rect -2 96 102 100
rect -2 92 52 96
rect 56 92 68 96
rect 72 92 102 96
rect -2 88 4 92
rect 8 88 28 92
rect 32 88 80 92
rect 84 88 102 92
rect 4 82 8 88
rect 18 82 22 83
rect 15 78 16 82
rect 20 78 22 82
rect 4 72 8 78
rect 18 72 22 78
rect 15 68 16 72
rect 20 68 22 72
rect 4 62 8 68
rect 18 62 22 68
rect 15 58 16 62
rect 20 58 22 62
rect 4 57 8 58
rect 4 22 8 23
rect 18 22 22 58
rect 15 18 16 22
rect 20 18 22 22
rect 4 12 8 18
rect 18 17 22 18
rect 28 62 32 83
rect 56 82 60 83
rect 39 78 40 82
rect 44 78 50 82
rect 46 66 50 78
rect 28 58 36 62
rect 40 58 41 62
rect 28 32 32 58
rect 46 32 50 62
rect 28 28 30 32
rect 34 28 35 32
rect 28 17 32 28
rect 46 22 50 28
rect 39 18 40 22
rect 44 18 50 22
rect 56 72 60 78
rect 56 38 60 68
rect 68 82 72 83
rect 92 82 96 83
rect 72 78 92 82
rect 68 72 72 78
rect 68 67 72 68
rect 56 22 60 34
rect 66 56 70 57
rect 66 38 70 52
rect 66 33 70 34
rect 78 32 82 73
rect 92 72 96 78
rect 86 58 87 62
rect 78 27 82 28
rect 92 48 96 68
rect 92 22 96 44
rect 60 18 80 22
rect 84 18 85 22
rect 56 17 60 18
rect 92 17 96 18
rect -2 8 4 12
rect 8 8 28 12
rect 32 8 68 12
rect 72 8 102 12
rect -2 4 40 8
rect 44 4 56 8
rect 60 4 80 8
rect 84 4 92 8
rect 96 4 102 8
rect -2 0 102 4
<< ntransistor >>
rect 11 6 13 25
rect 23 6 25 25
rect 35 15 37 24
rect 63 15 65 24
rect 75 15 77 24
rect 87 15 89 25
<< ptransistor >>
rect 11 55 13 94
rect 23 55 25 94
rect 35 75 37 94
rect 63 66 65 85
rect 75 65 77 85
rect 87 66 89 86
<< polycontact >>
rect 36 58 40 62
rect 46 62 50 66
rect 82 58 86 62
rect 66 52 70 56
rect 92 44 96 48
rect 56 34 60 38
rect 66 34 70 38
rect 30 28 34 32
rect 46 28 50 32
rect 78 28 82 32
<< ndcontact >>
rect 4 18 8 22
rect 4 8 8 12
rect 16 18 20 22
rect 40 18 44 22
rect 56 18 60 22
rect 80 18 84 22
rect 92 18 96 22
rect 28 8 32 12
rect 68 8 72 12
<< pdcontact >>
rect 4 88 8 92
rect 4 78 8 82
rect 4 68 8 72
rect 4 58 8 62
rect 16 78 20 82
rect 16 68 20 72
rect 16 58 20 62
rect 28 88 32 92
rect 80 88 84 92
rect 40 78 44 82
rect 56 78 60 82
rect 56 68 60 72
rect 68 78 72 82
rect 68 68 72 72
rect 92 78 96 82
rect 92 68 96 72
<< psubstratepcontact >>
rect 40 4 44 8
rect 56 4 60 8
rect 80 4 84 8
rect 92 4 96 8
<< nsubstratencontact >>
rect 52 92 56 96
rect 68 92 72 96
<< psubstratepdiff >>
rect 39 8 61 9
rect 39 4 40 8
rect 44 4 56 8
rect 60 4 61 8
rect 79 8 97 9
rect 39 3 61 4
rect 79 4 80 8
rect 84 4 92 8
rect 96 4 97 8
rect 79 3 97 4
<< nsubstratendiff >>
rect 51 96 73 97
rect 51 92 52 96
rect 56 92 68 96
rect 72 92 73 96
rect 51 91 73 92
<< labels >>
rlabel metal1 20 50 20 50 6 q
rlabel metal1 30 50 30 50 6 cmd
rlabel metal1 50 6 50 6 6 vss
rlabel metal1 50 94 50 94 6 vdd
rlabel metal1 80 50 80 50 6 i
<< end >>
