magic
tech scmos
timestamp 1179385857
<< checkpaint >>
rect -22 -25 78 105
<< ab >>
rect 0 0 56 80
<< pwell >>
rect -4 -7 60 36
<< nwell >>
rect -4 36 60 87
<< polysilicon >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 39 62 41 67
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 39 39 41 42
rect 9 38 41 39
rect 9 37 27 38
rect 9 30 11 37
rect 19 30 21 37
rect 26 34 27 37
rect 31 34 36 38
rect 40 34 41 38
rect 26 33 41 34
rect 29 30 31 33
rect 39 30 41 33
rect 9 15 11 20
rect 19 11 21 16
rect 29 11 31 16
rect 39 11 41 16
<< ndiffusion >>
rect 2 25 9 30
rect 2 21 3 25
rect 7 21 9 25
rect 2 20 9 21
rect 11 29 19 30
rect 11 25 13 29
rect 17 25 19 29
rect 11 20 19 25
rect 14 16 19 20
rect 21 21 29 30
rect 21 17 23 21
rect 27 17 29 21
rect 21 16 29 17
rect 31 29 39 30
rect 31 25 33 29
rect 37 25 39 29
rect 31 22 39 25
rect 31 18 33 22
rect 37 18 39 22
rect 31 16 39 18
rect 41 29 48 30
rect 41 25 43 29
rect 47 25 48 29
rect 41 21 48 25
rect 41 17 43 21
rect 47 17 48 21
rect 41 16 48 17
<< pdiffusion >>
rect 2 69 9 70
rect 2 65 3 69
rect 7 65 9 69
rect 2 62 9 65
rect 2 58 3 62
rect 7 58 9 62
rect 2 42 9 58
rect 11 54 19 70
rect 11 50 13 54
rect 17 50 19 54
rect 11 47 19 50
rect 11 43 13 47
rect 17 43 19 47
rect 11 42 19 43
rect 21 69 29 70
rect 21 65 23 69
rect 27 65 29 69
rect 21 61 29 65
rect 21 57 23 61
rect 27 57 29 61
rect 21 42 29 57
rect 31 62 36 70
rect 31 54 39 62
rect 31 50 33 54
rect 37 50 39 54
rect 31 47 39 50
rect 31 43 33 47
rect 37 43 39 47
rect 31 42 39 43
rect 41 61 48 62
rect 41 57 43 61
rect 47 57 48 61
rect 41 54 48 57
rect 41 50 43 54
rect 47 50 48 54
rect 41 42 48 50
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect -2 69 58 78
rect -2 68 3 69
rect 2 65 3 68
rect 7 68 23 69
rect 7 65 8 68
rect 2 62 8 65
rect 2 58 3 62
rect 7 58 8 62
rect 27 68 58 69
rect 23 61 27 65
rect 23 56 27 57
rect 42 61 48 68
rect 42 57 43 61
rect 47 57 48 61
rect 13 54 17 55
rect 13 47 17 50
rect 10 43 13 47
rect 33 54 38 55
rect 37 50 38 54
rect 42 54 48 57
rect 42 50 43 54
rect 47 50 48 54
rect 33 47 38 50
rect 17 43 33 46
rect 37 43 38 47
rect 10 42 38 43
rect 10 30 14 42
rect 42 38 47 47
rect 25 34 27 38
rect 31 34 36 38
rect 40 34 47 38
rect 10 29 38 30
rect 3 25 7 26
rect 10 25 13 29
rect 17 26 33 29
rect 17 25 18 26
rect 37 25 38 29
rect 33 22 38 25
rect 3 12 7 21
rect 23 21 27 22
rect 37 18 38 22
rect 33 17 38 18
rect 43 29 47 30
rect 43 21 47 25
rect 23 12 27 17
rect 43 12 47 17
rect -2 2 58 12
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
<< ntransistor >>
rect 9 20 11 30
rect 19 16 21 30
rect 29 16 31 30
rect 39 16 41 30
<< ptransistor >>
rect 9 42 11 70
rect 19 42 21 70
rect 29 42 31 70
rect 39 42 41 62
<< polycontact >>
rect 27 34 31 38
rect 36 34 40 38
<< ndcontact >>
rect 3 21 7 25
rect 13 25 17 29
rect 23 17 27 21
rect 33 25 37 29
rect 33 18 37 22
rect 43 25 47 29
rect 43 17 47 21
<< pdcontact >>
rect 3 65 7 69
rect 3 58 7 62
rect 13 50 17 54
rect 13 43 17 47
rect 23 65 27 69
rect 23 57 27 61
rect 33 50 37 54
rect 33 43 37 47
rect 43 57 47 61
rect 43 50 47 54
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
<< psubstratepdiff >>
rect 0 2 56 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 56 2
rect 0 -3 56 -2
<< nsubstratendiff >>
rect 0 82 56 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 56 82
rect 0 77 56 78
<< labels >>
rlabel metal1 12 36 12 36 6 z
rlabel metal1 20 28 20 28 6 z
rlabel metal1 20 44 20 44 6 z
rlabel metal1 28 6 28 6 6 vss
rlabel ndcontact 36 20 36 20 6 z
rlabel metal1 28 28 28 28 6 z
rlabel polycontact 28 36 28 36 6 a
rlabel metal1 36 36 36 36 6 a
rlabel metal1 28 44 28 44 6 z
rlabel pdcontact 36 52 36 52 6 z
rlabel metal1 28 74 28 74 6 vdd
rlabel metal1 44 40 44 40 6 a
<< end >>
