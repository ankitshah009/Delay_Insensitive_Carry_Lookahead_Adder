magic
tech scmos
timestamp 1185094829
<< checkpaint >>
rect -22 -22 92 122
<< ab >>
rect 0 0 70 100
<< pwell >>
rect -4 -4 74 48
<< nwell >>
rect -4 48 74 104
<< metal1 >>
rect -2 96 72 100
rect -2 92 4 96
rect 8 92 13 96
rect 17 92 23 96
rect 27 92 33 96
rect 37 92 43 96
rect 47 92 53 96
rect 57 92 62 96
rect 66 92 72 96
rect -2 88 72 92
rect -2 8 72 12
rect -2 4 4 8
rect 8 4 13 8
rect 17 4 23 8
rect 27 4 33 8
rect 37 4 43 8
rect 47 4 53 8
rect 57 4 62 8
rect 66 4 72 8
rect -2 0 72 4
<< psubstratepcontact >>
rect 4 4 8 8
rect 13 4 17 8
rect 23 4 27 8
rect 33 4 37 8
rect 43 4 47 8
rect 53 4 57 8
rect 62 4 66 8
<< nsubstratencontact >>
rect 4 92 8 96
rect 13 92 17 96
rect 23 92 27 96
rect 33 92 37 96
rect 43 92 47 96
rect 53 92 57 96
rect 62 92 66 96
<< psubstratepdiff >>
rect 3 8 67 39
rect 3 4 4 8
rect 8 4 13 8
rect 17 4 23 8
rect 27 4 33 8
rect 37 4 43 8
rect 47 4 53 8
rect 57 4 62 8
rect 66 4 67 8
rect 3 3 67 4
<< nsubstratendiff >>
rect 3 96 67 97
rect 3 92 4 96
rect 8 92 13 96
rect 17 92 23 96
rect 27 92 33 96
rect 37 92 43 96
rect 47 92 53 96
rect 57 92 62 96
rect 66 92 67 96
rect 3 55 67 92
<< labels >>
rlabel psubstratepcontact 35 6 35 6 6 vss
rlabel nsubstratencontact 35 94 35 94 6 vdd
<< end >>
