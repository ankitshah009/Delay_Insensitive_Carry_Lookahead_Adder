.subckt aon21v0x05 a1 a2 b vdd vss z
*   SPICE3 file   created from aon21v0x05.ext -      technology: scmos
m00 vdd    w1     z      vdd p w=12u  l=2.3636u ad=81.2727p pd=29.4545u as=72p      ps=38u
m01 n1     b      w1     vdd p w=16u  l=2.3636u ad=73.3333p pd=31.3333u as=106p     ps=46u
m02 vdd    a2     n1     vdd p w=16u  l=2.3636u ad=108.364p pd=39.2727u as=73.3333p ps=31.3333u
m03 n1     a1     vdd    vdd p w=16u  l=2.3636u ad=73.3333p pd=31.3333u as=108.364p ps=39.2727u
m04 vss    w1     z      vss n w=6u   l=2.3636u ad=59.0526p pd=27.1579u as=42p      ps=26u
m05 w1     b      vss    vss n w=6u   l=2.3636u ad=24.4615p pd=13.8462u as=59.0526p ps=27.1579u
m06 w2     a2     w1     vss n w=7u   l=2.3636u ad=17.5p    pd=12u      as=28.5385p ps=16.1538u
m07 vss    a1     w2     vss n w=7u   l=2.3636u ad=68.8947p pd=31.6842u as=17.5p    ps=12u
C0  w1     b      0.240f
C1  z      vdd    0.015f
C2  a1     a2     0.096f
C3  a1     vdd    0.047f
C4  a2     b      0.146f
C5  vss    z      0.098f
C6  b      vdd    0.055f
C7  n1     w1     0.017f
C8  vss    a1     0.015f
C9  n1     a2     0.021f
C10 vss    b      0.017f
C11 n1     vdd    0.197f
C12 z      b      0.017f
C13 w1     a2     0.070f
C14 w1     vdd    0.096f
C15 a1     b      0.093f
C16 vss    n1     0.003f
C17 a2     vdd    0.014f
C18 vss    w1     0.221f
C19 n1     a1     0.108f
C20 z      w1     0.082f
C21 vss    a2     0.053f
C22 w1     a1     0.025f
C23 n1     b      0.111f
C24 vss    vdd    0.006f
C25 z      a2     0.012f
C27 z      vss    0.013f
C28 w1     vss    0.035f
C29 a1     vss    0.029f
C30 a2     vss    0.025f
C31 b      vss    0.025f
.ends
