magic
tech scmos
timestamp 1179387151
<< checkpaint >>
rect -22 -25 62 105
<< ab >>
rect 0 0 40 80
<< pwell >>
rect -4 -7 44 36
<< nwell >>
rect -4 36 44 87
<< polysilicon >>
rect 22 70 24 74
rect 29 70 31 74
rect 9 61 11 65
rect 9 40 11 49
rect 22 47 24 52
rect 19 46 25 47
rect 19 42 20 46
rect 24 42 25 46
rect 19 41 25 42
rect 9 39 15 40
rect 9 35 10 39
rect 14 35 15 39
rect 9 34 15 35
rect 9 25 11 34
rect 19 25 21 41
rect 29 39 31 52
rect 29 38 35 39
rect 29 34 30 38
rect 34 34 35 38
rect 29 33 35 34
rect 29 25 31 33
rect 9 15 11 19
rect 19 15 21 19
rect 29 15 31 19
<< ndiffusion >>
rect 2 24 9 25
rect 2 20 3 24
rect 7 20 9 24
rect 2 19 9 20
rect 11 24 19 25
rect 11 20 13 24
rect 17 20 19 24
rect 11 19 19 20
rect 21 24 29 25
rect 21 20 23 24
rect 27 20 29 24
rect 21 19 29 20
rect 31 24 38 25
rect 31 20 33 24
rect 37 20 38 24
rect 31 19 38 20
<< pdiffusion >>
rect 13 69 22 70
rect 13 65 15 69
rect 19 65 22 69
rect 13 61 22 65
rect 2 60 9 61
rect 2 56 3 60
rect 7 56 9 60
rect 2 55 9 56
rect 4 49 9 55
rect 11 52 22 61
rect 24 52 29 70
rect 31 63 36 70
rect 31 62 38 63
rect 31 58 33 62
rect 37 58 38 62
rect 31 57 38 58
rect 31 52 36 57
rect 11 49 19 52
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect -2 69 42 78
rect -2 68 15 69
rect 14 65 15 68
rect 19 68 42 69
rect 19 65 20 68
rect 2 60 15 62
rect 2 56 3 60
rect 7 58 15 60
rect 18 58 33 62
rect 37 58 38 62
rect 2 55 7 56
rect 2 25 6 55
rect 18 54 22 58
rect 10 50 22 54
rect 10 39 14 50
rect 26 46 30 55
rect 17 42 20 46
rect 24 42 30 46
rect 10 31 14 35
rect 25 34 30 38
rect 34 33 38 47
rect 10 27 27 31
rect 2 24 7 25
rect 23 24 27 27
rect 2 20 3 24
rect 2 17 7 20
rect 12 20 13 24
rect 17 20 18 24
rect 12 12 18 20
rect 23 19 27 20
rect 32 20 33 24
rect 37 20 38 24
rect 32 12 38 20
rect -2 2 42 12
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
<< ntransistor >>
rect 9 19 11 25
rect 19 19 21 25
rect 29 19 31 25
<< ptransistor >>
rect 9 49 11 61
rect 22 52 24 70
rect 29 52 31 70
<< polycontact >>
rect 20 42 24 46
rect 10 35 14 39
rect 30 34 34 38
<< ndcontact >>
rect 3 20 7 24
rect 13 20 17 24
rect 23 20 27 24
rect 33 20 37 24
<< pdcontact >>
rect 15 65 19 69
rect 3 56 7 60
rect 33 58 37 62
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
<< psubstratepdiff >>
rect 0 2 40 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 40 2
rect 0 -3 40 -2
<< nsubstratendiff >>
rect 0 82 40 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 40 82
rect 0 77 40 78
<< labels >>
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 40 12 40 6 zn
rlabel metal1 12 60 12 60 6 z
rlabel metal1 20 6 20 6 6 vss
rlabel metal1 25 25 25 25 6 zn
rlabel metal1 28 36 28 36 6 b
rlabel metal1 20 44 20 44 6 a
rlabel metal1 28 52 28 52 6 a
rlabel metal1 20 74 20 74 6 vdd
rlabel metal1 36 40 36 40 6 b
rlabel metal1 28 60 28 60 6 zn
<< end >>
