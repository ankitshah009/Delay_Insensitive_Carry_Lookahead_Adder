magic
tech scmos
timestamp 1179385222
<< checkpaint >>
rect -22 -22 94 94
<< ab >>
rect 0 0 72 72
<< pwell >>
rect -4 -4 76 32
<< nwell >>
rect -4 32 76 76
<< polysilicon >>
rect 9 60 11 65
rect 21 60 23 65
rect 61 62 63 67
rect 39 54 41 59
rect 49 54 51 59
rect 9 45 11 48
rect 9 44 15 45
rect 9 40 10 44
rect 14 40 15 44
rect 9 39 15 40
rect 9 18 11 39
rect 21 35 23 48
rect 61 43 63 46
rect 60 42 66 43
rect 60 38 61 42
rect 65 38 66 42
rect 39 35 41 38
rect 17 34 23 35
rect 17 30 18 34
rect 22 30 23 34
rect 17 29 23 30
rect 33 34 41 35
rect 33 30 34 34
rect 38 31 41 34
rect 49 35 51 38
rect 60 37 66 38
rect 49 34 55 35
rect 38 30 45 31
rect 33 29 45 30
rect 49 30 50 34
rect 54 30 55 34
rect 49 29 55 30
rect 21 26 23 29
rect 43 26 45 29
rect 53 26 55 29
rect 60 26 62 37
rect 21 15 23 20
rect 9 7 11 12
rect 43 15 45 20
rect 53 14 55 19
rect 60 14 62 19
<< ndiffusion >>
rect 13 20 21 26
rect 23 25 30 26
rect 23 21 25 25
rect 29 21 30 25
rect 23 20 30 21
rect 34 20 43 26
rect 45 25 53 26
rect 45 21 47 25
rect 51 21 53 25
rect 45 20 53 21
rect 13 18 19 20
rect 2 17 9 18
rect 2 13 3 17
rect 7 13 9 17
rect 2 12 9 13
rect 11 12 19 18
rect 13 8 19 12
rect 13 4 14 8
rect 18 4 19 8
rect 13 3 19 4
rect 34 8 41 20
rect 48 19 53 20
rect 55 19 60 26
rect 62 24 69 26
rect 62 20 64 24
rect 68 20 69 24
rect 62 19 69 20
rect 34 4 36 8
rect 40 4 41 8
rect 34 3 41 4
<< pdiffusion >>
rect 13 68 19 69
rect 13 64 14 68
rect 18 64 19 68
rect 13 60 19 64
rect 53 61 61 62
rect 4 54 9 60
rect 2 53 9 54
rect 2 49 3 53
rect 7 49 9 53
rect 2 48 9 49
rect 11 48 21 60
rect 23 54 28 60
rect 53 57 54 61
rect 58 57 61 61
rect 53 54 61 57
rect 23 53 30 54
rect 23 49 25 53
rect 29 49 30 53
rect 23 48 30 49
rect 34 44 39 54
rect 32 43 39 44
rect 32 39 33 43
rect 37 39 39 43
rect 32 38 39 39
rect 41 51 49 54
rect 41 47 43 51
rect 47 47 49 51
rect 41 38 49 47
rect 51 46 61 54
rect 63 59 68 62
rect 63 58 70 59
rect 63 54 65 58
rect 69 54 70 58
rect 63 51 70 54
rect 63 47 65 51
rect 69 47 70 51
rect 63 46 70 47
rect 51 38 58 46
<< metal1 >>
rect -2 68 74 72
rect -2 64 14 68
rect 18 64 36 68
rect 40 64 44 68
rect 48 64 74 68
rect 54 61 58 64
rect 2 53 7 54
rect 2 49 3 53
rect 2 48 7 49
rect 10 53 22 59
rect 54 56 58 57
rect 64 54 65 58
rect 69 54 70 58
rect 25 53 29 54
rect 2 17 6 48
rect 10 44 14 53
rect 64 51 70 54
rect 10 39 14 40
rect 18 35 22 43
rect 10 34 22 35
rect 10 30 18 34
rect 10 29 22 30
rect 25 34 29 49
rect 33 43 38 51
rect 42 47 43 51
rect 47 47 65 51
rect 69 47 70 51
rect 37 39 46 43
rect 33 37 46 39
rect 57 42 70 43
rect 57 38 61 42
rect 65 38 70 42
rect 25 30 34 34
rect 38 30 39 34
rect 10 21 14 29
rect 25 25 29 30
rect 42 25 46 37
rect 49 30 50 34
rect 54 30 60 34
rect 42 21 47 25
rect 51 21 52 25
rect 25 20 29 21
rect 56 17 60 30
rect 66 29 70 38
rect 2 13 3 17
rect 7 13 60 17
rect 64 24 68 25
rect 64 8 68 20
rect -2 4 14 8
rect 18 4 25 8
rect 29 4 36 8
rect 40 4 56 8
rect 60 4 64 8
rect 68 4 74 8
rect -2 0 74 4
<< ntransistor >>
rect 21 20 23 26
rect 43 20 45 26
rect 9 12 11 18
rect 53 19 55 26
rect 60 19 62 26
<< ptransistor >>
rect 9 48 11 60
rect 21 48 23 60
rect 39 38 41 54
rect 49 38 51 54
rect 61 46 63 62
<< polycontact >>
rect 10 40 14 44
rect 61 38 65 42
rect 18 30 22 34
rect 34 30 38 34
rect 50 30 54 34
<< ndcontact >>
rect 25 21 29 25
rect 47 21 51 25
rect 3 13 7 17
rect 14 4 18 8
rect 64 20 68 24
rect 36 4 40 8
<< pdcontact >>
rect 14 64 18 68
rect 3 49 7 53
rect 54 57 58 61
rect 25 49 29 53
rect 33 39 37 43
rect 43 47 47 51
rect 65 54 69 58
rect 65 47 69 51
<< psubstratepcontact >>
rect 25 4 29 8
rect 56 4 60 8
rect 64 4 68 8
<< nsubstratencontact >>
rect 36 64 40 68
rect 44 64 48 68
<< psubstratepdiff >>
rect 24 8 30 9
rect 24 4 25 8
rect 29 4 30 8
rect 24 3 30 4
rect 55 8 69 9
rect 55 4 56 8
rect 60 4 64 8
rect 68 4 69 8
rect 55 3 69 4
<< nsubstratendiff >>
rect 35 68 49 69
rect 35 64 36 68
rect 40 64 44 68
rect 48 64 49 68
rect 35 63 49 64
<< labels >>
rlabel polycontact 37 32 37 32 6 bn
rlabel polycontact 52 32 52 32 6 a2n
rlabel metal1 12 28 12 28 6 b
rlabel metal1 4 33 4 33 6 a2n
rlabel metal1 12 52 12 52 6 a2
rlabel metal1 27 37 27 37 6 bn
rlabel metal1 20 36 20 36 6 b
rlabel metal1 20 56 20 56 6 a2
rlabel metal1 36 4 36 4 6 vss
rlabel metal1 32 32 32 32 6 bn
rlabel metal1 44 32 44 32 6 z
rlabel pdcontact 36 40 36 40 6 z
rlabel metal1 36 68 36 68 6 vdd
rlabel metal1 31 15 31 15 6 a2n
rlabel metal1 54 32 54 32 6 a2n
rlabel metal1 60 40 60 40 6 a1
rlabel metal1 68 36 68 36 6 a1
rlabel metal1 56 49 56 49 6 n1
rlabel metal1 67 52 67 52 6 n1
<< end >>
