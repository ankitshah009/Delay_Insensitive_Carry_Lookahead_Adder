magic
tech scmos
timestamp 1179387803
<< checkpaint >>
rect -22 -25 142 105
<< ab >>
rect 0 0 120 80
<< pwell >>
rect -4 -7 124 36
<< nwell >>
rect -4 36 124 87
<< polysilicon >>
rect 17 67 19 72
rect 29 67 31 72
rect 39 67 41 72
rect 49 67 51 72
rect 77 70 79 74
rect 2 54 8 55
rect 2 50 3 54
rect 7 50 8 54
rect 2 49 8 50
rect 6 45 8 49
rect 89 65 91 70
rect 99 65 101 70
rect 109 65 111 70
rect 77 51 79 54
rect 65 50 79 51
rect 17 45 19 48
rect 6 43 19 45
rect 9 25 11 43
rect 29 38 31 48
rect 39 39 41 48
rect 49 45 51 48
rect 65 46 66 50
rect 70 49 79 50
rect 70 46 71 49
rect 65 45 71 46
rect 45 44 51 45
rect 45 40 46 44
rect 50 40 51 44
rect 89 41 91 49
rect 45 39 51 40
rect 55 40 91 41
rect 99 40 101 49
rect 17 37 31 38
rect 17 33 18 37
rect 22 36 31 37
rect 35 38 41 39
rect 22 33 23 36
rect 35 34 36 38
rect 40 34 41 38
rect 35 33 41 34
rect 17 32 23 33
rect 20 25 22 32
rect 39 31 41 33
rect 30 25 32 29
rect 39 28 42 31
rect 40 25 42 28
rect 47 25 49 39
rect 55 36 56 40
rect 60 39 91 40
rect 95 39 101 40
rect 109 39 111 49
rect 60 36 61 39
rect 55 35 61 36
rect 65 34 71 35
rect 65 30 66 34
rect 70 30 71 34
rect 65 29 71 30
rect 69 26 71 29
rect 81 23 83 39
rect 95 35 96 39
rect 100 35 101 39
rect 95 34 101 35
rect 99 29 101 34
rect 105 38 111 39
rect 105 34 106 38
rect 110 34 111 38
rect 105 33 111 34
rect 91 23 93 28
rect 99 26 103 29
rect 101 23 103 26
rect 108 23 110 33
rect 9 8 11 16
rect 20 12 22 16
rect 30 8 32 16
rect 40 11 42 16
rect 47 11 49 16
rect 9 6 32 8
rect 69 8 71 19
rect 81 12 83 16
rect 91 8 93 16
rect 101 11 103 16
rect 108 11 110 16
rect 69 6 93 8
<< ndiffusion >>
rect 62 25 69 26
rect 2 24 9 25
rect 2 20 3 24
rect 7 20 9 24
rect 2 19 9 20
rect 4 16 9 19
rect 11 21 20 25
rect 11 17 14 21
rect 18 17 20 21
rect 11 16 20 17
rect 22 21 30 25
rect 22 17 24 21
rect 28 17 30 21
rect 22 16 30 17
rect 32 22 40 25
rect 32 18 34 22
rect 38 18 40 22
rect 32 16 40 18
rect 42 16 47 25
rect 49 16 57 25
rect 62 21 63 25
rect 67 21 69 25
rect 62 19 69 21
rect 71 23 79 26
rect 71 19 81 23
rect 51 15 57 16
rect 51 11 52 15
rect 56 11 57 15
rect 51 10 57 11
rect 73 17 81 19
rect 73 13 74 17
rect 78 16 81 17
rect 83 22 91 23
rect 83 18 85 22
rect 89 18 91 22
rect 83 16 91 18
rect 93 22 101 23
rect 93 18 95 22
rect 99 18 101 22
rect 93 16 101 18
rect 103 16 108 23
rect 110 16 118 23
rect 78 13 79 16
rect 73 12 79 13
rect 112 12 118 16
rect 112 8 113 12
rect 117 8 118 12
rect 112 7 118 8
<< pdiffusion >>
rect 21 72 27 73
rect 21 68 22 72
rect 26 68 27 72
rect 21 67 27 68
rect 81 72 87 73
rect 81 70 82 72
rect 12 54 17 67
rect 10 53 17 54
rect 10 49 11 53
rect 15 49 17 53
rect 10 48 17 49
rect 19 48 29 67
rect 31 53 39 67
rect 31 49 33 53
rect 37 49 39 53
rect 31 48 39 49
rect 41 54 49 67
rect 41 50 43 54
rect 47 50 49 54
rect 41 48 49 50
rect 51 63 56 67
rect 72 64 77 70
rect 70 63 77 64
rect 51 62 58 63
rect 51 58 53 62
rect 57 58 58 62
rect 70 59 71 63
rect 75 59 77 63
rect 70 58 77 59
rect 51 57 58 58
rect 51 48 56 57
rect 72 54 77 58
rect 79 68 82 70
rect 86 68 87 72
rect 79 65 87 68
rect 79 54 89 65
rect 81 49 89 54
rect 91 54 99 65
rect 91 50 93 54
rect 97 50 99 54
rect 91 49 99 50
rect 101 55 109 65
rect 101 51 103 55
rect 107 51 109 55
rect 101 49 109 51
rect 111 63 118 65
rect 111 59 113 63
rect 117 59 118 63
rect 111 58 118 59
rect 111 49 116 58
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect 118 78 122 82
rect -2 72 122 78
rect -2 68 22 72
rect 26 68 82 72
rect 86 68 122 72
rect 2 58 15 63
rect 26 58 53 62
rect 57 58 58 62
rect 70 59 71 63
rect 75 59 113 63
rect 117 59 118 63
rect 2 54 7 58
rect 26 54 30 58
rect 2 50 3 54
rect 2 49 7 50
rect 11 53 30 54
rect 15 50 30 53
rect 11 43 15 49
rect 3 39 15 43
rect 3 24 7 39
rect 18 37 22 39
rect 26 38 30 50
rect 33 53 37 54
rect 42 50 43 54
rect 47 50 58 54
rect 33 46 37 49
rect 33 44 50 46
rect 33 42 46 44
rect 26 34 36 38
rect 40 34 41 38
rect 18 31 22 33
rect 10 25 22 31
rect 46 30 50 40
rect 26 26 50 30
rect 54 40 58 50
rect 66 50 70 55
rect 66 42 79 46
rect 54 36 56 40
rect 60 36 61 40
rect 26 21 30 26
rect 54 22 58 36
rect 66 34 70 42
rect 84 39 88 59
rect 93 54 97 55
rect 102 51 103 55
rect 107 51 118 55
rect 93 47 97 50
rect 93 43 110 47
rect 66 29 70 30
rect 76 35 96 39
rect 100 35 101 39
rect 106 38 110 43
rect 76 25 80 35
rect 106 31 110 34
rect 3 19 7 20
rect 13 17 14 21
rect 18 17 19 21
rect 23 17 24 21
rect 28 17 30 21
rect 33 18 34 22
rect 38 18 58 22
rect 62 21 63 25
rect 67 21 80 25
rect 85 27 110 31
rect 85 22 89 27
rect 114 22 118 51
rect 94 18 95 22
rect 99 18 118 22
rect 85 17 89 18
rect 13 12 19 17
rect 51 12 52 15
rect -2 11 52 12
rect 56 12 57 15
rect 73 13 74 17
rect 78 13 79 17
rect 73 12 79 13
rect 56 11 113 12
rect -2 8 113 11
rect 117 8 122 12
rect -2 2 122 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 122 2
<< ntransistor >>
rect 9 16 11 25
rect 20 16 22 25
rect 30 16 32 25
rect 40 16 42 25
rect 47 16 49 25
rect 69 19 71 26
rect 81 16 83 23
rect 91 16 93 23
rect 101 16 103 23
rect 108 16 110 23
<< ptransistor >>
rect 17 48 19 67
rect 29 48 31 67
rect 39 48 41 67
rect 49 48 51 67
rect 77 54 79 70
rect 89 49 91 65
rect 99 49 101 65
rect 109 49 111 65
<< polycontact >>
rect 3 50 7 54
rect 66 46 70 50
rect 46 40 50 44
rect 18 33 22 37
rect 36 34 40 38
rect 56 36 60 40
rect 66 30 70 34
rect 96 35 100 39
rect 106 34 110 38
<< ndcontact >>
rect 3 20 7 24
rect 14 17 18 21
rect 24 17 28 21
rect 34 18 38 22
rect 63 21 67 25
rect 52 11 56 15
rect 74 13 78 17
rect 85 18 89 22
rect 95 18 99 22
rect 113 8 117 12
<< pdcontact >>
rect 22 68 26 72
rect 11 49 15 53
rect 33 49 37 53
rect 43 50 47 54
rect 53 58 57 62
rect 71 59 75 63
rect 82 68 86 72
rect 93 50 97 54
rect 103 51 107 55
rect 113 59 117 63
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
rect 90 -2 94 2
rect 98 -2 102 2
rect 106 -2 110 2
rect 114 -2 118 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
rect 90 78 94 82
rect 98 78 102 82
rect 106 78 110 82
rect 114 78 118 82
<< psubstratepdiff >>
rect 0 2 120 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 120 2
rect 0 -3 120 -2
<< nsubstratendiff >>
rect 0 82 120 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect 118 78 120 82
rect 0 77 120 78
<< labels >>
rlabel polycontact 38 36 38 36 6 bn
rlabel polycontact 48 42 48 42 6 an
rlabel polycontact 58 38 58 38 6 iz
rlabel polysilicon 109 25 109 25 6 zn
rlabel polycontact 98 37 98 37 6 cn
rlabel metal1 12 28 12 28 6 a
rlabel metal1 5 31 5 31 6 bn
rlabel metal1 13 46 13 46 6 bn
rlabel metal1 4 56 4 56 6 b
rlabel metal1 12 60 12 60 6 b
rlabel ndcontact 26 19 26 19 6 an
rlabel metal1 20 32 20 32 6 a
rlabel metal1 33 36 33 36 6 bn
rlabel metal1 35 48 35 48 6 an
rlabel metal1 60 6 60 6 6 vss
rlabel metal1 45 20 45 20 6 iz
rlabel metal1 48 36 48 36 6 an
rlabel metal1 68 44 68 44 6 c
rlabel metal1 50 52 50 52 6 iz
rlabel metal1 56 36 56 36 6 iz
rlabel metal1 42 60 42 60 6 bn
rlabel metal1 60 74 60 74 6 vdd
rlabel metal1 71 23 71 23 6 cn
rlabel metal1 87 24 87 24 6 zn
rlabel metal1 76 44 76 44 6 c
rlabel metal1 100 20 100 20 6 z
rlabel metal1 108 20 108 20 6 z
rlabel polycontact 108 37 108 37 6 zn
rlabel metal1 88 37 88 37 6 cn
rlabel metal1 116 40 116 40 6 z
rlabel metal1 95 49 95 49 6 zn
rlabel metal1 94 61 94 61 6 cn
<< end >>
