magic
tech scmos
timestamp 1179387188
<< checkpaint >>
rect -22 -22 126 94
<< ab >>
rect 0 0 104 72
<< pwell >>
rect -4 -4 108 32
<< nwell >>
rect -4 32 108 76
<< polysilicon >>
rect 9 66 11 70
rect 19 66 21 70
rect 29 62 31 67
rect 39 62 41 67
rect 49 62 51 67
rect 56 62 58 67
rect 66 62 68 67
rect 73 62 75 67
rect 83 56 85 61
rect 90 56 92 61
rect 9 35 11 38
rect 19 35 21 38
rect 29 35 31 38
rect 39 35 41 38
rect 49 35 51 38
rect 9 34 41 35
rect 9 33 32 34
rect 9 26 11 33
rect 19 26 21 33
rect 29 30 32 33
rect 36 33 41 34
rect 45 34 51 35
rect 36 30 37 33
rect 29 29 37 30
rect 45 30 46 34
rect 50 30 51 34
rect 45 29 51 30
rect 56 35 58 38
rect 66 35 68 38
rect 56 34 68 35
rect 56 30 63 34
rect 67 30 68 34
rect 56 29 68 30
rect 73 35 75 38
rect 83 35 85 38
rect 90 35 92 38
rect 73 33 85 35
rect 89 34 95 35
rect 29 26 31 29
rect 9 9 11 14
rect 46 24 48 29
rect 56 24 58 29
rect 73 27 75 33
rect 89 30 90 34
rect 94 30 95 34
rect 89 29 95 30
rect 72 26 78 27
rect 72 22 73 26
rect 77 22 78 26
rect 72 21 78 22
rect 19 2 21 6
rect 29 2 31 6
rect 46 2 48 6
rect 56 2 58 6
<< ndiffusion >>
rect 2 25 9 26
rect 2 21 3 25
rect 7 21 9 25
rect 2 20 9 21
rect 4 14 9 20
rect 11 19 19 26
rect 11 15 13 19
rect 17 15 19 19
rect 11 14 19 15
rect 13 6 19 14
rect 21 25 29 26
rect 21 21 23 25
rect 27 21 29 25
rect 21 18 29 21
rect 21 14 23 18
rect 27 14 29 18
rect 21 6 29 14
rect 31 24 44 26
rect 31 12 46 24
rect 31 8 33 12
rect 37 8 46 12
rect 31 6 46 8
rect 48 17 56 24
rect 48 13 50 17
rect 54 13 56 17
rect 48 6 56 13
rect 58 18 65 24
rect 58 14 60 18
rect 64 14 65 18
rect 58 11 65 14
rect 58 7 60 11
rect 64 7 65 11
rect 58 6 65 7
<< pdiffusion >>
rect 2 65 9 66
rect 2 61 3 65
rect 7 61 9 65
rect 2 58 9 61
rect 2 54 3 58
rect 7 54 9 58
rect 2 38 9 54
rect 11 58 19 66
rect 11 54 13 58
rect 17 54 19 58
rect 11 51 19 54
rect 11 47 13 51
rect 17 47 19 51
rect 11 38 19 47
rect 21 62 27 66
rect 21 61 29 62
rect 21 57 23 61
rect 27 57 29 61
rect 21 38 29 57
rect 31 58 39 62
rect 31 54 33 58
rect 37 54 39 58
rect 31 51 39 54
rect 31 47 33 51
rect 37 47 39 51
rect 31 38 39 47
rect 41 61 49 62
rect 41 57 43 61
rect 47 57 49 61
rect 41 53 49 57
rect 41 49 43 53
rect 47 49 49 53
rect 41 38 49 49
rect 51 38 56 62
rect 58 52 66 62
rect 58 48 60 52
rect 64 48 66 52
rect 58 44 66 48
rect 58 40 60 44
rect 64 40 66 44
rect 58 38 66 40
rect 68 38 73 62
rect 75 56 81 62
rect 75 55 83 56
rect 75 51 77 55
rect 81 51 83 55
rect 75 38 83 51
rect 85 38 90 56
rect 92 51 97 56
rect 92 50 99 51
rect 92 46 94 50
rect 98 46 99 50
rect 92 43 99 46
rect 92 39 94 43
rect 98 39 99 43
rect 92 38 99 39
<< metal1 >>
rect -2 68 106 72
rect -2 65 86 68
rect -2 64 3 65
rect 2 61 3 64
rect 7 64 86 65
rect 90 64 94 68
rect 98 64 106 68
rect 7 61 8 64
rect 2 58 8 61
rect 23 61 27 64
rect 2 54 3 58
rect 7 54 8 58
rect 13 58 17 59
rect 43 61 47 64
rect 23 56 27 57
rect 33 58 39 59
rect 13 51 17 54
rect 9 47 13 50
rect 37 54 39 58
rect 33 51 39 54
rect 17 47 33 50
rect 37 47 39 51
rect 43 53 47 57
rect 77 55 81 64
rect 43 48 47 49
rect 60 52 64 53
rect 77 50 81 51
rect 94 50 98 51
rect 9 46 39 47
rect 18 35 22 46
rect 60 44 64 48
rect 2 34 22 35
rect 37 40 60 42
rect 94 43 98 46
rect 64 40 94 42
rect 37 39 94 40
rect 37 38 98 39
rect 37 34 41 38
rect 2 30 27 34
rect 31 30 32 34
rect 36 30 41 34
rect 45 30 46 34
rect 50 30 55 34
rect 62 30 63 34
rect 67 30 90 34
rect 94 30 95 34
rect 2 25 7 30
rect 2 21 3 25
rect 2 20 7 21
rect 23 25 27 30
rect 13 19 17 20
rect 13 8 17 15
rect 23 18 27 21
rect 37 22 41 30
rect 49 26 55 30
rect 49 22 73 26
rect 77 22 78 26
rect 89 22 95 30
rect 37 18 45 22
rect 23 13 27 14
rect 41 17 45 18
rect 41 13 50 17
rect 54 13 55 17
rect 59 14 60 18
rect 64 14 65 18
rect 33 12 37 13
rect 59 11 65 14
rect 74 13 78 22
rect 59 8 60 11
rect -2 7 60 8
rect 64 8 65 11
rect 64 7 86 8
rect -2 4 86 7
rect 90 4 94 8
rect 98 4 106 8
rect -2 0 106 4
<< ntransistor >>
rect 9 14 11 26
rect 19 6 21 26
rect 29 6 31 26
rect 46 6 48 24
rect 56 6 58 24
<< ptransistor >>
rect 9 38 11 66
rect 19 38 21 66
rect 29 38 31 62
rect 39 38 41 62
rect 49 38 51 62
rect 56 38 58 62
rect 66 38 68 62
rect 73 38 75 62
rect 83 38 85 56
rect 90 38 92 56
<< polycontact >>
rect 32 30 36 34
rect 46 30 50 34
rect 63 30 67 34
rect 90 30 94 34
rect 73 22 77 26
<< ndcontact >>
rect 3 21 7 25
rect 13 15 17 19
rect 23 21 27 25
rect 23 14 27 18
rect 33 8 37 12
rect 50 13 54 17
rect 60 14 64 18
rect 60 7 64 11
<< pdcontact >>
rect 3 61 7 65
rect 3 54 7 58
rect 13 54 17 58
rect 13 47 17 51
rect 23 57 27 61
rect 33 54 37 58
rect 33 47 37 51
rect 43 57 47 61
rect 43 49 47 53
rect 60 48 64 52
rect 60 40 64 44
rect 77 51 81 55
rect 94 46 98 50
rect 94 39 98 43
<< psubstratepcontact >>
rect 86 4 90 8
rect 94 4 98 8
<< nsubstratencontact >>
rect 86 64 90 68
rect 94 64 98 68
<< psubstratepdiff >>
rect 85 8 99 24
rect 85 4 86 8
rect 90 4 94 8
rect 98 4 99 8
rect 85 3 99 4
<< nsubstratendiff >>
rect 85 68 99 69
rect 85 64 86 68
rect 90 64 94 68
rect 98 64 99 68
rect 85 63 99 64
<< labels >>
rlabel polycontact 33 32 33 32 6 zn
rlabel metal1 12 32 12 32 6 z
rlabel metal1 4 28 4 28 6 z
rlabel metal1 12 48 12 48 6 z
rlabel metal1 20 40 20 40 6 z
rlabel metal1 36 52 36 52 6 z
rlabel metal1 28 48 28 48 6 z
rlabel metal1 52 4 52 4 6 vss
rlabel metal1 48 15 48 15 6 zn
rlabel metal1 60 24 60 24 6 a
rlabel metal1 52 28 52 28 6 a
rlabel metal1 36 32 36 32 6 zn
rlabel metal1 52 68 52 68 6 vdd
rlabel metal1 76 16 76 16 6 a
rlabel metal1 68 24 68 24 6 a
rlabel metal1 68 32 68 32 6 b
rlabel metal1 76 32 76 32 6 b
rlabel metal1 62 45 62 45 6 zn
rlabel metal1 92 28 92 28 6 b
rlabel metal1 84 32 84 32 6 b
rlabel metal1 96 44 96 44 6 zn
<< end >>
