magic
tech scmos
timestamp 1185038962
<< checkpaint >>
rect -22 -24 202 124
<< ab >>
rect 0 0 180 100
<< pwell >>
rect -2 -4 182 49
<< nwell >>
rect -2 49 182 104
<< polysilicon >>
rect 11 95 13 98
rect 23 95 25 98
rect 35 83 37 86
rect 47 83 49 86
rect 83 77 85 80
rect 95 77 97 80
rect 107 77 109 80
rect 119 77 121 80
rect 155 95 157 98
rect 167 95 169 98
rect 131 77 133 80
rect 71 71 73 74
rect 11 43 13 55
rect 23 43 25 55
rect 35 53 37 65
rect 47 63 49 65
rect 47 62 53 63
rect 47 58 48 62
rect 52 58 53 62
rect 47 57 53 58
rect 29 52 37 53
rect 29 48 30 52
rect 34 48 37 52
rect 71 53 73 55
rect 83 53 85 55
rect 71 52 85 53
rect 71 51 78 52
rect 29 47 37 48
rect 77 48 78 51
rect 82 51 85 52
rect 95 53 97 55
rect 95 52 103 53
rect 95 51 98 52
rect 82 48 83 51
rect 77 47 83 48
rect 97 48 98 51
rect 102 48 103 52
rect 97 47 103 48
rect 11 41 25 43
rect 37 42 43 43
rect 37 41 38 42
rect 11 39 38 41
rect 11 37 25 39
rect 37 38 38 39
rect 42 38 43 42
rect 37 37 43 38
rect 47 42 53 43
rect 47 38 48 42
rect 52 38 53 42
rect 47 37 53 38
rect 63 42 69 43
rect 63 38 64 42
rect 68 41 69 42
rect 107 41 109 55
rect 119 43 121 55
rect 131 53 133 55
rect 127 52 133 53
rect 127 48 128 52
rect 132 48 133 52
rect 127 47 133 48
rect 155 43 157 55
rect 167 43 169 55
rect 68 39 109 41
rect 68 38 69 39
rect 63 37 69 38
rect 11 25 13 37
rect 23 25 25 37
rect 29 32 37 33
rect 29 28 30 32
rect 34 28 37 32
rect 47 29 49 37
rect 97 34 103 35
rect 77 32 83 33
rect 77 29 78 32
rect 29 27 37 28
rect 35 25 37 27
rect 71 28 78 29
rect 82 29 83 32
rect 97 31 98 34
rect 95 30 98 31
rect 102 30 103 34
rect 95 29 103 30
rect 82 28 85 29
rect 71 27 85 28
rect 95 27 97 29
rect 107 27 109 39
rect 117 42 123 43
rect 117 38 118 42
rect 122 41 123 42
rect 137 42 143 43
rect 137 41 138 42
rect 122 39 138 41
rect 122 38 123 39
rect 117 37 123 38
rect 137 38 138 39
rect 142 38 143 42
rect 137 37 143 38
rect 147 42 169 43
rect 147 38 148 42
rect 152 38 169 42
rect 147 37 169 38
rect 127 32 133 33
rect 127 29 128 32
rect 119 28 128 29
rect 132 28 133 32
rect 119 27 133 28
rect 71 25 73 27
rect 83 25 85 27
rect 35 12 37 15
rect 47 12 49 15
rect 71 14 73 17
rect 119 25 121 27
rect 131 25 133 27
rect 155 25 157 37
rect 167 25 169 37
rect 83 12 85 15
rect 95 12 97 15
rect 107 12 109 15
rect 119 12 121 15
rect 131 14 133 17
rect 11 2 13 5
rect 23 2 25 5
rect 155 2 157 5
rect 167 2 169 5
<< ndiffusion >>
rect 39 25 47 29
rect 3 22 11 25
rect 3 18 4 22
rect 8 18 11 22
rect 3 12 11 18
rect 3 8 4 12
rect 8 8 11 12
rect 3 5 11 8
rect 13 22 23 25
rect 13 18 16 22
rect 20 18 23 22
rect 13 5 23 18
rect 25 15 35 25
rect 37 15 47 25
rect 49 22 57 29
rect 87 25 95 27
rect 49 18 52 22
rect 56 18 57 22
rect 49 15 57 18
rect 63 22 71 25
rect 63 18 64 22
rect 68 18 71 22
rect 63 17 71 18
rect 73 17 83 25
rect 25 12 33 15
rect 75 15 83 17
rect 85 15 95 25
rect 97 24 107 27
rect 97 20 100 24
rect 104 20 107 24
rect 97 15 107 20
rect 109 25 117 27
rect 135 32 143 33
rect 135 28 138 32
rect 142 28 143 32
rect 135 27 143 28
rect 135 25 141 27
rect 109 15 119 25
rect 121 17 131 25
rect 133 17 141 25
rect 151 21 155 25
rect 121 15 129 17
rect 75 12 81 15
rect 123 12 129 15
rect 25 8 28 12
rect 32 8 33 12
rect 25 5 33 8
rect 75 8 76 12
rect 80 8 81 12
rect 75 7 81 8
rect 123 8 124 12
rect 128 8 129 12
rect 123 7 129 8
rect 147 12 155 21
rect 147 8 148 12
rect 152 8 155 12
rect 147 5 155 8
rect 157 22 167 25
rect 157 18 160 22
rect 164 18 167 22
rect 157 5 167 18
rect 169 22 177 25
rect 169 18 172 22
rect 176 18 177 22
rect 169 12 177 18
rect 169 8 172 12
rect 176 8 177 12
rect 169 5 177 8
<< pdiffusion >>
rect 3 92 11 95
rect 3 88 4 92
rect 8 88 11 92
rect 3 82 11 88
rect 3 78 4 82
rect 8 78 11 82
rect 3 72 11 78
rect 3 68 4 72
rect 8 68 11 72
rect 3 62 11 68
rect 3 58 4 62
rect 8 58 11 62
rect 3 55 11 58
rect 13 82 23 95
rect 13 78 16 82
rect 20 78 23 82
rect 13 72 23 78
rect 13 68 16 72
rect 20 68 23 72
rect 13 62 23 68
rect 13 58 16 62
rect 20 58 23 62
rect 13 55 23 58
rect 25 92 33 95
rect 25 88 28 92
rect 32 88 33 92
rect 25 83 33 88
rect 51 92 57 93
rect 51 88 52 92
rect 56 88 57 92
rect 51 83 57 88
rect 75 92 81 93
rect 75 88 76 92
rect 80 88 81 92
rect 123 92 129 93
rect 25 65 35 83
rect 37 72 47 83
rect 37 68 40 72
rect 44 68 47 72
rect 37 65 47 68
rect 49 65 57 83
rect 75 77 81 88
rect 123 88 124 92
rect 128 88 129 92
rect 123 77 129 88
rect 147 92 155 95
rect 147 88 148 92
rect 152 88 155 92
rect 147 82 155 88
rect 147 78 148 82
rect 152 78 155 82
rect 75 71 83 77
rect 25 55 33 65
rect 63 62 71 71
rect 63 58 64 62
rect 68 58 71 62
rect 63 55 71 58
rect 73 55 83 71
rect 85 72 95 77
rect 85 68 88 72
rect 92 68 95 72
rect 85 55 95 68
rect 97 62 107 77
rect 97 58 100 62
rect 104 58 107 62
rect 97 55 107 58
rect 109 72 119 77
rect 109 68 112 72
rect 116 68 119 72
rect 109 62 119 68
rect 109 58 112 62
rect 116 58 119 62
rect 109 55 119 58
rect 121 55 131 77
rect 133 61 141 77
rect 147 72 155 78
rect 147 68 148 72
rect 152 68 155 72
rect 147 67 155 68
rect 133 60 143 61
rect 133 56 138 60
rect 142 56 143 60
rect 133 55 143 56
rect 151 55 155 67
rect 157 82 167 95
rect 157 78 160 82
rect 164 78 167 82
rect 157 72 167 78
rect 157 68 160 72
rect 164 68 167 72
rect 157 62 167 68
rect 157 58 160 62
rect 164 58 167 62
rect 157 55 167 58
rect 169 92 177 95
rect 169 88 172 92
rect 176 88 177 92
rect 169 82 177 88
rect 169 78 172 82
rect 176 78 177 82
rect 169 72 177 78
rect 169 68 172 72
rect 176 68 177 72
rect 169 62 177 68
rect 169 58 172 62
rect 176 58 177 62
rect 169 55 177 58
<< metal1 >>
rect -2 96 182 101
rect -2 92 64 96
rect 68 92 88 96
rect 92 92 100 96
rect 104 92 112 96
rect 116 92 136 96
rect 140 92 182 96
rect -2 88 4 92
rect 8 88 28 92
rect 32 88 52 92
rect 56 88 76 92
rect 80 88 124 92
rect 128 88 148 92
rect 152 88 172 92
rect 176 88 182 92
rect -2 87 182 88
rect 3 82 9 87
rect 3 78 4 82
rect 8 78 9 82
rect 3 72 9 78
rect 15 82 21 83
rect 147 82 153 87
rect 159 82 165 83
rect 15 78 16 82
rect 20 78 23 82
rect 15 77 23 78
rect 17 73 23 77
rect 3 68 4 72
rect 8 68 9 72
rect 3 62 9 68
rect 15 72 23 73
rect 15 68 16 72
rect 20 68 23 72
rect 15 67 23 68
rect 17 63 23 67
rect 3 58 4 62
rect 8 58 9 62
rect 3 57 9 58
rect 15 62 23 63
rect 15 58 16 62
rect 20 58 23 62
rect 15 57 23 58
rect 17 23 23 57
rect 3 22 9 23
rect 3 18 4 22
rect 8 18 9 22
rect 3 13 9 18
rect 15 22 23 23
rect 15 18 16 22
rect 20 18 23 22
rect 27 78 132 82
rect 27 53 33 78
rect 39 72 45 73
rect 87 72 93 73
rect 111 72 117 73
rect 39 68 40 72
rect 44 68 45 72
rect 39 67 45 68
rect 50 68 83 72
rect 27 52 35 53
rect 27 48 30 52
rect 34 48 35 52
rect 27 47 35 48
rect 27 33 33 47
rect 39 43 43 67
rect 50 63 54 68
rect 47 62 54 63
rect 47 58 48 62
rect 52 58 54 62
rect 63 62 69 63
rect 63 58 64 62
rect 68 58 69 62
rect 47 57 53 58
rect 63 57 69 58
rect 48 43 52 57
rect 64 43 68 57
rect 77 52 83 68
rect 87 68 88 72
rect 92 68 112 72
rect 116 68 117 72
rect 87 67 93 68
rect 111 67 117 68
rect 112 63 116 67
rect 99 62 105 63
rect 77 48 78 52
rect 82 48 83 52
rect 37 42 43 43
rect 37 38 38 42
rect 42 38 43 42
rect 37 37 43 38
rect 47 42 53 43
rect 47 38 48 42
rect 52 38 53 42
rect 47 37 53 38
rect 63 42 69 43
rect 63 38 64 42
rect 68 38 69 42
rect 63 37 69 38
rect 27 32 35 33
rect 27 28 30 32
rect 34 28 35 32
rect 27 27 35 28
rect 27 18 33 27
rect 39 22 43 37
rect 64 23 68 37
rect 77 32 83 48
rect 77 28 78 32
rect 82 28 83 32
rect 51 22 57 23
rect 39 18 52 22
rect 56 18 57 22
rect 15 17 21 18
rect 51 17 57 18
rect 63 22 69 23
rect 63 18 64 22
rect 68 18 69 22
rect 77 18 83 28
rect 88 58 100 62
rect 104 58 105 62
rect 88 22 92 58
rect 99 57 105 58
rect 111 62 117 63
rect 111 58 112 62
rect 116 58 117 62
rect 111 57 117 58
rect 128 53 132 78
rect 147 78 148 82
rect 152 78 153 82
rect 147 72 153 78
rect 147 68 148 72
rect 152 68 153 72
rect 147 67 153 68
rect 157 78 160 82
rect 164 78 165 82
rect 157 77 165 78
rect 171 82 177 87
rect 171 78 172 82
rect 176 78 177 82
rect 157 73 163 77
rect 157 72 165 73
rect 157 68 160 72
rect 164 68 165 72
rect 157 67 165 68
rect 171 72 177 78
rect 171 68 172 72
rect 176 68 177 72
rect 157 63 163 67
rect 157 62 165 63
rect 137 60 143 61
rect 137 56 138 60
rect 142 56 143 60
rect 137 55 143 56
rect 157 58 160 62
rect 164 58 165 62
rect 157 57 165 58
rect 171 62 177 68
rect 171 58 172 62
rect 176 58 177 62
rect 171 57 177 58
rect 97 52 103 53
rect 127 52 133 53
rect 97 48 98 52
rect 102 48 128 52
rect 132 48 133 52
rect 97 47 103 48
rect 127 47 133 48
rect 117 42 123 43
rect 108 38 118 42
rect 122 38 123 42
rect 97 34 103 35
rect 108 34 112 38
rect 117 37 123 38
rect 97 30 98 34
rect 102 30 112 34
rect 128 33 132 47
rect 138 43 142 55
rect 137 42 143 43
rect 137 38 138 42
rect 142 38 143 42
rect 137 37 143 38
rect 147 42 153 43
rect 147 38 148 42
rect 152 38 153 42
rect 147 37 153 38
rect 138 33 142 37
rect 127 32 133 33
rect 97 29 103 30
rect 127 28 128 32
rect 132 28 133 32
rect 127 27 133 28
rect 137 32 143 33
rect 137 28 138 32
rect 142 28 143 32
rect 137 27 143 28
rect 99 24 105 25
rect 99 22 100 24
rect 88 20 100 22
rect 104 22 105 24
rect 148 22 152 37
rect 104 20 152 22
rect 88 18 152 20
rect 157 23 163 57
rect 157 22 165 23
rect 157 18 160 22
rect 164 18 165 22
rect 63 17 69 18
rect 159 17 165 18
rect 171 22 177 23
rect 171 18 172 22
rect 176 18 177 22
rect 171 13 177 18
rect -2 12 182 13
rect -2 8 4 12
rect 8 8 28 12
rect 32 8 76 12
rect 80 8 124 12
rect 128 8 148 12
rect 152 8 172 12
rect 176 8 182 12
rect -2 4 40 8
rect 44 4 52 8
rect 56 4 64 8
rect 68 4 88 8
rect 92 4 100 8
rect 104 4 112 8
rect 116 4 182 8
rect -2 -1 182 4
<< ntransistor >>
rect 11 5 13 25
rect 23 5 25 25
rect 35 15 37 25
rect 47 15 49 29
rect 71 17 73 25
rect 83 15 85 25
rect 95 15 97 27
rect 107 15 109 27
rect 119 15 121 25
rect 131 17 133 25
rect 155 5 157 25
rect 167 5 169 25
<< ptransistor >>
rect 11 55 13 95
rect 23 55 25 95
rect 35 65 37 83
rect 47 65 49 83
rect 71 55 73 71
rect 83 55 85 77
rect 95 55 97 77
rect 107 55 109 77
rect 119 55 121 77
rect 131 55 133 77
rect 155 55 157 95
rect 167 55 169 95
<< polycontact >>
rect 48 58 52 62
rect 30 48 34 52
rect 78 48 82 52
rect 98 48 102 52
rect 38 38 42 42
rect 48 38 52 42
rect 64 38 68 42
rect 128 48 132 52
rect 30 28 34 32
rect 78 28 82 32
rect 98 30 102 34
rect 118 38 122 42
rect 138 38 142 42
rect 148 38 152 42
rect 128 28 132 32
<< ndcontact >>
rect 4 18 8 22
rect 4 8 8 12
rect 16 18 20 22
rect 52 18 56 22
rect 64 18 68 22
rect 100 20 104 24
rect 138 28 142 32
rect 28 8 32 12
rect 76 8 80 12
rect 124 8 128 12
rect 148 8 152 12
rect 160 18 164 22
rect 172 18 176 22
rect 172 8 176 12
<< pdcontact >>
rect 4 88 8 92
rect 4 78 8 82
rect 4 68 8 72
rect 4 58 8 62
rect 16 78 20 82
rect 16 68 20 72
rect 16 58 20 62
rect 28 88 32 92
rect 52 88 56 92
rect 76 88 80 92
rect 40 68 44 72
rect 124 88 128 92
rect 148 88 152 92
rect 148 78 152 82
rect 64 58 68 62
rect 88 68 92 72
rect 100 58 104 62
rect 112 68 116 72
rect 112 58 116 62
rect 148 68 152 72
rect 138 56 142 60
rect 160 78 164 82
rect 160 68 164 72
rect 160 58 164 62
rect 172 88 176 92
rect 172 78 176 82
rect 172 68 176 72
rect 172 58 176 62
<< psubstratepcontact >>
rect 40 4 44 8
rect 52 4 56 8
rect 64 4 68 8
rect 88 4 92 8
rect 100 4 104 8
rect 112 4 116 8
<< nsubstratencontact >>
rect 64 92 68 96
rect 88 92 92 96
rect 100 92 104 96
rect 112 92 116 96
rect 136 92 140 96
<< psubstratepdiff >>
rect 39 8 69 9
rect 39 4 40 8
rect 44 4 52 8
rect 56 4 64 8
rect 68 4 69 8
rect 87 8 117 9
rect 39 3 69 4
rect 87 4 88 8
rect 92 4 100 8
rect 104 4 112 8
rect 116 4 117 8
rect 87 3 117 4
<< nsubstratendiff >>
rect 63 96 69 97
rect 63 92 64 96
rect 68 92 69 96
rect 87 96 117 97
rect 63 85 69 92
rect 87 92 88 96
rect 92 92 100 96
rect 104 92 112 96
rect 116 92 117 96
rect 135 96 141 97
rect 87 91 117 92
rect 135 92 136 96
rect 140 92 141 96
rect 135 85 141 92
<< labels >>
rlabel metal1 30 50 30 50 6 a
rlabel metal1 20 50 20 50 6 cout
rlabel metal1 30 50 30 50 6 a
rlabel metal1 20 50 20 50 6 cout
rlabel psubstratepcontact 90 6 90 6 6 vss
rlabel psubstratepcontact 90 6 90 6 6 vss
rlabel metal1 80 45 80 45 6 b
rlabel metal1 80 45 80 45 6 b
rlabel nsubstratencontact 90 94 90 94 6 vdd
rlabel nsubstratencontact 90 94 90 94 6 vdd
rlabel metal1 160 50 160 50 6 sout
rlabel metal1 160 50 160 50 6 sout
<< end >>
