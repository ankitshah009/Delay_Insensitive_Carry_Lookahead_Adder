magic
tech scmos
timestamp 1179386805
<< checkpaint >>
rect -22 -22 78 94
<< ab >>
rect 0 0 56 72
<< pwell >>
rect -4 -4 60 32
<< nwell >>
rect -4 32 60 76
<< polysilicon >>
rect 12 65 14 70
rect 19 65 21 70
rect 29 65 31 70
rect 36 65 38 70
rect 12 35 14 38
rect 19 35 21 38
rect 29 35 31 38
rect 36 35 38 38
rect 9 34 15 35
rect 9 30 10 34
rect 14 30 15 34
rect 9 29 15 30
rect 19 34 32 35
rect 19 30 27 34
rect 31 30 32 34
rect 19 29 32 30
rect 36 34 49 35
rect 36 30 44 34
rect 48 30 49 34
rect 36 29 49 30
rect 9 19 11 29
rect 19 19 21 29
rect 29 19 31 29
rect 39 26 41 29
rect 39 8 41 13
rect 9 2 11 6
rect 19 2 21 6
rect 29 2 31 6
<< ndiffusion >>
rect 34 19 39 26
rect 2 11 9 19
rect 2 7 3 11
rect 7 7 9 11
rect 2 6 9 7
rect 11 18 19 19
rect 11 14 13 18
rect 17 14 19 18
rect 11 6 19 14
rect 21 11 29 19
rect 21 7 23 11
rect 27 7 29 11
rect 21 6 29 7
rect 31 18 39 19
rect 31 14 33 18
rect 37 14 39 18
rect 31 13 39 14
rect 41 18 49 26
rect 41 14 43 18
rect 47 14 49 18
rect 41 13 49 14
rect 31 6 36 13
<< pdiffusion >>
rect 4 64 12 65
rect 4 60 6 64
rect 10 60 12 64
rect 4 56 12 60
rect 4 52 6 56
rect 10 52 12 56
rect 4 38 12 52
rect 14 38 19 65
rect 21 50 29 65
rect 21 46 23 50
rect 27 46 29 50
rect 21 43 29 46
rect 21 39 23 43
rect 27 39 29 43
rect 21 38 29 39
rect 31 38 36 65
rect 38 59 43 65
rect 38 58 46 59
rect 38 54 40 58
rect 44 54 46 58
rect 38 51 46 54
rect 38 47 40 51
rect 44 47 46 51
rect 38 38 46 47
<< metal1 >>
rect -2 68 58 72
rect -2 64 48 68
rect 52 64 58 68
rect 6 56 10 60
rect 6 51 10 52
rect 40 58 44 64
rect 40 51 44 54
rect 22 46 23 50
rect 27 46 31 50
rect 40 46 44 47
rect 22 43 28 46
rect 2 39 23 43
rect 27 39 28 43
rect 2 18 6 39
rect 33 38 47 42
rect 10 34 22 35
rect 33 34 39 38
rect 14 30 22 34
rect 26 30 27 34
rect 31 30 39 34
rect 43 30 44 34
rect 48 30 49 34
rect 10 29 22 30
rect 17 26 22 29
rect 43 26 49 30
rect 17 22 49 26
rect 43 18 47 19
rect 2 14 13 18
rect 17 14 33 18
rect 37 14 39 18
rect 2 8 3 11
rect -2 7 3 8
rect 7 8 8 11
rect 22 8 23 11
rect 7 7 23 8
rect 27 8 28 11
rect 43 8 47 14
rect 27 7 48 8
rect -2 4 48 7
rect 52 4 58 8
rect -2 0 58 4
<< ntransistor >>
rect 9 6 11 19
rect 19 6 21 19
rect 29 6 31 19
rect 39 13 41 26
<< ptransistor >>
rect 12 38 14 65
rect 19 38 21 65
rect 29 38 31 65
rect 36 38 38 65
<< polycontact >>
rect 10 30 14 34
rect 27 30 31 34
rect 44 30 48 34
<< ndcontact >>
rect 3 7 7 11
rect 13 14 17 18
rect 23 7 27 11
rect 33 14 37 18
rect 43 14 47 18
<< pdcontact >>
rect 6 60 10 64
rect 6 52 10 56
rect 23 46 27 50
rect 23 39 27 43
rect 40 54 44 58
rect 40 47 44 51
<< psubstratepcontact >>
rect 48 4 52 8
<< nsubstratencontact >>
rect 48 64 52 68
<< psubstratepdiff >>
rect 47 8 53 9
rect 47 4 48 8
rect 52 4 53 8
rect 47 3 53 4
<< nsubstratendiff >>
rect 47 68 53 69
rect 47 64 48 68
rect 52 64 53 68
rect 47 63 53 64
<< labels >>
rlabel metal1 4 32 4 32 6 z
rlabel metal1 20 16 20 16 6 z
rlabel metal1 12 16 12 16 6 z
rlabel metal1 20 28 20 28 6 a
rlabel metal1 28 4 28 4 6 vss
rlabel ndcontact 36 16 36 16 6 z
rlabel metal1 28 16 28 16 6 z
rlabel metal1 28 24 28 24 6 a
rlabel metal1 36 24 36 24 6 a
rlabel metal1 36 36 36 36 6 b
rlabel metal1 28 48 28 48 6 z
rlabel metal1 28 68 28 68 6 vdd
rlabel metal1 44 24 44 24 6 a
rlabel metal1 44 40 44 40 6 b
<< end >>
