.subckt nr2v0x1 a b vdd vss z
*   SPICE3 file   created from nr2v0x1.ext -      technology: scmos
m00 w1     b      z      vdd p w=28u  l=2.3636u ad=70p      pd=33u      as=166p     ps=70u
m01 vdd    a      w1     vdd p w=28u  l=2.3636u ad=252p     pd=74u      as=70p      ps=33u
m02 z      b      vss    vss n w=8u   l=2.3636u ad=40.5p    pd=20u      as=87p      ps=40u
m03 vss    a      z      vss n w=8u   l=2.3636u ad=87p      pd=40u      as=40.5p    ps=20u
C0  b      vdd    0.023f
C1  vss    z      0.155f
C2  vss    b      0.017f
C3  z      b      0.118f
C4  w1     vdd    0.005f
C5  a      vdd    0.018f
C6  vss    a      0.036f
C7  w1     b      0.007f
C8  z      a      0.043f
C9  vss    vdd    0.004f
C10 a      b      0.125f
C11 z      vdd    0.053f
C13 z      vss    0.015f
C14 a      vss    0.021f
C15 b      vss    0.019f
.ends
