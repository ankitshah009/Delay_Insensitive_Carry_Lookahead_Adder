magic
tech scmos
timestamp 1180600737
<< checkpaint >>
rect -22 -22 122 122
<< ab >>
rect 0 0 100 100
<< pwell >>
rect -4 -4 104 48
<< nwell >>
rect -4 48 104 104
<< polysilicon >>
rect 11 94 13 98
rect 23 94 25 98
rect 35 94 37 98
rect 47 94 49 98
rect 75 94 77 98
rect 87 94 89 98
rect 11 53 13 56
rect 23 53 25 56
rect 35 53 37 56
rect 47 53 49 56
rect 75 53 77 56
rect 87 53 89 56
rect 11 51 19 53
rect 23 51 29 53
rect 35 52 43 53
rect 35 51 38 52
rect 17 43 19 51
rect 27 43 29 51
rect 37 48 38 51
rect 42 48 43 52
rect 37 47 43 48
rect 47 52 53 53
rect 47 48 48 52
rect 52 48 53 52
rect 47 47 53 48
rect 75 52 81 53
rect 75 48 76 52
rect 80 48 81 52
rect 75 47 81 48
rect 17 42 23 43
rect 17 38 18 42
rect 22 38 23 42
rect 17 37 23 38
rect 27 42 33 43
rect 27 38 28 42
rect 32 38 33 42
rect 27 37 33 38
rect 17 29 19 37
rect 27 29 29 37
rect 37 29 39 47
rect 47 29 49 47
rect 15 27 19 29
rect 23 27 29 29
rect 35 27 39 29
rect 43 27 49 29
rect 15 24 17 27
rect 23 24 25 27
rect 35 24 37 27
rect 43 24 45 27
rect 79 25 81 47
rect 87 52 93 53
rect 87 48 88 52
rect 92 48 93 52
rect 87 47 93 48
rect 87 25 89 47
rect 15 2 17 6
rect 23 2 25 6
rect 35 2 37 6
rect 43 2 45 6
rect 79 2 81 6
rect 87 2 89 6
<< ndiffusion >>
rect 7 12 15 24
rect 7 8 8 12
rect 12 8 15 12
rect 7 6 15 8
rect 17 6 23 24
rect 25 22 35 24
rect 25 18 28 22
rect 32 18 35 22
rect 25 6 35 18
rect 37 6 43 24
rect 45 12 53 24
rect 71 22 79 25
rect 71 18 72 22
rect 76 18 79 22
rect 45 8 48 12
rect 52 8 53 12
rect 45 6 53 8
rect 71 6 79 18
rect 81 6 87 25
rect 89 22 97 25
rect 89 18 92 22
rect 96 18 97 22
rect 89 12 97 18
rect 89 8 92 12
rect 96 8 97 12
rect 89 6 97 8
<< pdiffusion >>
rect 3 82 11 94
rect 3 78 4 82
rect 8 78 11 82
rect 3 56 11 78
rect 13 72 23 94
rect 13 68 16 72
rect 20 68 23 72
rect 13 56 23 68
rect 25 82 35 94
rect 25 78 28 82
rect 32 78 35 82
rect 25 56 35 78
rect 37 72 47 94
rect 37 68 40 72
rect 44 68 47 72
rect 37 56 47 68
rect 49 82 57 94
rect 49 78 52 82
rect 56 78 57 82
rect 49 56 57 78
rect 67 82 75 94
rect 67 78 68 82
rect 72 78 75 82
rect 67 56 75 78
rect 77 82 87 94
rect 77 78 80 82
rect 84 78 87 82
rect 77 56 87 78
rect 89 92 97 94
rect 89 88 92 92
rect 96 88 97 92
rect 89 82 97 88
rect 89 78 92 82
rect 96 78 97 82
rect 89 72 97 78
rect 89 68 92 72
rect 96 68 97 72
rect 89 56 97 68
<< metal1 >>
rect -2 92 102 100
rect -2 88 92 92
rect 96 88 102 92
rect 68 82 72 88
rect 3 78 4 82
rect 8 78 28 82
rect 32 78 52 82
rect 56 78 57 82
rect 68 77 72 78
rect 80 82 84 83
rect 8 72 12 73
rect 8 68 16 72
rect 20 68 21 72
rect 8 22 12 68
rect 18 42 22 63
rect 18 27 22 38
rect 28 42 32 73
rect 80 72 84 78
rect 39 68 40 72
rect 44 68 84 72
rect 92 82 96 88
rect 92 72 96 78
rect 92 67 96 68
rect 28 27 32 38
rect 38 52 42 63
rect 38 27 42 48
rect 48 52 52 63
rect 78 52 82 63
rect 75 48 76 52
rect 80 48 82 52
rect 48 27 52 48
rect 78 27 82 48
rect 88 52 92 63
rect 88 27 92 48
rect 92 22 96 23
rect 8 18 28 22
rect 32 18 72 22
rect 76 18 77 22
rect 8 17 12 18
rect 92 12 96 18
rect -2 8 8 12
rect 12 8 48 12
rect 52 10 92 12
rect 52 8 60 10
rect -2 6 60 8
rect 64 8 92 10
rect 96 8 102 12
rect 64 6 102 8
rect -2 0 102 6
<< ntransistor >>
rect 15 6 17 24
rect 23 6 25 24
rect 35 6 37 24
rect 43 6 45 24
rect 79 6 81 25
rect 87 6 89 25
<< ptransistor >>
rect 11 56 13 94
rect 23 56 25 94
rect 35 56 37 94
rect 47 56 49 94
rect 75 56 77 94
rect 87 56 89 94
<< polycontact >>
rect 38 48 42 52
rect 48 48 52 52
rect 76 48 80 52
rect 18 38 22 42
rect 28 38 32 42
rect 88 48 92 52
<< ndcontact >>
rect 8 8 12 12
rect 28 18 32 22
rect 72 18 76 22
rect 48 8 52 12
rect 92 18 96 22
rect 92 8 96 12
<< pdcontact >>
rect 4 78 8 82
rect 16 68 20 72
rect 28 78 32 82
rect 40 68 44 72
rect 52 78 56 82
rect 68 78 72 82
rect 80 78 84 82
rect 92 88 96 92
rect 92 78 96 82
rect 92 68 96 72
<< psubstratepcontact >>
rect 60 6 64 10
<< psubstratepdiff >>
rect 59 10 65 16
rect 59 6 60 10
rect 64 6 65 10
rect 59 5 65 6
<< labels >>
rlabel metal1 10 45 10 45 6 nq
rlabel ndcontact 30 20 30 20 6 nq
rlabel metal1 20 20 20 20 6 nq
rlabel metal1 20 45 20 45 6 i5
rlabel metal1 30 50 30 50 6 i4
rlabel metal1 50 6 50 6 6 vss
rlabel metal1 50 20 50 20 6 nq
rlabel metal1 40 20 40 20 6 nq
rlabel metal1 40 45 40 45 6 i3
rlabel metal1 50 45 50 45 6 i2
rlabel metal1 50 94 50 94 6 vdd
rlabel metal1 70 20 70 20 6 nq
rlabel metal1 60 20 60 20 6 nq
rlabel metal1 80 45 80 45 6 i1
rlabel metal1 90 45 90 45 6 i0
<< end >>
