magic
tech scmos
timestamp 1179385415
<< checkpaint >>
rect -22 -25 78 105
<< ab >>
rect 0 0 56 80
<< pwell >>
rect -4 -7 60 36
<< nwell >>
rect -4 36 60 87
<< polysilicon >>
rect 9 69 11 74
rect 19 69 21 74
rect 31 70 33 74
rect 41 70 43 74
rect 31 47 33 50
rect 41 47 43 50
rect 31 46 37 47
rect 9 39 11 45
rect 19 39 21 45
rect 31 42 32 46
rect 36 42 37 46
rect 31 41 37 42
rect 41 46 47 47
rect 41 42 42 46
rect 46 42 47 46
rect 41 41 47 42
rect 9 38 15 39
rect 9 34 10 38
rect 14 34 15 38
rect 9 33 15 34
rect 19 38 25 39
rect 19 34 20 38
rect 24 34 25 38
rect 19 33 25 34
rect 13 30 15 33
rect 20 30 22 33
rect 32 30 34 41
rect 41 36 43 41
rect 39 33 43 36
rect 39 30 41 33
rect 13 6 15 10
rect 20 6 22 10
rect 32 8 34 13
rect 39 8 41 13
<< ndiffusion >>
rect 8 22 13 30
rect 6 21 13 22
rect 6 17 7 21
rect 11 17 13 21
rect 6 16 13 17
rect 8 10 13 16
rect 15 10 20 30
rect 22 13 32 30
rect 34 13 39 30
rect 41 22 46 30
rect 41 21 48 22
rect 41 17 43 21
rect 47 17 48 21
rect 41 16 48 17
rect 41 13 46 16
rect 22 12 30 13
rect 22 10 25 12
rect 24 8 25 10
rect 29 8 30 12
rect 24 7 30 8
<< pdiffusion >>
rect 23 69 31 70
rect 2 68 9 69
rect 2 64 3 68
rect 7 64 9 68
rect 2 61 9 64
rect 2 57 3 61
rect 7 57 9 61
rect 2 45 9 57
rect 11 62 19 69
rect 11 58 13 62
rect 17 58 19 62
rect 11 55 19 58
rect 11 51 13 55
rect 17 51 19 55
rect 11 45 19 51
rect 21 65 24 69
rect 28 65 31 69
rect 21 50 31 65
rect 33 62 41 70
rect 33 58 35 62
rect 39 58 41 62
rect 33 50 41 58
rect 43 69 50 70
rect 43 65 45 69
rect 49 65 50 69
rect 43 62 50 65
rect 43 58 45 62
rect 49 58 50 62
rect 43 50 50 58
rect 21 45 29 50
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect -2 69 58 78
rect -2 68 24 69
rect 2 64 3 68
rect 7 64 8 68
rect 23 65 24 68
rect 28 68 45 69
rect 28 65 29 68
rect 44 65 45 68
rect 49 68 58 69
rect 49 65 50 68
rect 2 61 8 64
rect 2 57 3 61
rect 7 57 8 61
rect 13 62 17 63
rect 44 62 50 65
rect 13 55 17 58
rect 2 51 13 54
rect 2 50 17 51
rect 23 58 35 62
rect 39 58 40 62
rect 44 58 45 62
rect 49 58 50 62
rect 2 21 6 50
rect 10 38 14 39
rect 23 38 27 58
rect 33 50 46 54
rect 42 46 46 50
rect 31 42 32 46
rect 36 42 38 46
rect 19 34 20 38
rect 24 34 30 38
rect 10 29 14 34
rect 10 25 22 29
rect 2 17 7 21
rect 11 17 12 21
rect 18 17 22 25
rect 26 21 30 34
rect 34 31 38 42
rect 42 41 46 42
rect 34 25 46 31
rect 26 17 43 21
rect 47 17 48 21
rect -2 8 25 12
rect 29 8 58 12
rect -2 2 58 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
<< ntransistor >>
rect 13 10 15 30
rect 20 10 22 30
rect 32 13 34 30
rect 39 13 41 30
<< ptransistor >>
rect 9 45 11 69
rect 19 45 21 69
rect 31 50 33 70
rect 41 50 43 70
<< polycontact >>
rect 32 42 36 46
rect 42 42 46 46
rect 10 34 14 38
rect 20 34 24 38
<< ndcontact >>
rect 7 17 11 21
rect 43 17 47 21
rect 25 8 29 12
<< pdcontact >>
rect 3 64 7 68
rect 3 57 7 61
rect 13 58 17 62
rect 13 51 17 55
rect 24 65 28 69
rect 35 58 39 62
rect 45 65 49 69
rect 45 58 49 62
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
<< psubstratepdiff >>
rect 0 2 56 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 56 2
rect 0 -3 56 -2
<< nsubstratendiff >>
rect 0 82 56 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 56 82
rect 0 77 56 78
<< labels >>
rlabel polycontact 22 36 22 36 6 an
rlabel metal1 4 32 4 32 6 z
rlabel metal1 20 20 20 20 6 b
rlabel metal1 12 32 12 32 6 b
rlabel metal1 12 52 12 52 6 z
rlabel metal1 28 6 28 6 6 vss
rlabel metal1 24 36 24 36 6 an
rlabel metal1 36 32 36 32 6 a2
rlabel metal1 36 52 36 52 6 a1
rlabel metal1 31 60 31 60 6 an
rlabel metal1 28 74 28 74 6 vdd
rlabel metal1 37 19 37 19 6 an
rlabel metal1 44 28 44 28 6 a2
rlabel polycontact 44 44 44 44 6 a1
<< end >>
