.subckt nr2av0x1 a b vdd vss z
*   SPICE3 file   created from nr2av0x1.ext -      technology: scmos
m00 vdd    vdd    w1     vdd p w=28u  l=2.3636u ad=182.667p pd=56.6667u as=196p     ps=70u
m01 w2     a      vdd    vdd p w=28u  l=2.3636u ad=196p     pd=70u      as=182.667p ps=56.6667u
m02 w3     w2     vdd    vdd p w=28u  l=2.3636u ad=176p     pd=50u      as=182.667p ps=56.6667u
m03 z      b      w3     vdd p w=28u  l=2.3636u ad=196p     pd=70u      as=176p     ps=50u
m04 vss    vdd    w4     vss n w=20u  l=2.3636u ad=138p     pd=48u      as=140p     ps=54u
m05 w2     a      vss    vss n w=20u  l=2.3636u ad=140p     pd=54u      as=138p     ps=48u
m06 z      w2     vss    vss n w=20u  l=2.3636u ad=136p     pd=42u      as=138p     ps=48u
m07 vss    b      z      vss n w=20u  l=2.3636u ad=138p     pd=48u      as=136p     ps=42u
C0  b      a      0.033f
C1  vss    z      0.090f
C2  w2     a      0.157f
C3  w3     vdd    0.010f
C4  vss    b      0.049f
C5  a      vdd    0.118f
C6  z      b      0.222f
C7  vss    w2     0.134f
C8  z      w2     0.122f
C9  vss    vdd    0.014f
C10 z      vdd    0.024f
C11 b      w2     0.104f
C12 b      vdd    0.022f
C13 w2     vdd    0.068f
C14 vss    a      0.036f
C15 z      w3     0.023f
C16 z      a      0.025f
C18 z      vss    0.006f
C19 b      vss    0.045f
C20 w2     vss    0.050f
C21 a      vss    0.049f
.ends
