magic
tech scmos
timestamp 1179386034
<< checkpaint >>
rect -22 -22 46 94
<< ab >>
rect 0 0 24 72
<< pwell >>
rect -4 -4 28 32
<< nwell >>
rect -4 32 28 76
<< polysilicon >>
rect 9 57 11 61
rect 9 35 11 39
rect 9 34 15 35
rect 9 30 10 34
rect 14 30 15 34
rect 9 29 15 30
rect 9 24 11 29
rect 9 11 11 15
<< ndiffusion >>
rect 2 23 9 24
rect 2 19 3 23
rect 7 19 9 23
rect 2 18 9 19
rect 4 15 9 18
rect 11 15 20 24
rect 13 8 20 15
rect 13 4 14 8
rect 18 4 20 8
rect 13 3 20 4
<< pdiffusion >>
rect 13 68 20 69
rect 13 64 14 68
rect 18 64 20 68
rect 13 57 20 64
rect 4 52 9 57
rect 2 51 9 52
rect 2 47 3 51
rect 7 47 9 51
rect 2 44 9 47
rect 2 40 3 44
rect 7 40 9 44
rect 2 39 9 40
rect 11 39 20 57
<< metal1 >>
rect -2 68 26 72
rect -2 64 4 68
rect 8 64 14 68
rect 18 64 26 68
rect 2 53 14 59
rect 2 51 7 53
rect 2 47 3 51
rect 2 44 7 47
rect 2 40 3 44
rect 2 39 7 40
rect 2 24 6 39
rect 18 35 22 59
rect 10 34 22 35
rect 14 30 22 34
rect 10 29 22 30
rect 2 23 7 24
rect 2 19 3 23
rect 2 13 14 19
rect 18 13 22 29
rect -2 4 4 8
rect 8 4 14 8
rect 18 4 26 8
rect -2 0 26 4
<< ntransistor >>
rect 9 15 11 24
<< ptransistor >>
rect 9 39 11 57
<< polycontact >>
rect 10 30 14 34
<< ndcontact >>
rect 3 19 7 23
rect 14 4 18 8
<< pdcontact >>
rect 14 64 18 68
rect 3 47 7 51
rect 3 40 7 44
<< psubstratepcontact >>
rect 4 4 8 8
<< nsubstratencontact >>
rect 4 64 8 68
<< psubstratepdiff >>
rect 3 8 9 9
rect 3 4 4 8
rect 8 4 9 8
rect 3 3 9 4
<< nsubstratendiff >>
rect 3 68 9 69
rect 3 64 4 68
rect 8 64 9 68
rect 3 63 9 64
<< labels >>
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 4 12 4 6 vss
rlabel metal1 12 16 12 16 6 z
rlabel polycontact 12 32 12 32 6 a
rlabel metal1 12 56 12 56 6 z
rlabel metal1 12 68 12 68 6 vdd
rlabel metal1 20 36 20 36 6 a
<< end >>
