magic
tech scmos
timestamp 1180600681
<< checkpaint >>
rect -22 -22 72 122
<< ab >>
rect 0 0 50 100
<< pwell >>
rect -4 -4 54 48
<< nwell >>
rect -4 48 54 104
<< polysilicon >>
rect 13 86 15 90
rect 25 85 27 89
rect 37 85 39 89
rect 13 63 15 66
rect 7 62 15 63
rect 7 58 8 62
rect 12 58 15 62
rect 7 57 15 58
rect 11 24 13 57
rect 25 43 27 65
rect 17 42 27 43
rect 17 38 18 42
rect 22 38 27 42
rect 17 37 27 38
rect 19 24 21 37
rect 37 33 39 65
rect 27 32 39 33
rect 27 28 28 32
rect 32 31 39 32
rect 32 28 33 31
rect 27 27 33 28
rect 27 24 29 27
rect 11 2 13 6
rect 19 2 21 6
rect 27 2 29 6
<< ndiffusion >>
rect 33 24 43 25
rect 3 12 11 24
rect 3 8 4 12
rect 8 8 11 12
rect 3 6 11 8
rect 13 6 19 24
rect 21 6 27 24
rect 29 22 43 24
rect 29 18 38 22
rect 42 18 43 22
rect 29 15 43 18
rect 29 6 34 15
<< pdiffusion >>
rect 5 92 11 93
rect 5 88 6 92
rect 10 88 11 92
rect 29 92 35 93
rect 5 86 11 88
rect 5 66 13 86
rect 15 85 23 86
rect 29 88 30 92
rect 34 88 35 92
rect 29 85 35 88
rect 15 82 25 85
rect 15 78 18 82
rect 22 78 25 82
rect 15 66 25 78
rect 20 65 25 66
rect 27 65 37 85
rect 39 82 47 85
rect 39 78 42 82
rect 46 78 47 82
rect 39 65 47 78
<< metal1 >>
rect -2 92 52 100
rect -2 88 6 92
rect 10 88 30 92
rect 34 88 52 92
rect 8 62 12 83
rect 17 78 18 82
rect 22 78 42 82
rect 46 78 47 82
rect 8 17 12 58
rect 18 42 22 73
rect 18 17 22 38
rect 28 32 32 73
rect 28 17 32 28
rect 38 22 42 78
rect 38 17 42 18
rect -2 8 4 12
rect 8 8 52 12
rect -2 0 52 8
<< ntransistor >>
rect 11 6 13 24
rect 19 6 21 24
rect 27 6 29 24
<< ptransistor >>
rect 13 66 15 86
rect 25 65 27 85
rect 37 65 39 85
<< polycontact >>
rect 8 58 12 62
rect 18 38 22 42
rect 28 28 32 32
<< ndcontact >>
rect 4 8 8 12
rect 38 18 42 22
<< pdcontact >>
rect 6 88 10 92
rect 30 88 34 92
rect 18 78 22 82
rect 42 78 46 82
<< labels >>
rlabel metal1 20 45 20 45 6 i1
rlabel metal1 10 50 10 50 6 i0
rlabel pdcontact 20 80 20 80 6 nq
rlabel metal1 25 6 25 6 6 vss
rlabel metal1 30 45 30 45 6 i2
rlabel metal1 25 94 25 94 6 vdd
rlabel metal1 30 80 30 80 6 nq
rlabel metal1 40 50 40 50 6 nq
<< end >>
