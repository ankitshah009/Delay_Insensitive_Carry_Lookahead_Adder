magic
tech scmos
timestamp 1182286859
<< checkpaint >>
rect -22 -22 190 94
<< ab >>
rect 0 0 168 72
<< pwell >>
rect -4 -4 172 32
<< nwell >>
rect -4 32 172 76
<< polysilicon >>
rect 9 65 11 70
rect 19 65 21 70
rect 29 68 53 70
rect 29 65 31 68
rect 39 65 41 68
rect 51 51 53 68
rect 62 66 64 70
rect 72 66 74 70
rect 82 66 84 70
rect 92 66 94 70
rect 112 66 114 70
rect 122 66 124 70
rect 132 66 134 70
rect 48 50 54 51
rect 48 46 49 50
rect 53 46 54 50
rect 48 45 54 46
rect 9 35 11 38
rect 19 35 21 38
rect 29 35 31 38
rect 39 35 41 38
rect 62 37 64 40
rect 72 37 74 40
rect 143 60 158 61
rect 143 59 153 60
rect 143 56 145 59
rect 152 56 153 59
rect 157 56 158 60
rect 152 55 158 56
rect 153 52 155 55
rect 143 38 145 42
rect 9 34 22 35
rect 9 33 17 34
rect 16 30 17 33
rect 21 30 22 34
rect 29 33 41 35
rect 61 35 74 37
rect 82 35 84 38
rect 92 35 94 38
rect 112 35 114 38
rect 122 35 124 38
rect 61 34 67 35
rect 16 29 22 30
rect 9 24 11 29
rect 16 27 28 29
rect 16 24 18 27
rect 26 24 28 27
rect 33 24 35 33
rect 61 31 62 34
rect 45 26 47 31
rect 55 30 62 31
rect 66 30 67 34
rect 79 34 108 35
rect 79 33 103 34
rect 79 31 81 33
rect 55 29 67 30
rect 55 26 57 29
rect 65 26 67 29
rect 75 29 81 31
rect 102 30 103 33
rect 107 30 108 34
rect 102 29 108 30
rect 112 34 118 35
rect 112 30 113 34
rect 117 30 118 34
rect 112 29 118 30
rect 122 34 128 35
rect 122 30 123 34
rect 127 30 128 34
rect 132 34 134 38
rect 132 33 146 34
rect 132 32 141 33
rect 122 29 128 30
rect 140 29 141 32
rect 145 29 146 33
rect 75 26 77 29
rect 85 28 91 29
rect 85 24 86 28
rect 90 25 91 28
rect 90 24 97 25
rect 85 23 97 24
rect 85 20 87 23
rect 95 20 97 23
rect 113 20 115 29
rect 122 25 124 29
rect 140 28 146 29
rect 140 25 142 28
rect 153 26 155 38
rect 120 23 124 25
rect 120 20 122 23
rect 130 20 132 25
rect 9 4 11 12
rect 16 8 18 12
rect 26 8 28 12
rect 33 4 35 12
rect 9 2 35 4
rect 45 4 47 12
rect 55 8 57 12
rect 65 8 67 12
rect 75 4 77 12
rect 45 2 77 4
rect 85 3 87 8
rect 95 3 97 8
rect 140 8 142 12
rect 113 2 115 7
rect 120 2 122 7
rect 130 4 132 7
rect 153 4 155 15
rect 130 2 155 4
<< ndiffusion >>
rect 37 24 45 26
rect 2 17 9 24
rect 2 13 3 17
rect 7 13 9 17
rect 2 12 9 13
rect 11 12 16 24
rect 18 23 26 24
rect 18 19 20 23
rect 24 19 26 23
rect 18 12 26 19
rect 28 12 33 24
rect 35 12 45 24
rect 47 25 55 26
rect 47 21 49 25
rect 53 21 55 25
rect 47 12 55 21
rect 57 18 65 26
rect 57 14 59 18
rect 63 14 65 18
rect 57 12 65 14
rect 67 25 75 26
rect 67 21 69 25
rect 73 21 75 25
rect 67 18 75 21
rect 67 14 69 18
rect 73 14 75 18
rect 67 12 75 14
rect 77 20 82 26
rect 148 25 153 26
rect 135 20 140 25
rect 77 17 85 20
rect 77 13 79 17
rect 83 13 85 17
rect 77 12 85 13
rect 37 8 43 12
rect 37 4 38 8
rect 42 4 43 8
rect 37 3 43 4
rect 80 8 85 12
rect 87 18 95 20
rect 87 14 89 18
rect 93 14 95 18
rect 87 8 95 14
rect 97 11 113 20
rect 97 8 103 11
rect 99 7 103 8
rect 107 7 113 11
rect 115 7 120 20
rect 122 18 130 20
rect 122 14 124 18
rect 128 14 130 18
rect 122 7 130 14
rect 132 19 140 20
rect 132 15 134 19
rect 138 15 140 19
rect 132 12 140 15
rect 142 18 153 25
rect 142 14 146 18
rect 150 15 153 18
rect 155 25 162 26
rect 155 21 157 25
rect 161 21 162 25
rect 155 20 162 21
rect 155 15 160 20
rect 150 14 151 15
rect 142 12 151 14
rect 132 7 137 12
rect 99 5 111 7
<< pdiffusion >>
rect 4 58 9 65
rect 2 57 9 58
rect 2 53 3 57
rect 7 53 9 57
rect 2 50 9 53
rect 2 46 3 50
rect 7 46 9 50
rect 2 45 9 46
rect 4 38 9 45
rect 11 50 19 65
rect 11 46 13 50
rect 17 46 19 50
rect 11 43 19 46
rect 11 39 13 43
rect 17 39 19 43
rect 11 38 19 39
rect 21 58 29 65
rect 21 54 23 58
rect 27 54 29 58
rect 21 38 29 54
rect 31 43 39 65
rect 31 39 33 43
rect 37 39 39 43
rect 31 38 39 39
rect 41 59 46 65
rect 41 58 49 59
rect 41 54 44 58
rect 48 54 49 58
rect 41 53 49 54
rect 41 38 46 53
rect 55 65 62 66
rect 55 61 56 65
rect 60 61 62 65
rect 55 58 62 61
rect 55 54 56 58
rect 60 54 62 58
rect 55 53 62 54
rect 56 40 62 53
rect 64 57 72 66
rect 64 53 66 57
rect 70 53 72 57
rect 64 50 72 53
rect 64 46 66 50
rect 70 46 72 50
rect 64 40 72 46
rect 74 65 82 66
rect 74 61 76 65
rect 80 61 82 65
rect 74 58 82 61
rect 74 54 76 58
rect 80 54 82 58
rect 74 40 82 54
rect 77 38 82 40
rect 84 43 92 66
rect 84 39 86 43
rect 90 39 92 43
rect 84 38 92 39
rect 94 65 101 66
rect 94 61 96 65
rect 100 61 101 65
rect 94 58 101 61
rect 107 59 112 66
rect 94 54 96 58
rect 100 54 101 58
rect 94 38 101 54
rect 105 58 112 59
rect 105 54 106 58
rect 110 54 112 58
rect 105 53 112 54
rect 107 38 112 53
rect 114 51 122 66
rect 114 47 116 51
rect 120 47 122 51
rect 114 38 122 47
rect 124 50 132 66
rect 124 46 126 50
rect 130 46 132 50
rect 124 43 132 46
rect 124 39 126 43
rect 130 39 132 43
rect 124 38 132 39
rect 134 65 141 66
rect 134 61 136 65
rect 140 61 141 65
rect 160 68 166 69
rect 160 64 161 68
rect 165 64 166 68
rect 134 56 141 61
rect 134 42 143 56
rect 145 52 150 56
rect 160 52 166 64
rect 145 47 153 52
rect 145 43 147 47
rect 151 43 153 47
rect 145 42 153 43
rect 134 38 141 42
rect 148 38 153 42
rect 155 38 166 52
<< metal1 >>
rect -2 68 170 72
rect -2 65 149 68
rect -2 64 56 65
rect 55 61 56 64
rect 60 64 76 65
rect 60 61 61 64
rect 55 58 61 61
rect 75 61 76 64
rect 80 64 96 65
rect 80 61 81 64
rect 75 58 81 61
rect 2 57 23 58
rect 2 53 3 57
rect 7 54 23 57
rect 27 54 44 58
rect 48 54 49 58
rect 55 54 56 58
rect 60 54 61 58
rect 66 57 70 58
rect 2 50 7 53
rect 75 54 76 58
rect 80 54 81 58
rect 95 61 96 64
rect 100 64 136 65
rect 100 61 101 64
rect 135 61 136 64
rect 140 64 149 65
rect 153 64 161 68
rect 165 64 170 68
rect 140 61 141 64
rect 95 58 101 61
rect 95 54 96 58
rect 100 54 101 58
rect 105 54 106 58
rect 110 54 138 58
rect 66 50 70 53
rect 2 46 3 50
rect 2 45 7 46
rect 12 46 13 50
rect 17 46 49 50
rect 53 46 66 50
rect 70 46 99 50
rect 2 26 6 45
rect 12 43 17 46
rect 12 39 13 43
rect 12 38 17 39
rect 32 39 33 43
rect 37 39 38 43
rect 85 42 86 43
rect 32 34 38 39
rect 48 39 86 42
rect 90 39 91 43
rect 48 38 91 39
rect 48 34 52 38
rect 16 30 17 34
rect 21 30 52 34
rect 57 30 62 34
rect 66 30 87 34
rect 2 23 24 26
rect 2 22 20 23
rect 48 25 52 30
rect 81 28 87 30
rect 48 21 49 25
rect 53 21 69 25
rect 73 21 74 25
rect 81 24 86 28
rect 90 24 91 28
rect 81 22 87 24
rect 20 18 24 19
rect 69 18 74 21
rect 95 18 99 46
rect 3 17 7 18
rect 20 14 59 18
rect 63 14 64 18
rect 73 14 74 18
rect 69 13 74 14
rect 79 17 83 18
rect 88 14 89 18
rect 93 14 99 18
rect 103 47 116 51
rect 120 47 121 51
rect 126 50 130 51
rect 103 34 107 47
rect 126 43 130 46
rect 103 18 107 30
rect 113 39 126 42
rect 113 38 130 39
rect 134 42 138 54
rect 152 56 153 60
rect 157 59 158 60
rect 157 56 166 59
rect 152 53 166 56
rect 147 47 151 48
rect 162 45 166 53
rect 147 42 151 43
rect 134 38 166 42
rect 113 34 117 38
rect 134 34 138 38
rect 145 34 158 35
rect 122 30 123 34
rect 127 30 138 34
rect 141 33 158 34
rect 113 26 117 30
rect 145 29 158 33
rect 141 28 151 29
rect 113 22 138 26
rect 145 22 151 28
rect 162 25 166 38
rect 134 19 138 22
rect 156 21 157 25
rect 161 21 166 25
rect 103 14 124 18
rect 128 14 129 18
rect 134 14 138 15
rect 145 14 146 18
rect 150 14 151 18
rect 3 8 7 13
rect 79 8 83 13
rect 102 8 103 11
rect -2 4 38 8
rect 42 7 103 8
rect 107 8 108 11
rect 145 8 151 14
rect 107 7 159 8
rect 42 4 159 7
rect 163 4 170 8
rect -2 0 170 4
<< ntransistor >>
rect 9 12 11 24
rect 16 12 18 24
rect 26 12 28 24
rect 33 12 35 24
rect 45 12 47 26
rect 55 12 57 26
rect 65 12 67 26
rect 75 12 77 26
rect 85 8 87 20
rect 95 8 97 20
rect 113 7 115 20
rect 120 7 122 20
rect 130 7 132 20
rect 140 12 142 25
rect 153 15 155 26
<< ptransistor >>
rect 9 38 11 65
rect 19 38 21 65
rect 29 38 31 65
rect 39 38 41 65
rect 62 40 64 66
rect 72 40 74 66
rect 82 38 84 66
rect 92 38 94 66
rect 112 38 114 66
rect 122 38 124 66
rect 132 38 134 66
rect 143 42 145 56
rect 153 38 155 52
<< polycontact >>
rect 49 46 53 50
rect 153 56 157 60
rect 17 30 21 34
rect 62 30 66 34
rect 103 30 107 34
rect 113 30 117 34
rect 123 30 127 34
rect 141 29 145 33
rect 86 24 90 28
<< ndcontact >>
rect 3 13 7 17
rect 20 19 24 23
rect 49 21 53 25
rect 59 14 63 18
rect 69 21 73 25
rect 69 14 73 18
rect 79 13 83 17
rect 38 4 42 8
rect 89 14 93 18
rect 103 7 107 11
rect 124 14 128 18
rect 134 15 138 19
rect 146 14 150 18
rect 157 21 161 25
<< pdcontact >>
rect 3 53 7 57
rect 3 46 7 50
rect 13 46 17 50
rect 13 39 17 43
rect 23 54 27 58
rect 33 39 37 43
rect 44 54 48 58
rect 56 61 60 65
rect 56 54 60 58
rect 66 53 70 57
rect 66 46 70 50
rect 76 61 80 65
rect 76 54 80 58
rect 86 39 90 43
rect 96 61 100 65
rect 96 54 100 58
rect 106 54 110 58
rect 116 47 120 51
rect 126 46 130 50
rect 126 39 130 43
rect 136 61 140 65
rect 161 64 165 68
rect 147 43 151 47
<< psubstratepcontact >>
rect 159 4 163 8
<< nsubstratencontact >>
rect 149 64 153 68
<< psubstratepdiff >>
rect 157 8 165 9
rect 157 4 159 8
rect 163 4 165 8
rect 157 3 165 4
<< nsubstratendiff >>
rect 145 68 156 69
rect 145 64 149 68
rect 153 64 156 68
rect 145 63 156 64
<< labels >>
rlabel polysilicon 52 57 52 57 6 cn
rlabel ntransistor 114 18 114 18 6 an
rlabel polycontact 105 32 105 32 6 iz
rlabel polycontact 125 32 125 32 6 bn
rlabel metal1 28 16 28 16 6 z
rlabel metal1 20 24 20 24 6 z
rlabel metal1 12 24 12 24 6 z
rlabel metal1 4 40 4 40 6 z
rlabel metal1 14 44 14 44 6 cn
rlabel metal1 12 56 12 56 6 z
rlabel metal1 20 56 20 56 6 z
rlabel metal1 28 56 28 56 6 z
rlabel metal1 36 16 36 16 6 z
rlabel metal1 44 16 44 16 6 z
rlabel metal1 52 16 52 16 6 z
rlabel ndcontact 60 16 60 16 6 z
rlabel metal1 60 32 60 32 6 c
rlabel metal1 35 36 35 36 6 zn
rlabel metal1 36 56 36 56 6 z
rlabel metal1 44 56 44 56 6 z
rlabel metal1 84 4 84 4 6 vss
rlabel metal1 71 19 71 19 6 zn
rlabel metal1 93 16 93 16 6 cn
rlabel metal1 61 23 61 23 6 zn
rlabel metal1 76 32 76 32 6 c
rlabel metal1 84 28 84 28 6 c
rlabel metal1 68 32 68 32 6 c
rlabel pdcontact 88 40 88 40 6 zn
rlabel metal1 55 48 55 48 6 cn
rlabel metal1 68 52 68 52 6 cn
rlabel metal1 84 68 84 68 6 vdd
rlabel metal1 116 16 116 16 6 iz
rlabel polycontact 115 32 115 32 6 an
rlabel metal1 128 44 128 44 6 an
rlabel polycontact 105 32 105 32 6 iz
rlabel metal1 112 49 112 49 6 iz
rlabel metal1 136 20 136 20 6 an
rlabel metal1 161 23 161 23 6 bn
rlabel metal1 148 28 148 28 6 a
rlabel metal1 156 32 156 32 6 a
rlabel metal1 130 32 130 32 6 bn
rlabel metal1 149 43 149 43 6 bn
rlabel metal1 164 52 164 52 6 b
rlabel metal1 156 56 156 56 6 b
rlabel metal1 121 56 121 56 6 bn
<< end >>
