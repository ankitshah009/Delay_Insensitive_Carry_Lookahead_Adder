.subckt xaoi21_x1 a1 a2 b vdd vss z
*   SPICE3 file   created from xaoi21_x1.ext -      technology: scmos
m00 an     a1     vdd    vdd p w=38u  l=2.3636u ad=204p     pd=62.6667u as=223p     ps=70u
m01 vdd    a2     an     vdd p w=38u  l=2.3636u ad=223p     pd=70u      as=204p     ps=62.6667u
m02 z      b      an     vdd p w=38u  l=2.3636u ad=190p     pd=48u      as=204p     ps=62.6667u
m03 w1     bn     z      vdd p w=38u  l=2.3636u ad=114p     pd=44u      as=190p     ps=48u
m04 vdd    an     w1     vdd p w=38u  l=2.3636u ad=223p     pd=70u      as=114p     ps=44u
m05 bn     b      vdd    vdd p w=38u  l=2.3636u ad=232p     pd=92u      as=223p     ps=70u
m06 w2     a1     vss    vss n w=24u  l=2.3636u ad=72p      pd=30u      as=220.098p ps=71.4146u
m07 an     a2     w2     vss n w=24u  l=2.3636u ad=120p     pd=34u      as=72p      ps=30u
m08 z      bn     an     vss n w=24u  l=2.3636u ad=120p     pd=39.8049u as=120p     ps=34u
m09 bn     an     z      vss n w=17u  l=2.3636u ad=85p      pd=27u      as=85p      ps=28.1951u
m10 vss    b      bn     vss n w=17u  l=2.3636u ad=155.902p pd=50.5854u as=85p      ps=27u
C0  z      bn     0.101f
C1  w1     an     0.022f
C2  w1     b      0.012f
C3  vss    a2     0.010f
C4  w2     a1     0.009f
C5  z      vdd    0.033f
C6  bn     an     0.339f
C7  bn     b      0.293f
C8  an     vdd    0.237f
C9  z      a2     0.066f
C10 an     a2     0.241f
C11 bn     a1     0.039f
C12 vdd    b      0.294f
C13 vss    z      0.071f
C14 vdd    a1     0.008f
C15 b      a2     0.032f
C16 vss    an     0.234f
C17 a2     a1     0.225f
C18 vss    b      0.011f
C19 z      an     0.394f
C20 w1     vdd    0.010f
C21 vss    a1     0.060f
C22 bn     vdd    0.019f
C23 z      b      0.076f
C24 w2     vss    0.010f
C25 z      a1     0.067f
C26 bn     a2     0.043f
C27 an     b      0.435f
C28 vdd    a2     0.035f
C29 an     a1     0.287f
C30 vss    bn     0.147f
C31 w2     an     0.012f
C32 b      a1     0.010f
C34 z      vss    0.019f
C35 bn     vss    0.049f
C36 an     vss    0.056f
C38 b      vss    0.050f
C39 a2     vss    0.028f
C40 a1     vss    0.033f
.ends
