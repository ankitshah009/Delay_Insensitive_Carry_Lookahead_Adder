magic
tech scmos
timestamp 1179385947
<< checkpaint >>
rect -22 -25 54 105
<< ab >>
rect 0 0 32 80
<< pwell >>
rect -4 -7 36 36
<< nwell >>
rect -4 36 36 87
<< polysilicon >>
rect 11 58 13 63
rect 21 58 23 63
rect 11 39 13 42
rect 21 39 23 42
rect 11 38 23 39
rect 11 34 18 38
rect 22 34 23 38
rect 11 33 23 34
rect 15 30 17 33
rect 15 17 17 22
<< ndiffusion >>
rect 8 29 15 30
rect 8 25 9 29
rect 13 25 15 29
rect 8 24 15 25
rect 10 22 15 24
rect 17 27 25 30
rect 17 23 19 27
rect 23 23 25 27
rect 17 22 25 23
<< pdiffusion >>
rect 2 57 11 58
rect 2 53 3 57
rect 7 53 11 57
rect 2 50 11 53
rect 2 46 3 50
rect 7 46 11 50
rect 2 42 11 46
rect 13 55 21 58
rect 13 51 15 55
rect 19 51 21 55
rect 13 48 21 51
rect 13 44 15 48
rect 19 44 21 48
rect 13 42 21 44
rect 23 57 30 58
rect 23 53 25 57
rect 29 53 30 57
rect 23 50 30 53
rect 23 46 25 50
rect 29 46 30 50
rect 23 42 30 46
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect -2 68 34 78
rect 3 57 7 68
rect 25 57 29 68
rect 3 50 7 53
rect 15 55 22 56
rect 19 51 22 55
rect 15 49 22 51
rect 25 50 29 53
rect 15 48 19 49
rect 3 45 7 46
rect 10 44 15 47
rect 25 45 29 46
rect 10 43 19 44
rect 10 30 14 43
rect 18 38 30 39
rect 22 34 30 38
rect 18 33 30 34
rect 9 29 14 30
rect 13 25 14 29
rect 9 24 14 25
rect 19 27 23 28
rect 26 25 30 33
rect 19 12 23 23
rect -2 2 34 12
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
<< ntransistor >>
rect 15 22 17 30
<< ptransistor >>
rect 11 42 13 58
rect 21 42 23 58
<< polycontact >>
rect 18 34 22 38
<< ndcontact >>
rect 9 25 13 29
rect 19 23 23 27
<< pdcontact >>
rect 3 53 7 57
rect 3 46 7 50
rect 15 51 19 55
rect 15 44 19 48
rect 25 53 29 57
rect 25 46 29 50
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
<< psubstratepdiff >>
rect 0 2 32 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 32 2
rect 0 -3 32 -2
<< nsubstratendiff >>
rect 0 82 32 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 32 82
rect 0 77 32 78
<< labels >>
rlabel metal1 12 36 12 36 6 z
rlabel metal1 16 6 16 6 6 vss
rlabel polycontact 20 36 20 36 6 a
rlabel metal1 20 52 20 52 6 z
rlabel metal1 16 74 16 74 6 vdd
rlabel metal1 28 32 28 32 6 a
<< end >>
