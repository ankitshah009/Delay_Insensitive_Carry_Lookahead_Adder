magic
tech scmos
timestamp 1179385099
<< checkpaint >>
rect -22 -25 78 105
<< ab >>
rect 0 0 56 80
<< pwell >>
rect -4 -7 60 36
<< nwell >>
rect -4 36 60 87
<< polysilicon >>
rect 9 64 11 69
rect 19 64 21 69
rect 29 64 31 69
rect 41 64 43 69
rect 19 47 21 58
rect 29 55 31 58
rect 29 54 37 55
rect 29 50 32 54
rect 36 50 37 54
rect 29 49 37 50
rect 19 46 25 47
rect 9 39 11 46
rect 19 42 20 46
rect 24 42 25 46
rect 19 41 25 42
rect 9 38 15 39
rect 9 34 10 38
rect 14 34 15 38
rect 9 33 15 34
rect 9 26 11 33
rect 22 23 24 41
rect 29 23 31 49
rect 41 32 43 58
rect 40 31 46 32
rect 40 28 41 31
rect 36 27 41 28
rect 45 27 46 31
rect 36 26 46 27
rect 36 23 38 26
rect 9 12 11 17
rect 22 12 24 17
rect 29 12 31 17
rect 36 12 38 17
<< ndiffusion >>
rect 4 23 9 26
rect 2 22 9 23
rect 2 18 3 22
rect 7 18 9 22
rect 2 17 9 18
rect 11 23 20 26
rect 11 17 22 23
rect 24 17 29 23
rect 31 17 36 23
rect 38 22 45 23
rect 38 18 40 22
rect 44 18 45 22
rect 38 17 45 18
rect 13 12 20 17
rect 13 8 14 12
rect 18 8 20 12
rect 13 7 20 8
<< pdiffusion >>
rect 33 72 39 73
rect 33 68 34 72
rect 38 68 39 72
rect 33 64 39 68
rect 4 59 9 64
rect 2 58 9 59
rect 2 54 3 58
rect 7 54 9 58
rect 2 51 9 54
rect 2 47 3 51
rect 7 47 9 51
rect 2 46 9 47
rect 11 63 19 64
rect 11 59 13 63
rect 17 59 19 63
rect 11 58 19 59
rect 21 63 29 64
rect 21 59 23 63
rect 27 59 29 63
rect 21 58 29 59
rect 31 58 41 64
rect 43 63 50 64
rect 43 59 45 63
rect 49 59 50 63
rect 43 58 50 59
rect 11 46 17 58
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect -2 72 58 78
rect -2 68 34 72
rect 38 68 58 72
rect 13 63 17 68
rect 2 58 7 63
rect 13 58 17 59
rect 22 59 23 63
rect 27 59 45 63
rect 49 59 50 63
rect 2 54 3 58
rect 22 54 26 59
rect 2 51 7 54
rect 2 47 3 51
rect 2 46 7 47
rect 10 50 26 54
rect 31 50 32 54
rect 36 50 47 54
rect 2 22 6 46
rect 10 38 14 50
rect 17 42 20 46
rect 24 42 31 46
rect 41 42 47 50
rect 25 34 31 42
rect 10 30 14 34
rect 41 31 47 38
rect 10 26 22 30
rect 25 27 41 30
rect 45 27 47 31
rect 25 26 47 27
rect 18 22 22 26
rect 2 18 3 22
rect 7 18 15 22
rect 18 18 40 22
rect 44 18 45 22
rect -2 8 14 12
rect 18 8 58 12
rect -2 2 58 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
<< ntransistor >>
rect 9 17 11 26
rect 22 17 24 23
rect 29 17 31 23
rect 36 17 38 23
<< ptransistor >>
rect 9 46 11 64
rect 19 58 21 64
rect 29 58 31 64
rect 41 58 43 64
<< polycontact >>
rect 32 50 36 54
rect 20 42 24 46
rect 10 34 14 38
rect 41 27 45 31
<< ndcontact >>
rect 3 18 7 22
rect 40 18 44 22
rect 14 8 18 12
<< pdcontact >>
rect 34 68 38 72
rect 3 54 7 58
rect 3 47 7 51
rect 13 59 17 63
rect 23 59 27 63
rect 45 59 49 63
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
<< psubstratepdiff >>
rect 0 2 56 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 56 2
rect 0 -3 56 -2
<< nsubstratendiff >>
rect 0 82 56 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 56 82
rect 0 77 56 78
<< labels >>
rlabel polycontact 12 36 12 36 6 zn
rlabel metal1 4 44 4 44 6 z
rlabel metal1 12 20 12 20 6 z
rlabel metal1 20 44 20 44 6 a
rlabel metal1 12 40 12 40 6 zn
rlabel metal1 28 6 28 6 6 vss
rlabel metal1 28 28 28 28 6 c
rlabel metal1 36 28 36 28 6 c
rlabel metal1 28 40 28 40 6 a
rlabel metal1 36 52 36 52 6 b
rlabel metal1 28 74 28 74 6 vdd
rlabel metal1 31 20 31 20 6 zn
rlabel metal1 44 32 44 32 6 c
rlabel metal1 44 48 44 48 6 b
rlabel metal1 36 61 36 61 6 zn
<< end >>
