magic
tech scmos
timestamp 1179386882
<< checkpaint >>
rect -22 -25 86 105
<< ab >>
rect 0 0 64 80
<< pwell >>
rect -4 -7 68 36
<< nwell >>
rect -4 36 68 87
<< polysilicon >>
rect 11 70 13 74
rect 18 70 20 74
rect 25 70 27 74
rect 35 70 37 74
rect 42 70 44 74
rect 49 70 51 74
rect 11 31 13 42
rect 18 39 20 42
rect 25 39 27 42
rect 35 39 37 42
rect 18 36 21 39
rect 25 37 37 39
rect 19 31 21 36
rect 35 31 37 37
rect 9 30 15 31
rect 9 26 10 30
rect 14 26 15 30
rect 9 25 15 26
rect 19 30 25 31
rect 19 26 20 30
rect 24 26 25 30
rect 19 25 25 26
rect 31 30 37 31
rect 31 26 32 30
rect 36 26 37 30
rect 42 33 44 42
rect 49 39 51 42
rect 49 38 58 39
rect 49 37 53 38
rect 52 34 53 37
rect 57 34 58 38
rect 52 33 58 34
rect 42 32 48 33
rect 42 28 43 32
rect 47 28 48 32
rect 42 27 48 28
rect 31 25 37 26
rect 9 22 11 25
rect 21 22 23 25
rect 31 22 33 25
rect 9 7 11 12
rect 21 7 23 12
rect 31 7 33 12
<< ndiffusion >>
rect 2 21 9 22
rect 2 17 3 21
rect 7 17 9 21
rect 2 16 9 17
rect 4 12 9 16
rect 11 12 21 22
rect 23 21 31 22
rect 23 17 25 21
rect 29 17 31 21
rect 23 12 31 17
rect 33 12 42 22
rect 13 8 14 12
rect 18 8 19 12
rect 13 7 19 8
rect 35 8 36 12
rect 40 8 42 12
rect 35 7 42 8
<< pdiffusion >>
rect 4 69 11 70
rect 4 65 5 69
rect 9 65 11 69
rect 4 62 11 65
rect 4 58 5 62
rect 9 58 11 62
rect 4 42 11 58
rect 13 42 18 70
rect 20 42 25 70
rect 27 62 35 70
rect 27 58 29 62
rect 33 58 35 62
rect 27 55 35 58
rect 27 51 29 55
rect 33 51 35 55
rect 27 42 35 51
rect 37 42 42 70
rect 44 42 49 70
rect 51 69 58 70
rect 51 65 53 69
rect 57 65 58 69
rect 51 62 58 65
rect 51 58 53 62
rect 57 58 58 62
rect 51 42 58 58
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect -2 69 66 78
rect -2 68 5 69
rect 4 65 5 68
rect 9 68 53 69
rect 9 65 10 68
rect 4 62 10 65
rect 52 65 53 68
rect 57 68 66 69
rect 57 65 58 68
rect 4 58 5 62
rect 9 58 10 62
rect 29 62 33 63
rect 52 62 58 65
rect 52 58 53 62
rect 57 58 58 62
rect 29 55 33 58
rect 2 51 29 54
rect 33 51 39 54
rect 2 50 39 51
rect 2 21 6 50
rect 10 42 55 46
rect 10 30 14 42
rect 51 38 55 42
rect 10 25 14 26
rect 18 34 47 38
rect 51 34 53 38
rect 57 34 58 38
rect 18 30 24 34
rect 43 32 47 34
rect 18 26 20 30
rect 31 26 32 30
rect 36 26 39 30
rect 47 28 55 30
rect 43 26 55 28
rect 18 25 24 26
rect 34 22 39 26
rect 2 17 3 21
rect 7 17 25 21
rect 29 17 30 21
rect 34 17 47 22
rect -2 8 14 12
rect 18 8 36 12
rect 40 8 66 12
rect -2 2 66 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
<< ntransistor >>
rect 9 12 11 22
rect 21 12 23 22
rect 31 12 33 22
<< ptransistor >>
rect 11 42 13 70
rect 18 42 20 70
rect 25 42 27 70
rect 35 42 37 70
rect 42 42 44 70
rect 49 42 51 70
<< polycontact >>
rect 10 26 14 30
rect 20 26 24 30
rect 32 26 36 30
rect 53 34 57 38
rect 43 28 47 32
<< ndcontact >>
rect 3 17 7 21
rect 25 17 29 21
rect 14 8 18 12
rect 36 8 40 12
<< pdcontact >>
rect 5 65 9 69
rect 5 58 9 62
rect 29 58 33 62
rect 29 51 33 55
rect 53 65 57 69
rect 53 58 57 62
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
<< psubstratepdiff >>
rect 0 2 64 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 64 2
rect 0 -3 64 -2
<< nsubstratendiff >>
rect 0 82 64 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 64 82
rect 0 77 64 78
<< labels >>
rlabel metal1 4 32 4 32 6 z
rlabel metal1 20 28 20 28 6 b
rlabel metal1 12 32 12 32 6 a
rlabel metal1 20 44 20 44 6 a
rlabel metal1 20 52 20 52 6 z
rlabel metal1 12 52 12 52 6 z
rlabel metal1 32 6 32 6 6 vss
rlabel metal1 36 24 36 24 6 c
rlabel metal1 28 36 28 36 6 b
rlabel metal1 28 44 28 44 6 a
rlabel metal1 36 36 36 36 6 b
rlabel metal1 36 44 36 44 6 a
rlabel metal1 36 52 36 52 6 z
rlabel metal1 28 52 28 52 6 z
rlabel metal1 32 74 32 74 6 vdd
rlabel metal1 44 20 44 20 6 c
rlabel metal1 44 36 44 36 6 b
rlabel metal1 44 44 44 44 6 a
rlabel metal1 52 28 52 28 6 b
rlabel metal1 52 44 52 44 6 a
<< end >>
