magic
tech scmos
timestamp 1179387791
<< checkpaint >>
rect -22 -22 190 94
<< ab >>
rect 0 0 168 72
<< pwell >>
rect -4 -4 172 32
<< nwell >>
rect -4 32 172 76
<< polysilicon >>
rect 11 66 13 70
rect 19 66 21 70
rect 27 66 29 70
rect 37 66 39 70
rect 44 66 46 70
rect 54 66 56 70
rect 75 66 77 70
rect 104 66 106 70
rect 114 66 116 70
rect 121 66 123 70
rect 131 66 133 70
rect 139 66 141 70
rect 147 66 149 70
rect 86 43 92 44
rect 86 39 87 43
rect 91 39 92 43
rect 86 38 92 39
rect 159 44 165 45
rect 159 40 160 44
rect 164 40 165 44
rect 159 39 165 40
rect 11 35 13 38
rect 19 35 21 38
rect 27 35 29 38
rect 37 35 39 38
rect 44 35 46 38
rect 54 35 56 38
rect 75 35 77 38
rect 86 35 88 38
rect 2 34 13 35
rect 2 30 3 34
rect 7 30 13 34
rect 2 29 13 30
rect 17 34 23 35
rect 17 30 18 34
rect 22 30 23 34
rect 17 29 23 30
rect 27 34 40 35
rect 27 30 35 34
rect 39 30 40 34
rect 44 32 48 35
rect 54 32 58 35
rect 27 29 40 30
rect 11 26 13 29
rect 19 26 21 29
rect 27 26 29 29
rect 37 26 39 29
rect 46 28 48 32
rect 46 27 52 28
rect 46 23 47 27
rect 51 23 52 27
rect 46 22 52 23
rect 46 19 48 22
rect 56 19 58 32
rect 62 34 77 35
rect 62 30 63 34
rect 67 30 77 34
rect 62 29 77 30
rect 83 33 88 35
rect 104 34 106 38
rect 92 33 106 34
rect 68 26 70 29
rect 11 7 13 12
rect 19 7 21 12
rect 27 7 29 12
rect 37 7 39 12
rect 83 18 85 33
rect 92 29 93 33
rect 97 29 106 33
rect 92 28 106 29
rect 104 25 106 28
rect 114 25 116 38
rect 121 35 123 38
rect 131 35 133 38
rect 139 35 141 38
rect 147 35 149 38
rect 159 35 161 39
rect 121 34 133 35
rect 121 30 122 34
rect 126 30 133 34
rect 121 29 133 30
rect 137 34 143 35
rect 137 30 138 34
rect 142 30 143 34
rect 137 29 143 30
rect 147 33 161 35
rect 121 25 123 29
rect 131 25 133 29
rect 139 25 141 29
rect 147 25 149 33
rect 79 17 85 18
rect 79 13 80 17
rect 84 13 85 17
rect 79 12 85 13
rect 68 8 70 12
rect 160 18 166 19
rect 160 14 161 18
rect 165 14 166 18
rect 160 13 166 14
rect 104 8 106 12
rect 46 2 48 7
rect 56 4 58 7
rect 114 4 116 12
rect 121 8 123 12
rect 131 8 133 12
rect 139 8 141 12
rect 147 8 149 12
rect 160 4 162 13
rect 56 2 162 4
<< ndiffusion >>
rect 3 12 11 26
rect 13 12 19 26
rect 21 12 27 26
rect 29 25 37 26
rect 29 21 31 25
rect 35 21 37 25
rect 29 12 37 21
rect 39 19 44 26
rect 60 19 68 26
rect 39 12 46 19
rect 3 8 9 12
rect 3 4 4 8
rect 8 4 9 8
rect 41 7 46 12
rect 48 17 56 19
rect 48 13 50 17
rect 54 13 56 17
rect 48 7 56 13
rect 58 15 61 19
rect 65 15 68 19
rect 58 12 68 15
rect 70 18 75 26
rect 70 17 77 18
rect 70 13 72 17
rect 76 13 77 17
rect 70 12 77 13
rect 58 8 61 12
rect 65 8 66 12
rect 97 17 104 25
rect 97 13 98 17
rect 102 13 104 17
rect 97 12 104 13
rect 106 24 114 25
rect 106 20 108 24
rect 112 20 114 24
rect 106 17 114 20
rect 106 13 108 17
rect 112 13 114 17
rect 106 12 114 13
rect 116 12 121 25
rect 123 18 131 25
rect 123 14 125 18
rect 129 14 131 18
rect 123 12 131 14
rect 133 12 139 25
rect 141 12 147 25
rect 149 24 158 25
rect 149 20 153 24
rect 157 20 158 24
rect 149 17 158 20
rect 149 13 153 17
rect 157 13 158 17
rect 149 12 158 13
rect 58 7 66 8
rect 3 3 9 4
<< pdiffusion >>
rect 3 65 11 66
rect 3 61 5 65
rect 9 61 11 65
rect 3 38 11 61
rect 13 38 19 66
rect 21 38 27 66
rect 29 50 37 66
rect 29 46 31 50
rect 35 46 37 50
rect 29 38 37 46
rect 39 38 44 66
rect 46 58 54 66
rect 46 54 48 58
rect 52 54 54 58
rect 46 38 54 54
rect 56 65 75 66
rect 56 61 59 65
rect 63 61 69 65
rect 73 61 75 65
rect 56 38 75 61
rect 77 44 82 66
rect 97 65 104 66
rect 97 61 98 65
rect 102 61 104 65
rect 77 43 84 44
rect 77 39 79 43
rect 83 39 84 43
rect 77 38 84 39
rect 97 38 104 61
rect 106 43 114 66
rect 106 39 108 43
rect 112 39 114 43
rect 106 38 114 39
rect 116 38 121 66
rect 123 50 131 66
rect 123 46 125 50
rect 129 46 131 50
rect 123 38 131 46
rect 133 38 139 66
rect 141 38 147 66
rect 149 59 155 66
rect 149 58 157 59
rect 149 54 151 58
rect 155 54 157 58
rect 149 38 157 54
<< metal1 >>
rect -2 68 170 72
rect -2 65 87 68
rect -2 64 5 65
rect 4 61 5 64
rect 9 64 59 65
rect 9 61 10 64
rect 58 61 59 64
rect 63 61 69 65
rect 73 64 87 65
rect 91 65 160 68
rect 91 64 98 65
rect 73 61 74 64
rect 97 61 98 64
rect 102 64 160 65
rect 164 64 170 68
rect 102 61 103 64
rect 151 58 155 64
rect 3 54 48 58
rect 52 54 148 58
rect 3 34 7 54
rect 144 50 148 54
rect 151 53 155 54
rect 3 17 7 30
rect 10 46 31 50
rect 35 46 125 50
rect 129 46 141 50
rect 144 46 164 50
rect 10 25 14 46
rect 25 38 75 42
rect 78 39 79 43
rect 83 39 87 43
rect 91 39 104 43
rect 25 35 30 38
rect 18 34 30 35
rect 71 34 75 38
rect 100 34 104 39
rect 107 39 108 43
rect 112 42 113 43
rect 137 42 141 46
rect 160 44 164 46
rect 112 39 134 42
rect 107 38 134 39
rect 137 38 150 42
rect 160 39 164 40
rect 130 34 134 38
rect 22 30 30 34
rect 34 30 35 34
rect 39 30 63 34
rect 67 30 68 34
rect 71 33 97 34
rect 71 30 93 33
rect 18 29 30 30
rect 100 30 122 34
rect 126 30 127 34
rect 130 30 138 34
rect 142 30 143 34
rect 93 28 97 29
rect 10 21 31 25
rect 35 21 36 25
rect 46 23 47 27
rect 51 26 52 27
rect 130 26 134 30
rect 51 25 89 26
rect 107 25 134 26
rect 51 24 134 25
rect 51 23 108 24
rect 46 22 108 23
rect 85 21 108 22
rect 107 20 108 21
rect 112 22 134 24
rect 112 20 113 22
rect 3 13 50 17
rect 54 13 55 17
rect 60 15 61 19
rect 65 15 66 19
rect 107 17 113 20
rect 146 18 150 38
rect 154 29 166 35
rect 60 12 66 15
rect 71 13 72 17
rect 76 13 80 17
rect 84 13 85 17
rect 97 13 98 17
rect 102 13 103 17
rect 107 13 108 17
rect 112 13 113 17
rect 124 14 125 18
rect 129 14 150 18
rect 153 24 157 25
rect 153 17 157 20
rect 161 18 166 29
rect 165 14 166 18
rect 161 13 166 14
rect 60 8 61 12
rect 65 8 66 12
rect 88 11 92 12
rect -2 4 4 8
rect 8 7 88 8
rect 97 8 103 13
rect 153 8 157 13
rect 92 7 170 8
rect 8 4 170 7
rect -2 0 170 4
<< ntransistor >>
rect 11 12 13 26
rect 19 12 21 26
rect 27 12 29 26
rect 37 12 39 26
rect 46 7 48 19
rect 56 7 58 19
rect 68 12 70 26
rect 104 12 106 25
rect 114 12 116 25
rect 121 12 123 25
rect 131 12 133 25
rect 139 12 141 25
rect 147 12 149 25
<< ptransistor >>
rect 11 38 13 66
rect 19 38 21 66
rect 27 38 29 66
rect 37 38 39 66
rect 44 38 46 66
rect 54 38 56 66
rect 75 38 77 66
rect 104 38 106 66
rect 114 38 116 66
rect 121 38 123 66
rect 131 38 133 66
rect 139 38 141 66
rect 147 38 149 66
<< polycontact >>
rect 87 39 91 43
rect 160 40 164 44
rect 3 30 7 34
rect 18 30 22 34
rect 35 30 39 34
rect 47 23 51 27
rect 63 30 67 34
rect 93 29 97 33
rect 122 30 126 34
rect 138 30 142 34
rect 80 13 84 17
rect 161 14 165 18
<< ndcontact >>
rect 31 21 35 25
rect 4 4 8 8
rect 50 13 54 17
rect 61 15 65 19
rect 72 13 76 17
rect 61 8 65 12
rect 98 13 102 17
rect 108 20 112 24
rect 108 13 112 17
rect 125 14 129 18
rect 153 20 157 24
rect 153 13 157 17
<< pdcontact >>
rect 5 61 9 65
rect 31 46 35 50
rect 48 54 52 58
rect 59 61 63 65
rect 69 61 73 65
rect 98 61 102 65
rect 79 39 83 43
rect 108 39 112 43
rect 125 46 129 50
rect 151 54 155 58
<< psubstratepcontact >>
rect 88 7 92 11
<< nsubstratencontact >>
rect 87 64 91 68
rect 160 64 164 68
<< psubstratepdiff >>
rect 87 11 93 24
rect 87 7 88 11
rect 92 7 93 11
rect 87 6 93 7
<< nsubstratendiff >>
rect 86 68 92 69
rect 86 64 87 68
rect 91 64 92 68
rect 159 68 165 69
rect 86 48 92 64
rect 159 64 160 68
rect 164 64 165 68
rect 159 63 165 64
<< labels >>
rlabel polysilicon 7 32 7 32 6 an
rlabel polycontact 49 25 49 25 6 bn
rlabel polycontact 82 15 82 15 6 cn
rlabel polycontact 89 41 89 41 6 cn
rlabel polysilicon 127 32 127 32 6 cn
rlabel polycontact 162 42 162 42 6 an
rlabel ptransistor 140 39 140 39 6 bn
rlabel metal1 12 32 12 32 6 z
rlabel polycontact 20 32 20 32 6 b
rlabel metal1 28 36 28 36 6 b
rlabel metal1 20 48 20 48 6 z
rlabel metal1 28 48 28 48 6 z
rlabel metal1 5 35 5 35 6 an
rlabel metal1 29 15 29 15 6 an
rlabel metal1 44 32 44 32 6 c
rlabel metal1 52 32 52 32 6 c
rlabel metal1 60 32 60 32 6 c
rlabel metal1 36 40 36 40 6 b
rlabel metal1 44 40 44 40 6 b
rlabel metal1 52 40 52 40 6 b
rlabel metal1 60 40 60 40 6 b
rlabel metal1 36 48 36 48 6 z
rlabel metal1 44 48 44 48 6 z
rlabel metal1 52 48 52 48 6 z
rlabel metal1 60 48 60 48 6 z
rlabel metal1 84 4 84 4 6 vss
rlabel metal1 78 15 78 15 6 cn
rlabel metal1 67 24 67 24 6 bn
rlabel metal1 76 32 76 32 6 b
rlabel metal1 84 32 84 32 6 b
rlabel metal1 92 32 92 32 6 b
rlabel metal1 68 40 68 40 6 b
rlabel metal1 68 48 68 48 6 z
rlabel metal1 76 48 76 48 6 z
rlabel metal1 84 48 84 48 6 z
rlabel metal1 92 48 92 48 6 z
rlabel metal1 84 68 84 68 6 vdd
rlabel metal1 132 16 132 16 6 z
rlabel metal1 110 19 110 19 6 bn
rlabel metal1 113 32 113 32 6 cn
rlabel metal1 120 40 120 40 6 bn
rlabel metal1 91 41 91 41 6 cn
rlabel metal1 100 48 100 48 6 z
rlabel metal1 108 48 108 48 6 z
rlabel metal1 116 48 116 48 6 z
rlabel metal1 124 48 124 48 6 z
rlabel metal1 132 48 132 48 6 z
rlabel metal1 140 16 140 16 6 z
rlabel metal1 164 24 164 24 6 a
rlabel metal1 148 28 148 28 6 z
rlabel metal1 156 32 156 32 6 a
rlabel metal1 136 32 136 32 6 bn
rlabel metal1 140 40 140 40 6 z
rlabel metal1 162 44 162 44 6 an
rlabel metal1 75 56 75 56 6 an
<< end >>
