magic
tech scmos
timestamp 1179385731
<< checkpaint >>
rect -22 -22 86 94
<< ab >>
rect 0 0 64 72
<< pwell >>
rect -4 -4 68 32
<< nwell >>
rect -4 32 68 76
<< polysilicon >>
rect 12 65 14 70
rect 22 65 24 70
rect 29 65 31 70
rect 39 65 41 70
rect 49 65 51 70
rect 12 35 14 38
rect 22 35 24 38
rect 9 34 24 35
rect 9 30 10 34
rect 14 30 24 34
rect 29 32 31 38
rect 39 35 41 38
rect 49 35 51 38
rect 9 29 24 30
rect 28 29 31 32
rect 35 34 41 35
rect 35 30 36 34
rect 40 30 41 34
rect 35 29 41 30
rect 48 34 55 35
rect 48 30 50 34
rect 54 30 55 34
rect 48 29 55 30
rect 9 24 11 29
rect 21 26 23 29
rect 28 26 30 29
rect 38 26 40 29
rect 48 26 50 29
rect 9 7 11 12
rect 21 9 23 14
rect 28 5 30 14
rect 38 9 40 14
rect 48 5 50 14
rect 28 3 50 5
<< ndiffusion >>
rect 13 24 21 26
rect 4 18 9 24
rect 2 17 9 18
rect 2 13 3 17
rect 7 13 9 17
rect 2 12 9 13
rect 11 14 21 24
rect 23 14 28 26
rect 30 25 38 26
rect 30 21 32 25
rect 36 21 38 25
rect 30 14 38 21
rect 40 19 48 26
rect 40 15 42 19
rect 46 15 48 19
rect 40 14 48 15
rect 50 19 58 26
rect 50 15 52 19
rect 56 15 58 19
rect 50 14 58 15
rect 11 12 19 14
rect 13 8 19 12
rect 13 4 14 8
rect 18 4 19 8
rect 13 3 19 4
<< pdiffusion >>
rect 7 59 12 65
rect 5 58 12 59
rect 5 54 6 58
rect 10 54 12 58
rect 5 51 12 54
rect 5 47 6 51
rect 10 47 12 51
rect 5 46 12 47
rect 7 38 12 46
rect 14 64 22 65
rect 14 60 16 64
rect 20 60 22 64
rect 14 57 22 60
rect 14 53 16 57
rect 20 53 22 57
rect 14 38 22 53
rect 24 38 29 65
rect 31 50 39 65
rect 31 46 33 50
rect 37 46 39 50
rect 31 43 39 46
rect 31 39 33 43
rect 37 39 39 43
rect 31 38 39 39
rect 41 59 49 65
rect 41 55 43 59
rect 47 55 49 59
rect 41 38 49 55
rect 51 64 58 65
rect 51 60 53 64
rect 57 60 58 64
rect 51 56 58 60
rect 51 52 53 56
rect 57 52 58 56
rect 51 38 58 52
<< metal1 >>
rect -2 64 66 72
rect 15 60 16 64
rect 20 60 21 64
rect 6 58 10 59
rect 6 51 10 54
rect 15 57 21 60
rect 15 53 16 57
rect 20 53 21 57
rect 24 55 43 59
rect 47 55 48 59
rect 53 56 57 60
rect 24 50 28 55
rect 53 51 57 52
rect 10 47 28 50
rect 6 46 28 47
rect 33 50 38 51
rect 37 46 38 50
rect 33 43 38 46
rect 2 35 6 43
rect 18 39 33 42
rect 37 39 38 43
rect 18 38 38 39
rect 42 43 46 51
rect 42 38 55 43
rect 2 34 14 35
rect 2 30 10 34
rect 2 29 14 30
rect 18 26 22 38
rect 49 34 55 38
rect 33 30 36 34
rect 40 30 45 34
rect 49 30 50 34
rect 54 30 55 34
rect 41 26 45 30
rect 18 25 37 26
rect 18 21 32 25
rect 36 21 37 25
rect 41 22 55 26
rect 41 17 42 19
rect 2 13 3 17
rect 7 15 42 17
rect 46 15 47 19
rect 7 13 47 15
rect 51 15 52 19
rect 56 15 57 19
rect 51 8 57 15
rect -2 4 14 8
rect 18 4 66 8
rect -2 0 66 4
<< ntransistor >>
rect 9 12 11 24
rect 21 14 23 26
rect 28 14 30 26
rect 38 14 40 26
rect 48 14 50 26
<< ptransistor >>
rect 12 38 14 65
rect 22 38 24 65
rect 29 38 31 65
rect 39 38 41 65
rect 49 38 51 65
<< polycontact >>
rect 10 30 14 34
rect 36 30 40 34
rect 50 30 54 34
<< ndcontact >>
rect 3 13 7 17
rect 32 21 36 25
rect 42 15 46 19
rect 52 15 56 19
rect 14 4 18 8
<< pdcontact >>
rect 6 54 10 58
rect 6 47 10 51
rect 16 60 20 64
rect 16 53 20 57
rect 33 46 37 50
rect 33 39 37 43
rect 43 55 47 59
rect 53 60 57 64
rect 53 52 57 56
<< labels >>
rlabel polycontact 12 32 12 32 6 a
rlabel metal1 4 36 4 36 6 a
rlabel metal1 8 52 8 52 6 n1
rlabel metal1 28 24 28 24 6 z
rlabel metal1 20 28 20 28 6 z
rlabel metal1 28 40 28 40 6 z
rlabel metal1 32 4 32 4 6 vss
rlabel metal1 24 15 24 15 6 n3
rlabel ndcontact 44 16 44 16 6 n3
rlabel metal1 36 32 36 32 6 c
rlabel metal1 44 24 44 24 6 c
rlabel pdcontact 36 48 36 48 6 z
rlabel metal1 44 48 44 48 6 b
rlabel metal1 36 57 36 57 6 n1
rlabel metal1 32 68 32 68 6 vdd
rlabel metal1 52 24 52 24 6 c
rlabel metal1 52 36 52 36 6 b
<< end >>
