magic
tech scmos
timestamp 1179386249
<< checkpaint >>
rect -22 -22 86 94
<< ab >>
rect 0 0 64 72
<< pwell >>
rect -4 -4 68 32
<< nwell >>
rect -4 32 68 76
<< polysilicon >>
rect 9 56 11 60
rect 19 58 21 63
rect 29 58 31 63
rect 39 60 41 64
rect 49 60 51 65
rect 9 34 11 40
rect 19 35 21 40
rect 29 35 31 40
rect 19 34 31 35
rect 9 33 15 34
rect 9 29 10 33
rect 14 29 15 33
rect 9 28 15 29
rect 19 30 26 34
rect 30 30 31 34
rect 19 29 31 30
rect 12 25 14 28
rect 19 25 21 29
rect 29 18 31 29
rect 39 27 41 40
rect 49 35 51 38
rect 45 34 51 35
rect 45 30 46 34
rect 50 30 51 34
rect 45 29 51 30
rect 35 26 41 27
rect 49 26 51 29
rect 35 22 36 26
rect 40 22 41 26
rect 35 21 41 22
rect 36 18 38 21
rect 49 11 51 15
rect 12 2 14 6
rect 19 2 21 6
rect 29 2 31 7
rect 36 2 38 7
<< ndiffusion >>
rect 4 11 12 25
rect 4 7 6 11
rect 10 7 12 11
rect 4 6 12 7
rect 14 6 19 25
rect 21 18 26 25
rect 43 18 49 26
rect 21 17 29 18
rect 21 13 23 17
rect 27 13 29 17
rect 21 7 29 13
rect 31 7 36 18
rect 38 16 49 18
rect 38 12 42 16
rect 46 15 49 16
rect 51 25 58 26
rect 51 21 53 25
rect 57 21 58 25
rect 51 20 58 21
rect 51 15 56 20
rect 46 12 47 15
rect 38 7 47 12
rect 21 6 26 7
<< pdiffusion >>
rect 34 58 39 60
rect 14 56 19 58
rect 2 55 9 56
rect 2 51 3 55
rect 7 51 9 55
rect 2 40 9 51
rect 11 50 19 56
rect 11 46 13 50
rect 17 46 19 50
rect 11 40 19 46
rect 21 57 29 58
rect 21 53 23 57
rect 27 53 29 57
rect 21 40 29 53
rect 31 57 39 58
rect 31 53 33 57
rect 37 53 39 57
rect 31 50 39 53
rect 31 46 33 50
rect 37 46 39 50
rect 31 40 39 46
rect 41 57 49 60
rect 41 53 43 57
rect 47 53 49 57
rect 41 50 49 53
rect 41 46 43 50
rect 47 46 49 50
rect 41 40 49 46
rect 43 38 49 40
rect 51 51 56 60
rect 51 50 58 51
rect 51 46 53 50
rect 57 46 58 50
rect 51 43 58 46
rect 51 39 53 43
rect 57 39 58 43
rect 51 38 58 39
<< metal1 >>
rect -2 68 66 72
rect -2 64 6 68
rect 10 64 66 68
rect 3 55 7 64
rect 22 57 28 64
rect 22 53 23 57
rect 27 53 28 57
rect 33 57 38 59
rect 37 53 38 57
rect 3 50 7 51
rect 33 50 38 53
rect 10 46 13 50
rect 17 46 33 50
rect 37 46 38 50
rect 42 57 48 64
rect 42 53 43 57
rect 47 53 48 57
rect 42 50 48 53
rect 42 46 43 50
rect 47 46 48 50
rect 53 50 57 51
rect 10 43 14 46
rect 2 39 14 43
rect 53 43 57 46
rect 2 18 6 39
rect 17 38 30 42
rect 26 34 30 38
rect 41 35 47 42
rect 10 33 14 34
rect 26 29 30 30
rect 34 34 50 35
rect 34 30 46 34
rect 34 29 50 30
rect 10 26 14 29
rect 53 26 57 39
rect 10 22 36 26
rect 40 25 57 26
rect 40 22 53 25
rect 53 20 57 21
rect 2 17 28 18
rect 2 14 23 17
rect 22 13 23 14
rect 27 13 28 17
rect 42 16 46 17
rect 5 8 6 11
rect -2 7 6 8
rect 10 8 11 11
rect 42 8 46 12
rect 10 7 52 8
rect -2 4 52 7
rect 56 4 66 8
rect -2 0 66 4
<< ntransistor >>
rect 12 6 14 25
rect 19 6 21 25
rect 29 7 31 18
rect 36 7 38 18
rect 49 15 51 26
<< ptransistor >>
rect 9 40 11 56
rect 19 40 21 58
rect 29 40 31 58
rect 39 40 41 60
rect 49 38 51 60
<< polycontact >>
rect 10 29 14 33
rect 26 30 30 34
rect 46 30 50 34
rect 36 22 40 26
<< ndcontact >>
rect 6 7 10 11
rect 23 13 27 17
rect 42 12 46 16
rect 53 21 57 25
<< pdcontact >>
rect 3 51 7 55
rect 13 46 17 50
rect 23 53 27 57
rect 33 53 37 57
rect 33 46 37 50
rect 43 53 47 57
rect 43 46 47 50
rect 53 46 57 50
rect 53 39 57 43
<< psubstratepcontact >>
rect 52 4 56 8
<< nsubstratencontact >>
rect 6 64 10 68
<< psubstratepdiff >>
rect 51 8 57 9
rect 51 4 52 8
rect 56 4 57 8
rect 51 3 57 4
<< nsubstratendiff >>
rect 3 68 13 69
rect 3 64 6 68
rect 10 64 13 68
rect 3 63 13 64
<< labels >>
rlabel ntransistor 13 18 13 18 6 an
rlabel polycontact 38 24 38 24 6 an
rlabel metal1 12 16 12 16 6 z
rlabel metal1 12 28 12 28 6 an
rlabel metal1 4 32 4 32 6 z
rlabel metal1 20 16 20 16 6 z
rlabel polycontact 28 32 28 32 6 b
rlabel metal1 20 40 20 40 6 b
rlabel metal1 20 48 20 48 6 z
rlabel metal1 28 48 28 48 6 z
rlabel metal1 32 4 32 4 6 vss
rlabel metal1 36 32 36 32 6 a
rlabel metal1 44 36 44 36 6 a
rlabel pdcontact 36 56 36 56 6 z
rlabel metal1 32 68 32 68 6 vdd
rlabel metal1 33 24 33 24 6 an
rlabel metal1 55 35 55 35 6 an
<< end >>
