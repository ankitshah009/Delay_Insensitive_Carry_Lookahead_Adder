magic
tech scmos
timestamp 1179385032
<< checkpaint >>
rect -22 -22 62 94
<< ab >>
rect 0 0 40 72
<< pwell >>
rect -4 -4 44 32
<< nwell >>
rect -4 32 44 76
<< polysilicon >>
rect 9 66 11 70
rect 20 54 22 59
rect 30 54 32 59
rect 9 35 11 38
rect 20 35 22 46
rect 30 43 32 46
rect 29 42 35 43
rect 29 38 30 42
rect 34 38 35 42
rect 29 37 35 38
rect 9 34 15 35
rect 9 30 10 34
rect 14 30 15 34
rect 9 29 15 30
rect 19 34 25 35
rect 19 30 20 34
rect 24 30 25 34
rect 19 29 25 30
rect 9 26 11 29
rect 22 21 24 29
rect 29 21 31 37
rect 9 7 11 12
rect 22 9 24 14
rect 29 9 31 14
<< ndiffusion >>
rect 2 25 9 26
rect 2 21 3 25
rect 7 21 9 25
rect 2 17 9 21
rect 2 13 3 17
rect 7 13 9 17
rect 2 12 9 13
rect 11 21 19 26
rect 11 14 22 21
rect 24 14 29 21
rect 31 19 38 21
rect 31 15 33 19
rect 37 15 38 19
rect 31 14 38 15
rect 11 12 19 14
rect 13 8 19 12
rect 13 4 14 8
rect 18 4 19 8
rect 13 3 19 4
<< pdiffusion >>
rect 4 51 9 66
rect 2 50 9 51
rect 2 46 3 50
rect 7 46 9 50
rect 2 43 9 46
rect 2 39 3 43
rect 7 39 9 43
rect 2 38 9 39
rect 11 65 18 66
rect 11 61 13 65
rect 17 61 18 65
rect 32 66 38 67
rect 32 62 33 66
rect 37 62 38 66
rect 32 61 38 62
rect 11 58 18 61
rect 11 54 13 58
rect 17 54 18 58
rect 34 54 38 61
rect 11 46 20 54
rect 22 51 30 54
rect 22 47 24 51
rect 28 47 30 51
rect 22 46 30 47
rect 32 46 38 54
rect 11 38 18 46
<< metal1 >>
rect -2 68 42 72
rect -2 65 23 68
rect -2 64 13 65
rect 12 61 13 64
rect 17 64 23 65
rect 27 66 42 68
rect 27 64 33 66
rect 17 61 18 64
rect 32 62 33 64
rect 37 64 42 66
rect 37 62 38 64
rect 12 58 18 61
rect 12 54 13 58
rect 17 54 18 58
rect 2 50 7 51
rect 2 46 3 50
rect 2 43 7 46
rect 2 39 3 43
rect 2 38 7 39
rect 10 47 24 51
rect 28 47 29 51
rect 2 26 6 38
rect 10 34 14 47
rect 25 38 30 42
rect 34 38 38 51
rect 17 30 20 34
rect 24 30 31 34
rect 10 26 14 30
rect 2 25 7 26
rect 2 21 3 25
rect 10 22 22 26
rect 25 22 31 30
rect 2 19 7 21
rect 18 19 22 22
rect 2 17 14 19
rect 2 13 3 17
rect 7 13 14 17
rect 18 15 33 19
rect 37 15 38 19
rect -2 4 14 8
rect 18 4 42 8
rect -2 0 42 4
<< ntransistor >>
rect 9 12 11 26
rect 22 14 24 21
rect 29 14 31 21
<< ptransistor >>
rect 9 38 11 66
rect 20 46 22 54
rect 30 46 32 54
<< polycontact >>
rect 30 38 34 42
rect 10 30 14 34
rect 20 30 24 34
<< ndcontact >>
rect 3 21 7 25
rect 3 13 7 17
rect 33 15 37 19
rect 14 4 18 8
<< pdcontact >>
rect 3 46 7 50
rect 3 39 7 43
rect 13 61 17 65
rect 33 62 37 66
rect 13 54 17 58
rect 24 47 28 51
<< nsubstratencontact >>
rect 23 64 27 68
<< nsubstratendiff >>
rect 22 68 28 69
rect 22 64 23 68
rect 27 64 28 68
rect 22 61 28 64
<< labels >>
rlabel polycontact 12 32 12 32 6 zn
rlabel metal1 4 32 4 32 6 z
rlabel metal1 12 16 12 16 6 z
rlabel metal1 12 36 12 36 6 zn
rlabel metal1 20 4 20 4 6 vss
rlabel metal1 20 32 20 32 6 a
rlabel metal1 28 28 28 28 6 a
rlabel metal1 28 40 28 40 6 b
rlabel metal1 19 49 19 49 6 zn
rlabel metal1 20 68 20 68 6 vdd
rlabel metal1 28 17 28 17 6 zn
rlabel metal1 36 48 36 48 6 b
<< end >>
