magic
tech scmos
timestamp 1179387436
<< checkpaint >>
rect -22 -22 102 94
<< ab >>
rect 0 0 80 72
<< pwell >>
rect -4 -4 84 32
<< nwell >>
rect -4 32 84 76
<< polysilicon >>
rect 9 66 11 70
rect 19 66 21 70
rect 29 66 31 70
rect 47 66 49 70
rect 9 35 11 38
rect 19 35 21 38
rect 29 36 31 39
rect 64 60 70 61
rect 64 57 65 60
rect 58 56 65 57
rect 69 56 70 60
rect 58 55 70 56
rect 58 52 60 55
rect 68 52 70 55
rect 29 35 39 36
rect 47 35 49 38
rect 58 35 60 38
rect 68 35 70 38
rect 9 34 15 35
rect 9 30 10 34
rect 14 30 15 34
rect 9 29 15 30
rect 19 34 25 35
rect 29 34 42 35
rect 19 30 20 34
rect 24 30 25 34
rect 36 30 37 34
rect 41 30 42 34
rect 19 29 25 30
rect 13 26 15 29
rect 20 26 22 29
rect 30 26 32 30
rect 36 29 42 30
rect 40 26 42 29
rect 47 34 54 35
rect 47 30 49 34
rect 53 30 54 34
rect 58 33 70 35
rect 47 29 54 30
rect 47 26 49 29
rect 63 26 65 33
rect 13 8 15 13
rect 20 8 22 13
rect 40 8 42 12
rect 47 8 49 12
rect 30 4 32 7
rect 63 4 65 13
rect 30 2 65 4
<< ndiffusion >>
rect 4 13 13 26
rect 15 13 20 26
rect 22 18 30 26
rect 22 14 24 18
rect 28 14 30 18
rect 22 13 30 14
rect 4 8 11 13
rect 4 4 6 8
rect 10 4 11 8
rect 25 7 30 13
rect 32 23 40 26
rect 32 19 34 23
rect 38 19 40 23
rect 32 12 40 19
rect 42 12 47 26
rect 49 18 63 26
rect 49 14 57 18
rect 61 14 63 18
rect 49 13 63 14
rect 65 25 72 26
rect 65 21 67 25
rect 71 21 72 25
rect 65 20 72 21
rect 65 13 70 20
rect 49 12 61 13
rect 32 7 37 12
rect 4 3 11 4
<< pdiffusion >>
rect 4 59 9 66
rect 2 58 9 59
rect 2 54 3 58
rect 7 54 9 58
rect 2 53 9 54
rect 4 38 9 53
rect 11 50 19 66
rect 11 46 13 50
rect 17 46 19 50
rect 11 38 19 46
rect 21 50 29 66
rect 21 46 23 50
rect 27 46 29 50
rect 21 39 29 46
rect 31 65 38 66
rect 31 61 33 65
rect 37 61 38 65
rect 31 55 38 61
rect 31 39 36 55
rect 42 51 47 66
rect 40 50 47 51
rect 40 46 41 50
rect 45 46 47 50
rect 40 45 47 46
rect 21 38 26 39
rect 42 38 47 45
rect 49 65 56 66
rect 49 61 51 65
rect 55 61 56 65
rect 72 68 78 69
rect 72 64 73 68
rect 77 64 78 68
rect 49 52 56 61
rect 72 52 78 64
rect 49 38 58 52
rect 60 50 68 52
rect 60 46 62 50
rect 66 46 68 50
rect 60 43 68 46
rect 60 39 62 43
rect 66 39 68 43
rect 60 38 68 39
rect 70 38 78 52
<< metal1 >>
rect -2 68 82 72
rect -2 65 62 68
rect -2 64 33 65
rect 32 61 33 64
rect 37 64 51 65
rect 37 61 38 64
rect 50 61 51 64
rect 55 64 62 65
rect 66 64 73 68
rect 77 64 82 68
rect 55 61 56 64
rect 2 54 3 58
rect 7 54 54 58
rect 64 56 65 60
rect 69 59 70 60
rect 69 56 78 59
rect 64 54 78 56
rect 2 50 17 51
rect 2 46 13 50
rect 2 45 17 46
rect 20 46 23 50
rect 27 46 41 50
rect 45 46 46 50
rect 2 18 6 45
rect 20 42 24 46
rect 50 43 54 54
rect 61 46 62 50
rect 66 46 67 50
rect 61 43 67 46
rect 10 38 24 42
rect 27 39 62 43
rect 66 39 71 43
rect 10 34 14 38
rect 27 34 31 39
rect 19 30 20 34
rect 24 30 31 34
rect 34 34 46 35
rect 34 30 37 34
rect 41 30 46 34
rect 10 26 14 30
rect 34 29 46 30
rect 49 34 54 35
rect 53 30 54 34
rect 49 29 54 30
rect 10 23 38 26
rect 10 22 34 23
rect 34 18 38 19
rect 2 14 24 18
rect 28 14 31 18
rect 42 13 46 29
rect 50 26 54 29
rect 50 22 63 26
rect 67 25 71 39
rect 74 37 78 54
rect 50 13 54 22
rect 67 20 71 21
rect 57 18 61 19
rect 57 8 61 14
rect -2 4 6 8
rect 10 4 72 8
rect 76 4 82 8
rect -2 0 82 4
<< ntransistor >>
rect 13 13 15 26
rect 20 13 22 26
rect 30 7 32 26
rect 40 12 42 26
rect 47 12 49 26
rect 63 13 65 26
<< ptransistor >>
rect 9 38 11 66
rect 19 38 21 66
rect 29 39 31 66
rect 47 38 49 66
rect 58 38 60 52
rect 68 38 70 52
<< polycontact >>
rect 65 56 69 60
rect 10 30 14 34
rect 20 30 24 34
rect 37 30 41 34
rect 49 30 53 34
<< ndcontact >>
rect 24 14 28 18
rect 6 4 10 8
rect 34 19 38 23
rect 57 14 61 18
rect 67 21 71 25
<< pdcontact >>
rect 3 54 7 58
rect 13 46 17 50
rect 23 46 27 50
rect 33 61 37 65
rect 41 46 45 50
rect 51 61 55 65
rect 73 64 77 68
rect 62 46 66 50
rect 62 39 66 43
<< psubstratepcontact >>
rect 72 4 76 8
<< nsubstratencontact >>
rect 62 64 66 68
<< psubstratepdiff >>
rect 71 8 77 9
rect 71 4 72 8
rect 76 4 77 8
rect 71 3 77 4
<< nsubstratendiff >>
rect 60 68 68 69
rect 60 64 62 68
rect 66 64 68 68
rect 60 63 68 64
<< labels >>
rlabel polycontact 12 32 12 32 6 an
rlabel polycontact 22 32 22 32 6 bn
rlabel metal1 12 16 12 16 6 z
rlabel metal1 4 36 4 36 6 z
rlabel polycontact 12 32 12 32 6 an
rlabel metal1 12 48 12 48 6 z
rlabel metal1 28 16 28 16 6 z
rlabel metal1 20 16 20 16 6 z
rlabel metal1 24 24 24 24 6 an
rlabel metal1 25 32 25 32 6 bn
rlabel metal1 36 32 36 32 6 a2
rlabel metal1 40 4 40 4 6 vss
rlabel metal1 44 24 44 24 6 a2
rlabel metal1 52 24 52 24 6 a1
rlabel metal1 33 48 33 48 6 an
rlabel metal1 28 56 28 56 6 bn
rlabel metal1 40 68 40 68 6 vdd
rlabel metal1 60 24 60 24 6 a1
rlabel metal1 69 31 69 31 6 bn
rlabel metal1 64 44 64 44 6 bn
rlabel metal1 49 41 49 41 6 bn
rlabel metal1 76 48 76 48 6 b
rlabel metal1 68 56 68 56 6 b
<< end >>
