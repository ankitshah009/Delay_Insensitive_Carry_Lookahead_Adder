magic
tech scmos
timestamp 1179387689
<< checkpaint >>
rect -22 -25 94 105
<< ab >>
rect 0 0 72 80
<< pwell >>
rect -4 -7 76 36
<< nwell >>
rect -4 36 76 87
<< polysilicon >>
rect 6 72 30 74
rect 6 63 8 72
rect 18 64 20 68
rect 28 64 30 72
rect 38 72 60 74
rect 38 64 40 72
rect 48 64 50 68
rect 58 64 60 72
rect 2 62 8 63
rect 2 58 3 62
rect 7 58 8 62
rect 2 57 8 58
rect 18 39 20 42
rect 8 38 20 39
rect 8 34 9 38
rect 13 37 20 38
rect 28 37 30 42
rect 38 38 40 42
rect 48 38 50 42
rect 58 39 60 42
rect 58 38 64 39
rect 48 37 54 38
rect 13 34 14 37
rect 28 35 34 37
rect 8 33 14 34
rect 12 30 14 33
rect 22 29 24 33
rect 32 29 34 35
rect 48 34 49 37
rect 42 33 49 34
rect 53 33 54 37
rect 58 34 59 38
rect 63 34 64 38
rect 58 33 64 34
rect 42 32 54 33
rect 42 29 44 32
rect 61 29 63 33
rect 12 14 14 19
rect 22 10 24 18
rect 32 14 34 18
rect 42 14 44 18
rect 61 10 63 18
rect 22 8 63 10
<< ndiffusion >>
rect 2 24 12 30
rect 2 20 3 24
rect 7 20 12 24
rect 2 19 12 20
rect 14 29 19 30
rect 14 27 22 29
rect 14 23 16 27
rect 20 23 22 27
rect 14 19 22 23
rect 17 18 22 19
rect 24 28 32 29
rect 24 24 26 28
rect 30 24 32 28
rect 24 18 32 24
rect 34 28 42 29
rect 34 24 36 28
rect 40 24 42 28
rect 34 18 42 24
rect 44 23 61 29
rect 44 19 55 23
rect 59 19 61 23
rect 44 18 61 19
rect 63 28 70 29
rect 63 24 65 28
rect 69 24 70 28
rect 63 23 70 24
rect 63 18 68 23
<< pdiffusion >>
rect 11 63 18 64
rect 11 59 12 63
rect 16 59 18 63
rect 11 42 18 59
rect 20 47 28 64
rect 20 43 22 47
rect 26 43 28 47
rect 20 42 28 43
rect 30 47 38 64
rect 30 43 32 47
rect 36 43 38 47
rect 30 42 38 43
rect 40 47 48 64
rect 40 43 42 47
rect 46 43 48 47
rect 40 42 48 43
rect 50 63 58 64
rect 50 59 52 63
rect 56 59 58 63
rect 50 42 58 59
rect 60 56 65 64
rect 60 55 67 56
rect 60 51 62 55
rect 66 51 67 55
rect 60 50 67 51
rect 60 42 65 50
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect -2 68 74 78
rect 11 63 17 68
rect 3 62 7 63
rect 11 59 12 63
rect 16 59 17 63
rect 51 63 57 68
rect 51 59 52 63
rect 56 59 57 63
rect 3 55 7 58
rect 3 51 62 55
rect 42 47 46 48
rect 2 39 6 47
rect 17 43 22 47
rect 26 43 27 47
rect 30 43 32 47
rect 36 43 38 47
rect 2 38 14 39
rect 2 34 9 38
rect 13 34 14 38
rect 2 33 14 34
rect 17 28 21 43
rect 30 41 38 43
rect 30 38 34 41
rect 42 38 46 43
rect 50 41 62 47
rect 58 39 62 41
rect 58 38 63 39
rect 16 27 21 28
rect 3 24 7 25
rect 20 23 21 27
rect 25 34 34 38
rect 38 34 46 38
rect 49 37 53 38
rect 25 28 31 34
rect 38 28 42 34
rect 58 34 59 38
rect 58 33 63 34
rect 49 31 53 33
rect 25 24 26 28
rect 30 24 31 28
rect 35 24 36 28
rect 40 24 42 28
rect 47 27 53 31
rect 66 29 70 55
rect 65 28 70 29
rect 16 22 21 23
rect 3 12 7 20
rect 17 21 21 22
rect 47 21 51 27
rect 69 24 70 28
rect 17 17 51 21
rect 55 23 59 24
rect 65 23 70 24
rect 55 12 59 19
rect -2 2 74 12
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
<< ntransistor >>
rect 12 19 14 30
rect 22 18 24 29
rect 32 18 34 29
rect 42 18 44 29
rect 61 18 63 29
<< ptransistor >>
rect 18 42 20 64
rect 28 42 30 64
rect 38 42 40 64
rect 48 42 50 64
rect 58 42 60 64
<< polycontact >>
rect 3 58 7 62
rect 9 34 13 38
rect 49 33 53 37
rect 59 34 63 38
<< ndcontact >>
rect 3 20 7 24
rect 16 23 20 27
rect 26 24 30 28
rect 36 24 40 28
rect 55 19 59 23
rect 65 24 69 28
<< pdcontact >>
rect 12 59 16 63
rect 22 43 26 47
rect 32 43 36 47
rect 42 43 46 47
rect 52 59 56 63
rect 62 51 66 55
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
<< psubstratepdiff >>
rect 0 2 72 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 72 2
rect 0 -3 72 -2
<< nsubstratendiff >>
rect 0 82 72 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 72 82
rect 0 77 72 78
<< labels >>
rlabel polycontact 5 60 5 60 6 bn
rlabel polycontact 51 35 51 35 6 an
rlabel metal1 4 40 4 40 6 a
rlabel metal1 5 57 5 57 6 bn
rlabel metal1 19 32 19 32 6 an
rlabel polycontact 12 36 12 36 6 a
rlabel metal1 22 45 22 45 6 an
rlabel metal1 36 6 36 6 6 vss
rlabel metal1 40 31 40 31 6 ai
rlabel metal1 28 32 28 32 6 z
rlabel metal1 36 44 36 44 6 z
rlabel metal1 36 74 36 74 6 vdd
rlabel metal1 51 32 51 32 6 an
rlabel metal1 52 44 52 44 6 b
rlabel metal1 44 41 44 41 6 ai
rlabel metal1 60 40 60 40 6 b
rlabel metal1 68 39 68 39 6 bn
rlabel metal1 36 53 36 53 6 bn
<< end >>
