magic
tech scmos
timestamp 1185039072
<< checkpaint >>
rect -22 -24 112 124
<< ab >>
rect 0 0 90 100
<< pwell >>
rect -2 -4 92 49
<< nwell >>
rect -2 49 92 104
<< polysilicon >>
rect 45 95 47 98
rect 57 95 59 98
rect 67 95 69 98
rect 77 95 79 98
rect 11 85 13 88
rect 23 85 25 88
rect 33 85 35 88
rect 11 43 13 55
rect 23 53 25 55
rect 33 53 35 55
rect 45 53 47 55
rect 21 51 25 53
rect 31 51 35 53
rect 43 51 47 53
rect 57 53 59 55
rect 67 53 69 55
rect 57 52 63 53
rect 21 43 23 51
rect 31 43 33 51
rect 43 43 45 51
rect 57 49 58 52
rect 7 42 13 43
rect 7 38 8 42
rect 12 38 13 42
rect 7 37 13 38
rect 17 42 23 43
rect 17 38 18 42
rect 22 38 23 42
rect 17 37 23 38
rect 27 42 33 43
rect 27 38 28 42
rect 32 38 33 42
rect 27 37 33 38
rect 37 42 45 43
rect 37 38 38 42
rect 42 38 45 42
rect 37 37 45 38
rect 11 35 13 37
rect 21 35 23 37
rect 31 35 33 37
rect 43 35 45 37
rect 55 48 58 49
rect 62 48 63 52
rect 55 47 63 48
rect 67 52 73 53
rect 67 48 68 52
rect 72 48 73 52
rect 67 47 73 48
rect 55 35 57 47
rect 67 39 69 47
rect 65 37 69 39
rect 77 43 79 55
rect 77 42 83 43
rect 77 38 78 42
rect 82 38 83 42
rect 77 37 83 38
rect 65 35 67 37
rect 77 35 79 37
rect 43 14 45 17
rect 55 14 57 17
rect 65 14 67 17
rect 77 14 79 17
rect 11 8 13 11
rect 21 8 23 11
rect 31 8 33 11
<< ndiffusion >>
rect 3 12 11 35
rect 3 8 4 12
rect 8 11 11 12
rect 13 11 21 35
rect 23 11 31 35
rect 33 22 43 35
rect 33 18 36 22
rect 40 18 43 22
rect 33 17 43 18
rect 45 22 55 35
rect 45 18 48 22
rect 52 18 55 22
rect 45 17 55 18
rect 57 17 65 35
rect 67 22 77 35
rect 67 18 70 22
rect 74 18 77 22
rect 67 17 77 18
rect 79 22 87 35
rect 79 18 82 22
rect 86 18 87 22
rect 79 17 87 18
rect 33 11 40 17
rect 59 11 63 17
rect 8 8 9 11
rect 58 10 64 11
rect 3 7 9 8
rect 58 6 59 10
rect 63 6 64 10
rect 58 5 64 6
<< pdiffusion >>
rect 26 96 32 97
rect 26 92 27 96
rect 31 92 32 96
rect 26 91 32 92
rect 27 85 31 91
rect 41 85 45 95
rect 3 82 11 85
rect 3 78 4 82
rect 8 78 11 82
rect 3 55 11 78
rect 13 82 23 85
rect 13 78 16 82
rect 20 78 23 82
rect 13 55 23 78
rect 25 55 33 85
rect 35 82 45 85
rect 35 78 38 82
rect 42 78 45 82
rect 35 55 45 78
rect 47 72 57 95
rect 47 68 50 72
rect 54 68 57 72
rect 47 55 57 68
rect 59 55 67 95
rect 69 55 77 95
rect 79 82 87 95
rect 79 78 82 82
rect 86 78 87 82
rect 79 55 87 78
<< metal1 >>
rect -2 96 92 101
rect -2 92 7 96
rect 11 92 15 96
rect 19 92 27 96
rect 31 92 92 96
rect -2 87 92 92
rect 3 82 9 87
rect 3 78 4 82
rect 8 78 9 82
rect 3 77 9 78
rect 15 82 21 83
rect 37 82 43 83
rect 81 82 87 83
rect 15 78 16 82
rect 20 78 38 82
rect 42 78 82 82
rect 86 78 87 82
rect 15 77 21 78
rect 37 77 43 78
rect 81 77 87 78
rect 47 72 55 73
rect 7 42 13 72
rect 7 38 8 42
rect 12 38 13 42
rect 7 18 13 38
rect 17 42 23 72
rect 17 38 18 42
rect 22 38 23 42
rect 17 18 23 38
rect 27 42 33 72
rect 27 38 28 42
rect 32 38 33 42
rect 27 28 33 38
rect 37 42 43 72
rect 37 38 38 42
rect 42 38 43 42
rect 37 37 43 38
rect 47 68 50 72
rect 54 68 55 72
rect 47 67 55 68
rect 47 33 53 67
rect 37 27 53 33
rect 57 52 63 62
rect 57 48 58 52
rect 62 48 63 52
rect 57 28 63 48
rect 67 52 73 72
rect 67 48 68 52
rect 72 48 73 52
rect 67 28 73 48
rect 77 42 83 72
rect 77 38 78 42
rect 82 38 83 42
rect 77 28 83 38
rect 37 23 43 27
rect 35 22 43 23
rect 35 18 36 22
rect 40 18 43 22
rect 35 17 43 18
rect 47 22 53 23
rect 69 22 75 23
rect 47 18 48 22
rect 52 18 70 22
rect 74 18 75 22
rect 47 17 53 18
rect 69 17 75 18
rect 81 22 87 23
rect 81 18 82 22
rect 86 18 87 22
rect 81 13 87 18
rect -2 12 92 13
rect -2 8 4 12
rect 8 10 92 12
rect 8 8 59 10
rect -2 6 59 8
rect 63 6 72 10
rect 76 6 80 10
rect 84 6 92 10
rect -2 -1 92 6
<< ntransistor >>
rect 11 11 13 35
rect 21 11 23 35
rect 31 11 33 35
rect 43 17 45 35
rect 55 17 57 35
rect 65 17 67 35
rect 77 17 79 35
<< ptransistor >>
rect 11 55 13 85
rect 23 55 25 85
rect 33 55 35 85
rect 45 55 47 95
rect 57 55 59 95
rect 67 55 69 95
rect 77 55 79 95
<< polycontact >>
rect 8 38 12 42
rect 18 38 22 42
rect 28 38 32 42
rect 38 38 42 42
rect 58 48 62 52
rect 68 48 72 52
rect 78 38 82 42
<< ndcontact >>
rect 4 8 8 12
rect 36 18 40 22
rect 48 18 52 22
rect 70 18 74 22
rect 82 18 86 22
rect 59 6 63 10
<< pdcontact >>
rect 27 92 31 96
rect 4 78 8 82
rect 16 78 20 82
rect 38 78 42 82
rect 50 68 54 72
rect 82 78 86 82
<< psubstratepcontact >>
rect 72 6 76 10
rect 80 6 84 10
<< nsubstratencontact >>
rect 7 92 11 96
rect 15 92 19 96
<< psubstratepdiff >>
rect 71 10 85 11
rect 71 6 72 10
rect 76 6 80 10
rect 84 6 85 10
rect 71 5 85 6
<< nsubstratendiff >>
rect 6 96 20 97
rect 6 92 7 96
rect 11 92 15 96
rect 19 92 20 96
rect 6 91 20 92
<< labels >>
rlabel metal1 10 45 10 45 6 i0
rlabel metal1 10 45 10 45 6 i0
rlabel metal1 30 50 30 50 6 i2
rlabel metal1 20 45 20 45 6 i1
rlabel metal1 30 50 30 50 6 i2
rlabel metal1 20 45 20 45 6 i1
rlabel metal1 45 6 45 6 6 vss
rlabel metal1 45 6 45 6 6 vss
rlabel metal1 40 25 40 25 6 nq
rlabel metal1 40 25 40 25 6 nq
rlabel metal1 50 50 50 50 6 nq
rlabel metal1 40 55 40 55 6 i6
rlabel metal1 50 50 50 50 6 nq
rlabel metal1 40 55 40 55 6 i6
rlabel metal1 45 94 45 94 6 vdd
rlabel metal1 45 94 45 94 6 vdd
rlabel polycontact 70 50 70 50 6 i4
rlabel metal1 60 45 60 45 6 i3
rlabel polycontact 70 50 70 50 6 i4
rlabel metal1 60 45 60 45 6 i3
rlabel metal1 80 50 80 50 6 i5
rlabel metal1 80 50 80 50 6 i5
<< end >>
