magic
tech scmos
timestamp 1185038949
<< checkpaint >>
rect -22 -24 102 124
<< ab >>
rect 0 0 80 100
<< pwell >>
rect -2 -4 82 49
<< nwell >>
rect -2 49 82 104
<< polysilicon >>
rect 11 95 13 98
rect 23 95 25 98
rect 35 95 37 98
rect 47 95 49 98
rect 59 95 61 98
rect 11 53 13 55
rect 11 52 19 53
rect 11 48 14 52
rect 18 48 19 52
rect 11 47 19 48
rect 23 43 25 55
rect 35 43 37 55
rect 47 43 49 55
rect 59 43 61 55
rect 3 42 61 43
rect 3 38 4 42
rect 8 38 61 42
rect 3 37 61 38
rect 11 32 19 33
rect 11 28 14 32
rect 18 28 19 32
rect 11 27 19 28
rect 11 25 13 27
rect 23 25 25 37
rect 35 25 37 37
rect 47 25 49 37
rect 59 25 61 37
rect 11 2 13 5
rect 23 2 25 5
rect 35 2 37 5
rect 47 2 49 5
rect 59 2 61 5
<< ndiffusion >>
rect 3 22 11 25
rect 3 18 4 22
rect 8 18 11 22
rect 3 5 11 18
rect 13 12 23 25
rect 13 8 16 12
rect 20 8 23 12
rect 13 5 23 8
rect 25 22 35 25
rect 25 18 28 22
rect 32 18 35 22
rect 25 5 35 18
rect 37 22 47 25
rect 37 18 40 22
rect 44 18 47 22
rect 37 12 47 18
rect 37 8 40 12
rect 44 8 47 12
rect 37 5 47 8
rect 49 22 59 25
rect 49 18 52 22
rect 56 18 59 22
rect 49 5 59 18
rect 61 22 69 25
rect 61 18 64 22
rect 68 18 69 22
rect 61 12 69 18
rect 61 8 64 12
rect 68 8 69 12
rect 61 5 69 8
<< pdiffusion >>
rect 3 82 11 95
rect 3 78 4 82
rect 8 78 11 82
rect 3 72 11 78
rect 3 68 4 72
rect 8 68 11 72
rect 3 62 11 68
rect 3 58 4 62
rect 8 58 11 62
rect 3 55 11 58
rect 13 92 23 95
rect 13 88 16 92
rect 20 88 23 92
rect 13 55 23 88
rect 25 82 35 95
rect 25 78 28 82
rect 32 78 35 82
rect 25 72 35 78
rect 25 68 28 72
rect 32 68 35 72
rect 25 62 35 68
rect 25 58 28 62
rect 32 58 35 62
rect 25 55 35 58
rect 37 92 47 95
rect 37 88 40 92
rect 44 88 47 92
rect 37 82 47 88
rect 37 78 40 82
rect 44 78 47 82
rect 37 72 47 78
rect 37 68 40 72
rect 44 68 47 72
rect 37 62 47 68
rect 37 58 40 62
rect 44 58 47 62
rect 37 55 47 58
rect 49 82 59 95
rect 49 78 52 82
rect 56 78 59 82
rect 49 72 59 78
rect 49 68 52 72
rect 56 68 59 72
rect 49 62 59 68
rect 49 58 52 62
rect 56 58 59 62
rect 49 55 59 58
rect 61 92 69 95
rect 61 88 64 92
rect 68 88 69 92
rect 61 82 69 88
rect 61 78 64 82
rect 68 78 69 82
rect 61 77 69 78
rect 61 55 65 77
<< metal1 >>
rect -2 92 82 101
rect -2 88 16 92
rect 20 88 40 92
rect 44 88 64 92
rect 68 88 82 92
rect -2 87 82 88
rect 3 82 9 83
rect 27 82 33 83
rect 3 78 4 82
rect 8 78 9 82
rect 3 77 9 78
rect 4 73 8 77
rect 3 72 9 73
rect 3 68 4 72
rect 8 68 9 72
rect 3 67 9 68
rect 4 63 8 67
rect 3 62 9 63
rect 3 58 4 62
rect 8 58 9 62
rect 3 57 9 58
rect 4 43 8 57
rect 17 53 23 82
rect 13 52 23 53
rect 13 48 14 52
rect 18 48 23 52
rect 13 47 23 48
rect 3 42 9 43
rect 3 38 4 42
rect 8 38 9 42
rect 3 37 9 38
rect 4 23 8 37
rect 17 33 23 47
rect 13 32 23 33
rect 13 28 14 32
rect 18 28 23 32
rect 13 27 23 28
rect 3 22 9 23
rect 3 18 4 22
rect 8 18 9 22
rect 17 18 23 27
rect 27 78 28 82
rect 32 78 33 82
rect 27 72 33 78
rect 27 68 28 72
rect 32 68 33 72
rect 27 62 33 68
rect 27 58 28 62
rect 32 58 33 62
rect 27 43 33 58
rect 39 82 45 87
rect 39 78 40 82
rect 44 78 45 82
rect 39 72 45 78
rect 39 68 40 72
rect 44 68 45 72
rect 39 62 45 68
rect 39 58 40 62
rect 44 58 45 62
rect 39 57 45 58
rect 51 82 57 83
rect 51 78 52 82
rect 56 78 57 82
rect 51 72 57 78
rect 51 68 52 72
rect 56 68 57 72
rect 51 62 57 68
rect 63 82 69 87
rect 63 78 64 82
rect 68 78 69 82
rect 63 71 69 78
rect 63 70 77 71
rect 63 66 72 70
rect 76 66 77 70
rect 63 65 77 66
rect 51 58 52 62
rect 56 58 57 62
rect 51 43 57 58
rect 71 60 77 65
rect 71 56 72 60
rect 76 56 77 60
rect 71 55 77 56
rect 27 37 57 43
rect 27 22 33 37
rect 27 18 28 22
rect 32 18 33 22
rect 3 17 9 18
rect 27 17 33 18
rect 39 22 45 23
rect 39 18 40 22
rect 44 18 45 22
rect 39 13 45 18
rect 51 22 57 37
rect 51 18 52 22
rect 56 18 57 22
rect 51 17 57 18
rect 63 36 77 37
rect 63 32 64 36
rect 68 32 72 36
rect 76 32 77 36
rect 63 31 77 32
rect 63 22 69 31
rect 63 18 64 22
rect 68 18 69 22
rect 63 13 69 18
rect -2 12 82 13
rect -2 8 16 12
rect 20 8 40 12
rect 44 8 64 12
rect 68 8 82 12
rect -2 -1 82 8
<< ntransistor >>
rect 11 5 13 25
rect 23 5 25 25
rect 35 5 37 25
rect 47 5 49 25
rect 59 5 61 25
<< ptransistor >>
rect 11 55 13 95
rect 23 55 25 95
rect 35 55 37 95
rect 47 55 49 95
rect 59 55 61 95
<< polycontact >>
rect 14 48 18 52
rect 4 38 8 42
rect 14 28 18 32
<< ndcontact >>
rect 4 18 8 22
rect 16 8 20 12
rect 28 18 32 22
rect 40 18 44 22
rect 40 8 44 12
rect 52 18 56 22
rect 64 18 68 22
rect 64 8 68 12
<< pdcontact >>
rect 4 78 8 82
rect 4 68 8 72
rect 4 58 8 62
rect 16 88 20 92
rect 28 78 32 82
rect 28 68 32 72
rect 28 58 32 62
rect 40 88 44 92
rect 40 78 44 82
rect 40 68 44 72
rect 40 58 44 62
rect 52 78 56 82
rect 52 68 56 72
rect 52 58 56 62
rect 64 88 68 92
rect 64 78 68 82
<< psubstratepcontact >>
rect 64 32 68 36
rect 72 32 76 36
<< nsubstratencontact >>
rect 72 66 76 70
rect 72 56 76 60
<< psubstratepdiff >>
rect 63 36 77 37
rect 63 32 64 36
rect 68 32 72 36
rect 76 32 77 36
rect 63 31 77 32
<< nsubstratendiff >>
rect 71 70 77 71
rect 71 66 72 70
rect 76 66 77 70
rect 71 60 77 66
rect 71 56 72 60
rect 76 56 77 60
rect 71 55 77 56
<< labels >>
rlabel metal1 30 50 30 50 6 q
rlabel metal1 30 50 30 50 6 q
rlabel metal1 20 50 20 50 6 i
rlabel metal1 20 50 20 50 6 i
rlabel metal1 40 6 40 6 6 vss
rlabel metal1 40 6 40 6 6 vss
rlabel metal1 40 94 40 94 6 vdd
rlabel metal1 40 94 40 94 6 vdd
<< end >>
