magic
tech scmos
timestamp 1179386040
<< checkpaint >>
rect -22 -22 46 94
<< ab >>
rect 0 0 24 72
<< pwell >>
rect -4 -4 28 32
<< nwell >>
rect -4 32 28 76
<< polysilicon >>
rect 9 66 11 70
rect 9 35 11 38
rect 9 34 15 35
rect 9 30 10 34
rect 14 30 15 34
rect 9 29 15 30
rect 9 26 11 29
rect 9 7 11 12
<< ndiffusion >>
rect 2 24 9 26
rect 2 20 3 24
rect 7 20 9 24
rect 2 17 9 20
rect 2 13 3 17
rect 7 13 9 17
rect 2 12 9 13
rect 11 12 20 26
rect 13 8 20 12
rect 13 4 14 8
rect 18 4 20 8
rect 13 3 20 4
<< pdiffusion >>
rect 13 68 20 69
rect 13 66 14 68
rect 4 53 9 66
rect 2 52 9 53
rect 2 48 3 52
rect 7 48 9 52
rect 2 45 9 48
rect 2 41 3 45
rect 7 41 9 45
rect 2 40 9 41
rect 4 38 9 40
rect 11 64 14 66
rect 18 64 20 68
rect 11 38 20 64
<< metal1 >>
rect -2 68 26 72
rect -2 64 14 68
rect 18 64 26 68
rect 2 53 14 59
rect 2 52 7 53
rect 2 48 3 52
rect 2 45 7 48
rect 2 41 3 45
rect 2 40 7 41
rect 2 25 6 40
rect 18 35 22 59
rect 10 34 22 35
rect 14 30 22 34
rect 10 29 22 30
rect 2 24 7 25
rect 2 20 3 24
rect 2 19 7 20
rect 2 17 14 19
rect 2 13 3 17
rect 7 13 14 17
rect 18 13 22 29
rect -2 4 14 8
rect 18 4 26 8
rect -2 0 26 4
<< ntransistor >>
rect 9 12 11 26
<< ptransistor >>
rect 9 38 11 66
<< polycontact >>
rect 10 30 14 34
<< ndcontact >>
rect 3 20 7 24
rect 3 13 7 17
rect 14 4 18 8
<< pdcontact >>
rect 3 48 7 52
rect 3 41 7 45
rect 14 64 18 68
<< labels >>
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 4 12 4 6 vss
rlabel metal1 12 16 12 16 6 z
rlabel polycontact 12 32 12 32 6 a
rlabel metal1 12 56 12 56 6 z
rlabel metal1 12 68 12 68 6 vdd
rlabel metal1 20 36 20 36 6 a
<< end >>
