.subckt nmx3_x1 cmd0 cmd1 i0 i1 i2 nq vdd vss
*   SPICE3 file   created from nmx3_x1.ext -      technology: scmos
m00 w1     i2     w2     vdd p w=19u  l=2.3636u ad=95p      pd=29.7838u as=114.339p ps=38u
m01 nq     cmd1   w1     vdd p w=18u  l=2.3636u ad=124.364p pd=41.2364u as=90p      ps=28.2162u
m02 w3     cmd1   vdd    vdd p w=14u  l=2.3636u ad=112p     pd=44u      as=123.812p ps=43.3125u
m03 w4     w3     nq     vdd p w=19u  l=2.3636u ad=57p      pd=25u      as=131.273p ps=43.5273u
m04 w2     i1     w4     vdd p w=19u  l=2.3636u ad=114.339p pd=38u      as=57p      ps=25u
m05 vdd    w5     w2     vdd p w=18u  l=2.3636u ad=159.188p pd=55.6875u as=108.321p ps=36u
m06 w6     cmd0   vdd    vdd p w=18u  l=2.3636u ad=54p      pd=24u      as=159.188p ps=55.6875u
m07 nq     i0     w6     vdd p w=18u  l=2.3636u ad=124.364p pd=41.2364u as=54p      ps=24u
m08 w3     cmd1   vss    vss n w=8u   l=2.3636u ad=64p      pd=32u      as=90.8p    ps=35.6u
m09 vdd    cmd0   w5     vdd p w=14u  l=2.3636u ad=123.812p pd=43.3125u as=112p     ps=44u
m10 w7     i2     w8     vss n w=12u  l=2.3636u ad=60p      pd=22u      as=82p      ps=31.3333u
m11 nq     w3     w7     vss n w=12u  l=2.3636u ad=100p     pd=37.3333u as=60p      ps=22u
m12 w9     cmd1   nq     vss n w=12u  l=2.3636u ad=36p      pd=18u      as=100p     ps=37.3333u
m13 w8     i1     w9     vss n w=12u  l=2.3636u ad=82p      pd=31.3333u as=36p      ps=18u
m14 vss    cmd0   w5     vss n w=8u   l=2.3636u ad=90.8p    pd=35.6u    as=64p      ps=32u
m15 vss    cmd0   w8     vss n w=12u  l=2.3636u ad=136.2p   pd=53.4u    as=82p      ps=31.3333u
m16 w10    w5     vss    vss n w=12u  l=2.3636u ad=36p      pd=18u      as=136.2p   ps=53.4u
m17 nq     i0     w10    vss n w=12u  l=2.3636u ad=100p     pd=37.3333u as=36p      ps=18u
C0  i0     i1     0.029f
C1  cmd0   w5     0.315f
C2  vdd    w3     0.046f
C3  w2     cmd1   0.106f
C4  w9     vss    0.004f
C5  w7     w8     0.019f
C6  vss    cmd0   0.017f
C7  nq     w2     0.167f
C8  w4     vdd    0.011f
C9  w8     w5     0.020f
C10 w5     i1     0.130f
C11 i0     cmd1   0.008f
C12 vdd    i2     0.008f
C13 cmd0   w3     0.026f
C14 w8     vss    0.293f
C15 w1     vdd    0.019f
C16 nq     i0     0.175f
C17 w8     w3     0.132f
C18 vss    i1     0.015f
C19 w5     cmd1   0.045f
C20 cmd0   i2     0.012f
C21 i1     w3     0.177f
C22 w8     i2     0.012f
C23 nq     w5     0.315f
C24 vss    cmd1   0.055f
C25 i1     i2     0.057f
C26 w3     cmd1   0.393f
C27 vss    nq     0.176f
C28 vdd    cmd0   0.017f
C29 nq     w3     0.149f
C30 cmd1   i2     0.184f
C31 w2     w3     0.070f
C32 i0     w5     0.309f
C33 vdd    i1     0.017f
C34 nq     i2     0.015f
C35 w10    vss    0.010f
C36 w9     w8     0.012f
C37 w8     cmd0   0.002f
C38 w4     w2     0.012f
C39 w6     vdd    0.011f
C40 vss    i0     0.022f
C41 cmd0   i1     0.077f
C42 i0     w3     0.015f
C43 vdd    cmd1   0.123f
C44 w2     i2     0.010f
C45 w7     vss    0.007f
C46 w8     i1     0.022f
C47 w1     w2     0.019f
C48 nq     vdd    0.266f
C49 vss    w5     0.075f
C50 cmd0   cmd1   0.030f
C51 w5     w3     0.038f
C52 w2     vdd    0.307f
C53 vss    w3     0.043f
C54 w8     cmd1   0.005f
C55 nq     cmd0   0.208f
C56 i1     cmd1   0.151f
C57 w5     i2     0.022f
C58 w8     nq     0.075f
C59 w2     cmd0   0.002f
C60 vdd    i0     0.023f
C61 nq     i1     0.105f
C62 vss    i2     0.008f
C63 w3     i2     0.165f
C64 i0     cmd0   0.345f
C65 vdd    w5     0.013f
C66 nq     cmd1   0.052f
C67 w2     i1     0.022f
C69 nq     vss    0.048f
C71 i0     vss    0.049f
C72 cmd0   vss    0.066f
C73 w5     vss    0.056f
C74 i1     vss    0.038f
C75 w3     vss    0.050f
C76 cmd1   vss    0.071f
C77 i2     vss    0.032f
.ends
