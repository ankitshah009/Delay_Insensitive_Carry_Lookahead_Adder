.subckt nxr2_x4 i0 i1 nq vdd vss
*   SPICE3 file   created from nxr2_x4.ext -      technology: scmos
m00 vdd    i0     w1     vdd p w=20u  l=2.3636u ad=131.2p   pd=39.2u    as=160p     ps=56u
m01 w2     i0     vdd    vdd p w=40u  l=2.3636u ad=200p     pd=50u      as=262.4p   ps=78.4u
m02 w3     w4     w2     vdd p w=40u  l=2.3636u ad=200p     pd=50u      as=200p     ps=50u
m03 w2     w1     w3     vdd p w=40u  l=2.3636u ad=200p     pd=50u      as=200p     ps=50u
m04 vdd    i1     w2     vdd p w=40u  l=2.3636u ad=262.4p   pd=78.4u    as=200p     ps=50u
m05 w4     i1     vdd    vdd p w=20u  l=2.3636u ad=172p     pd=60u      as=131.2p   ps=39.2u
m06 nq     w3     vdd    vdd p w=40u  l=2.3636u ad=200p     pd=50u      as=262.4p   ps=78.4u
m07 vdd    w3     nq     vdd p w=40u  l=2.3636u ad=262.4p   pd=78.4u    as=200p     ps=50u
m08 vss    i0     w1     vss n w=10u  l=2.3636u ad=66.4p    pd=23.2u    as=80p      ps=36u
m09 w5     i0     vss    vss n w=20u  l=2.3636u ad=100p     pd=30u      as=132.8p   ps=46.4u
m10 w3     i1     w5     vss n w=20u  l=2.3636u ad=100p     pd=30u      as=100p     ps=30u
m11 w6     w1     w3     vss n w=20u  l=2.3636u ad=100p     pd=30u      as=100p     ps=30u
m12 vss    w4     w6     vss n w=20u  l=2.3636u ad=132.8p   pd=46.4u    as=100p     ps=30u
m13 w4     i1     vss    vss n w=10u  l=2.3636u ad=140p     pd=56u      as=66.4p    ps=23.2u
m14 nq     w3     vss    vss n w=20u  l=2.3636u ad=100p     pd=30u      as=132.8p   ps=46.4u
m15 vss    w3     nq     vss n w=20u  l=2.3636u ad=132.8p   pd=46.4u    as=100p     ps=30u
C0  i1     i0     0.035f
C1  w2     vdd    0.253f
C2  w1     w4     0.125f
C3  vss    w3     0.471f
C4  w4     i0     0.050f
C5  w1     vdd    0.014f
C6  nq     w2     0.005f
C7  vss    i1     0.082f
C8  i0     vdd    0.096f
C9  vss    w4     0.050f
C10 w3     i1     0.352f
C11 w2     w1     0.005f
C12 w3     w4     0.331f
C13 vss    vdd    0.005f
C14 w5     vss    0.023f
C15 w3     vdd    0.081f
C16 w2     i0     0.039f
C17 i1     w4     0.528f
C18 vss    nq     0.111f
C19 w5     w3     0.019f
C20 i1     vdd    0.130f
C21 w1     i0     0.246f
C22 nq     w3     0.241f
C23 w4     vdd    0.031f
C24 w3     w2     0.155f
C25 nq     i1     0.070f
C26 vss    w1     0.053f
C27 w3     w1     0.085f
C28 w2     i1     0.016f
C29 nq     w4     0.077f
C30 vss    i0     0.060f
C31 w6     vss    0.023f
C32 w3     i0     0.333f
C33 nq     vdd    0.328f
C34 w2     w4     0.027f
C35 i1     w1     0.090f
C36 w6     w3     0.019f
C38 nq     vss    0.018f
C39 w3     vss    0.077f
C40 i1     vss    0.058f
C41 w1     vss    0.050f
C42 w4     vss    0.055f
C43 i0     vss    0.042f
.ends
