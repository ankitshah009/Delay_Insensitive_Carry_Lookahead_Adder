magic
tech scmos
timestamp 1179386302
<< checkpaint >>
rect -22 -22 54 94
<< ab >>
rect 0 0 32 72
<< pwell >>
rect -4 -4 36 32
<< nwell >>
rect -4 32 36 76
<< polysilicon >>
rect 9 66 11 70
rect 19 66 21 70
rect 9 35 11 42
rect 19 39 21 42
rect 19 38 30 39
rect 9 34 15 35
rect 9 30 10 34
rect 14 30 15 34
rect 9 29 15 30
rect 19 34 25 38
rect 29 34 30 38
rect 19 33 30 34
rect 12 26 14 29
rect 19 26 21 33
rect 12 2 14 6
rect 19 2 21 6
<< ndiffusion >>
rect 7 18 12 26
rect 5 17 12 18
rect 5 13 6 17
rect 10 13 12 17
rect 5 12 12 13
rect 7 6 12 12
rect 14 6 19 26
rect 21 18 30 26
rect 21 14 25 18
rect 29 14 30 18
rect 21 11 30 14
rect 21 7 25 11
rect 29 7 30 11
rect 21 6 30 7
<< pdiffusion >>
rect 2 65 9 66
rect 2 61 3 65
rect 7 61 9 65
rect 2 58 9 61
rect 2 54 3 58
rect 7 54 9 58
rect 2 42 9 54
rect 11 58 19 66
rect 11 54 13 58
rect 17 54 19 58
rect 11 51 19 54
rect 11 47 13 51
rect 17 47 19 51
rect 11 42 19 47
rect 21 65 29 66
rect 21 61 23 65
rect 27 61 29 65
rect 21 58 29 61
rect 21 54 23 58
rect 27 54 29 58
rect 21 42 29 54
<< metal1 >>
rect -2 65 34 72
rect -2 64 3 65
rect 2 61 3 64
rect 7 64 23 65
rect 7 61 8 64
rect 2 58 8 61
rect 22 61 23 64
rect 27 64 34 65
rect 27 61 28 64
rect 2 54 3 58
rect 7 54 8 58
rect 13 58 17 59
rect 22 58 28 61
rect 22 54 23 58
rect 27 54 28 58
rect 13 51 17 54
rect 2 47 13 51
rect 2 46 17 47
rect 2 45 14 46
rect 2 13 6 45
rect 18 38 30 43
rect 18 37 25 38
rect 10 34 14 35
rect 29 34 30 38
rect 25 33 30 34
rect 10 27 14 30
rect 26 29 30 33
rect 10 21 22 27
rect 25 18 29 19
rect 10 13 11 17
rect 25 11 29 14
rect -2 7 25 8
rect 29 7 34 8
rect -2 0 34 7
<< ntransistor >>
rect 12 6 14 26
rect 19 6 21 26
<< ptransistor >>
rect 9 42 11 66
rect 19 42 21 66
<< polycontact >>
rect 10 30 14 34
rect 25 34 29 38
<< ndcontact >>
rect 6 13 10 17
rect 25 14 29 18
rect 25 7 29 11
<< pdcontact >>
rect 3 61 7 65
rect 3 54 7 58
rect 13 54 17 58
rect 13 47 17 51
rect 23 61 27 65
rect 23 54 27 58
<< labels >>
rlabel metal1 4 32 4 32 6 z
rlabel metal1 12 28 12 28 6 b
rlabel metal1 12 48 12 48 6 z
rlabel metal1 16 4 16 4 6 vss
rlabel metal1 20 24 20 24 6 b
rlabel metal1 20 40 20 40 6 a
rlabel metal1 16 68 16 68 6 vdd
rlabel polycontact 28 36 28 36 6 a
<< end >>
