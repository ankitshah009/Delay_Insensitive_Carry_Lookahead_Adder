magic
tech scmos
timestamp 1179386595
<< checkpaint >>
rect -22 -22 94 94
<< ab >>
rect 0 0 72 72
<< pwell >>
rect -4 -4 76 32
<< nwell >>
rect -4 32 76 76
<< polysilicon >>
rect 10 68 62 70
rect 10 59 12 68
rect 20 59 22 64
rect 30 59 32 64
rect 40 59 42 64
rect 50 59 52 64
rect 60 59 62 68
rect 10 31 12 39
rect 20 35 22 39
rect 30 35 32 39
rect 40 35 42 39
rect 50 35 52 39
rect 60 35 62 39
rect 20 34 26 35
rect 10 29 16 31
rect 20 30 21 34
rect 25 30 26 34
rect 20 29 26 30
rect 30 34 42 35
rect 30 30 34 34
rect 38 30 42 34
rect 30 29 42 30
rect 46 34 52 35
rect 46 30 47 34
rect 51 30 52 34
rect 46 29 52 30
rect 56 34 63 35
rect 56 30 58 34
rect 62 30 63 34
rect 56 29 63 30
rect 14 26 16 29
rect 22 26 24 29
rect 30 26 32 29
rect 40 26 42 29
rect 48 26 50 29
rect 56 26 58 29
rect 14 2 16 6
rect 22 2 24 6
rect 30 2 32 6
rect 40 2 42 6
rect 48 2 50 6
rect 56 2 58 6
<< ndiffusion >>
rect 6 11 14 26
rect 6 7 8 11
rect 12 7 14 11
rect 6 6 14 7
rect 16 6 22 26
rect 24 6 30 26
rect 32 18 40 26
rect 32 14 34 18
rect 38 14 40 18
rect 32 6 40 14
rect 42 6 48 26
rect 50 6 56 26
rect 58 18 66 26
rect 58 14 60 18
rect 64 14 66 18
rect 58 11 66 14
rect 58 7 60 11
rect 64 7 66 11
rect 58 6 66 7
<< pdiffusion >>
rect 2 58 10 59
rect 2 54 3 58
rect 7 54 10 58
rect 2 51 10 54
rect 2 47 3 51
rect 7 47 10 51
rect 2 39 10 47
rect 12 58 20 59
rect 12 54 14 58
rect 18 54 20 58
rect 12 51 20 54
rect 12 47 14 51
rect 18 47 20 51
rect 12 39 20 47
rect 22 58 30 59
rect 22 54 24 58
rect 28 54 30 58
rect 22 39 30 54
rect 32 58 40 59
rect 32 54 34 58
rect 38 54 40 58
rect 32 51 40 54
rect 32 47 34 51
rect 38 47 40 51
rect 32 39 40 47
rect 42 58 50 59
rect 42 54 44 58
rect 48 54 50 58
rect 42 39 50 54
rect 52 58 60 59
rect 52 54 54 58
rect 58 54 60 58
rect 52 51 60 54
rect 52 47 54 51
rect 58 47 60 51
rect 52 39 60 47
rect 62 58 70 59
rect 62 54 65 58
rect 69 54 70 58
rect 62 39 70 54
<< metal1 >>
rect -2 64 74 72
rect 3 58 7 64
rect 3 51 7 54
rect 14 58 18 59
rect 23 58 29 64
rect 23 54 24 58
rect 28 54 29 58
rect 34 58 38 59
rect 43 58 49 64
rect 43 54 44 58
rect 48 54 49 58
rect 54 58 58 59
rect 64 58 70 64
rect 64 54 65 58
rect 69 54 70 58
rect 14 51 18 54
rect 3 46 7 47
rect 10 47 14 51
rect 34 51 38 54
rect 18 47 34 50
rect 54 51 58 54
rect 38 47 54 50
rect 10 46 58 47
rect 10 18 14 46
rect 22 38 52 42
rect 22 35 26 38
rect 18 34 26 35
rect 46 34 52 38
rect 66 35 70 51
rect 18 30 21 34
rect 25 30 26 34
rect 18 29 26 30
rect 33 30 34 34
rect 38 30 39 34
rect 46 30 47 34
rect 51 30 52 34
rect 58 34 70 35
rect 62 30 70 34
rect 33 26 39 30
rect 58 29 70 30
rect 33 22 47 26
rect 10 14 34 18
rect 38 14 39 18
rect 59 14 60 18
rect 64 14 65 18
rect 59 11 65 14
rect 7 8 8 11
rect -2 7 8 8
rect 12 8 13 11
rect 59 8 60 11
rect 12 7 60 8
rect 64 8 65 11
rect 64 7 74 8
rect -2 0 74 7
<< ntransistor >>
rect 14 6 16 26
rect 22 6 24 26
rect 30 6 32 26
rect 40 6 42 26
rect 48 6 50 26
rect 56 6 58 26
<< ptransistor >>
rect 10 39 12 59
rect 20 39 22 59
rect 30 39 32 59
rect 40 39 42 59
rect 50 39 52 59
rect 60 39 62 59
<< polycontact >>
rect 21 30 25 34
rect 34 30 38 34
rect 47 30 51 34
rect 58 30 62 34
<< ndcontact >>
rect 8 7 12 11
rect 34 14 38 18
rect 60 14 64 18
rect 60 7 64 11
<< pdcontact >>
rect 3 54 7 58
rect 3 47 7 51
rect 14 54 18 58
rect 14 47 18 51
rect 24 54 28 58
rect 34 54 38 58
rect 34 47 38 51
rect 44 54 48 58
rect 54 54 58 58
rect 54 47 58 51
rect 65 54 69 58
<< labels >>
rlabel metal1 20 16 20 16 6 z
rlabel metal1 20 32 20 32 6 b
rlabel metal1 12 36 12 36 6 z
rlabel metal1 20 48 20 48 6 z
rlabel metal1 36 4 36 4 6 vss
rlabel ndcontact 36 16 36 16 6 z
rlabel metal1 28 16 28 16 6 z
rlabel metal1 36 28 36 28 6 c
rlabel metal1 28 40 28 40 6 b
rlabel metal1 36 40 36 40 6 b
rlabel metal1 28 48 28 48 6 z
rlabel metal1 36 52 36 52 6 z
rlabel metal1 36 68 36 68 6 vdd
rlabel metal1 44 24 44 24 6 c
rlabel metal1 44 40 44 40 6 b
rlabel metal1 44 48 44 48 6 z
rlabel metal1 52 48 52 48 6 z
rlabel polycontact 60 32 60 32 6 a
rlabel metal1 68 40 68 40 6 a
<< end >>
