magic
tech scmos
timestamp 1179385977
<< checkpaint >>
rect -22 -25 86 105
<< ab >>
rect 0 0 64 80
<< pwell >>
rect -4 -7 68 36
<< nwell >>
rect -4 36 68 87
<< polysilicon >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 39 70 41 74
rect 49 58 51 63
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 39 39 41 42
rect 9 38 41 39
rect 9 37 36 38
rect 22 34 36 37
rect 40 34 41 38
rect 22 33 41 34
rect 49 39 51 42
rect 49 38 55 39
rect 49 34 50 38
rect 54 34 55 38
rect 49 33 55 34
rect 22 30 24 33
rect 32 30 34 33
rect 22 9 24 14
rect 32 9 34 14
<< ndiffusion >>
rect 14 27 22 30
rect 14 23 16 27
rect 20 23 22 27
rect 14 19 22 23
rect 14 15 16 19
rect 20 15 22 19
rect 14 14 22 15
rect 24 29 32 30
rect 24 25 26 29
rect 30 25 32 29
rect 24 22 32 25
rect 24 18 26 22
rect 30 18 32 22
rect 24 14 32 18
rect 34 27 42 30
rect 34 23 36 27
rect 40 23 42 27
rect 34 19 42 23
rect 34 15 36 19
rect 40 15 42 19
rect 34 14 42 15
<< pdiffusion >>
rect 2 69 9 70
rect 2 65 3 69
rect 7 65 9 69
rect 2 62 9 65
rect 2 58 3 62
rect 7 58 9 62
rect 2 42 9 58
rect 11 54 19 70
rect 11 50 13 54
rect 17 50 19 54
rect 11 47 19 50
rect 11 43 13 47
rect 17 43 19 47
rect 11 42 19 43
rect 21 69 29 70
rect 21 65 23 69
rect 27 65 29 69
rect 21 62 29 65
rect 21 58 23 62
rect 27 58 29 62
rect 21 42 29 58
rect 31 54 39 70
rect 31 50 33 54
rect 37 50 39 54
rect 31 47 39 50
rect 31 43 33 47
rect 37 43 39 47
rect 31 42 39 43
rect 41 58 47 70
rect 41 57 49 58
rect 41 53 43 57
rect 47 53 49 57
rect 41 42 49 53
rect 51 55 56 58
rect 51 54 58 55
rect 51 50 53 54
rect 57 50 58 54
rect 51 47 58 50
rect 51 43 53 47
rect 57 43 58 47
rect 51 42 58 43
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect -2 69 66 78
rect -2 68 3 69
rect 2 65 3 68
rect 7 68 23 69
rect 7 65 8 68
rect 2 62 8 65
rect 2 58 3 62
rect 7 58 8 62
rect 22 65 23 68
rect 27 68 66 69
rect 27 65 28 68
rect 22 62 28 65
rect 22 58 23 62
rect 27 58 28 62
rect 43 57 47 68
rect 13 54 17 55
rect 13 47 17 50
rect 9 43 13 46
rect 33 54 38 55
rect 37 50 38 54
rect 43 52 47 53
rect 53 54 62 55
rect 33 47 38 50
rect 17 43 33 46
rect 37 46 38 47
rect 57 50 62 54
rect 53 49 62 50
rect 53 47 57 49
rect 37 43 53 46
rect 9 42 57 43
rect 26 29 30 42
rect 35 34 36 38
rect 40 34 50 38
rect 54 34 55 38
rect 16 27 20 28
rect 16 19 20 23
rect 26 22 30 25
rect 26 17 30 18
rect 36 27 40 28
rect 49 26 55 34
rect 36 19 40 23
rect 16 12 20 15
rect 36 12 40 15
rect -2 2 66 12
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
<< ntransistor >>
rect 22 14 24 30
rect 32 14 34 30
<< ptransistor >>
rect 9 42 11 70
rect 19 42 21 70
rect 29 42 31 70
rect 39 42 41 70
rect 49 42 51 58
<< polycontact >>
rect 36 34 40 38
rect 50 34 54 38
<< ndcontact >>
rect 16 23 20 27
rect 16 15 20 19
rect 26 25 30 29
rect 26 18 30 22
rect 36 23 40 27
rect 36 15 40 19
<< pdcontact >>
rect 3 65 7 69
rect 3 58 7 62
rect 13 50 17 54
rect 13 43 17 47
rect 23 65 27 69
rect 23 58 27 62
rect 33 50 37 54
rect 33 43 37 47
rect 43 53 47 57
rect 53 50 57 54
rect 53 43 57 47
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
<< psubstratepdiff >>
rect 0 2 64 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 64 2
rect 0 -3 64 -2
<< nsubstratendiff >>
rect 0 82 64 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 64 82
rect 0 77 64 78
<< labels >>
rlabel metal1 12 44 12 44 6 z
rlabel metal1 28 32 28 32 6 z
rlabel metal1 20 44 20 44 6 z
rlabel metal1 32 6 32 6 6 vss
rlabel metal1 44 36 44 36 6 a
rlabel metal1 44 44 44 44 6 z
rlabel metal1 36 48 36 48 6 z
rlabel metal1 32 74 32 74 6 vdd
rlabel metal1 52 32 52 32 6 a
rlabel metal1 52 44 52 44 6 z
rlabel metal1 60 52 60 52 6 z
<< end >>
