magic
tech scmos
timestamp 1179387652
<< checkpaint >>
rect -22 -22 158 94
<< ab >>
rect 0 0 136 72
<< pwell >>
rect -4 -4 140 32
<< nwell >>
rect -4 32 140 76
<< polysilicon >>
rect 20 66 22 70
rect 30 66 32 70
rect 45 66 47 70
rect 55 66 57 70
rect 85 66 87 70
rect 95 66 97 70
rect 105 66 107 70
rect 115 66 117 70
rect 125 66 127 70
rect 71 59 77 60
rect 65 51 67 56
rect 71 55 72 59
rect 76 55 77 59
rect 71 54 77 55
rect 75 51 77 54
rect 20 35 22 38
rect 30 35 32 38
rect 45 35 47 38
rect 55 35 57 38
rect 9 34 51 35
rect 9 30 10 34
rect 14 33 51 34
rect 14 30 21 33
rect 9 29 21 30
rect 9 26 11 29
rect 19 26 21 29
rect 39 26 41 33
rect 49 26 51 33
rect 55 34 61 35
rect 55 30 56 34
rect 60 30 61 34
rect 65 33 67 38
rect 75 33 77 38
rect 85 35 87 38
rect 95 35 97 38
rect 105 35 107 38
rect 85 34 97 35
rect 65 31 80 33
rect 55 29 61 30
rect 59 26 61 29
rect 66 26 68 31
rect 78 26 80 31
rect 85 30 86 34
rect 90 33 97 34
rect 101 34 107 35
rect 90 30 91 33
rect 85 29 91 30
rect 101 30 102 34
rect 106 30 107 34
rect 101 29 107 30
rect 115 35 117 38
rect 125 35 127 38
rect 115 34 127 35
rect 115 30 122 34
rect 126 30 127 34
rect 115 29 127 30
rect 85 26 87 29
rect 115 26 117 29
rect 125 26 127 29
rect 9 11 11 15
rect 19 4 21 9
rect 39 7 41 12
rect 49 7 51 12
rect 59 2 61 7
rect 66 2 68 7
rect 115 8 117 12
rect 125 8 127 12
rect 78 2 80 7
rect 85 2 87 7
<< ndiffusion >>
rect 2 20 9 26
rect 2 16 3 20
rect 7 16 9 20
rect 2 15 9 16
rect 11 25 19 26
rect 11 21 13 25
rect 17 21 19 25
rect 11 15 19 21
rect 14 9 19 15
rect 21 14 28 26
rect 21 10 23 14
rect 27 10 28 14
rect 32 25 39 26
rect 32 21 33 25
rect 37 21 39 25
rect 32 18 39 21
rect 32 14 33 18
rect 37 14 39 18
rect 32 12 39 14
rect 41 25 49 26
rect 41 21 43 25
rect 47 21 49 25
rect 41 12 49 21
rect 51 25 59 26
rect 51 21 53 25
rect 57 21 59 25
rect 51 18 59 21
rect 51 14 53 18
rect 57 14 59 18
rect 51 12 59 14
rect 21 9 28 10
rect 54 7 59 12
rect 61 7 66 26
rect 68 8 78 26
rect 68 7 71 8
rect 70 4 71 7
rect 75 7 78 8
rect 80 7 85 26
rect 87 19 92 26
rect 87 18 94 19
rect 87 14 89 18
rect 93 14 94 18
rect 87 13 94 14
rect 87 7 92 13
rect 108 17 115 26
rect 108 13 109 17
rect 113 13 115 17
rect 108 12 115 13
rect 117 25 125 26
rect 117 21 119 25
rect 123 21 125 25
rect 117 18 125 21
rect 117 14 119 18
rect 123 14 125 18
rect 117 12 125 14
rect 127 17 134 26
rect 127 13 129 17
rect 133 13 134 17
rect 127 12 134 13
rect 75 4 76 7
rect 70 3 76 4
<< pdiffusion >>
rect 13 65 20 66
rect 13 61 14 65
rect 18 61 20 65
rect 13 58 20 61
rect 13 54 14 58
rect 18 54 20 58
rect 13 38 20 54
rect 22 50 30 66
rect 22 46 24 50
rect 28 46 30 50
rect 22 43 30 46
rect 22 39 24 43
rect 28 39 30 43
rect 22 38 30 39
rect 32 65 45 66
rect 32 61 36 65
rect 40 61 45 65
rect 32 58 45 61
rect 32 54 36 58
rect 40 54 45 58
rect 32 38 45 54
rect 47 58 55 66
rect 47 54 49 58
rect 53 54 55 58
rect 47 51 55 54
rect 47 47 49 51
rect 53 47 55 51
rect 47 38 55 47
rect 57 51 62 66
rect 80 51 85 66
rect 57 50 65 51
rect 57 46 59 50
rect 63 46 65 50
rect 57 43 65 46
rect 57 39 59 43
rect 63 39 65 43
rect 57 38 65 39
rect 67 43 75 51
rect 67 39 69 43
rect 73 39 75 43
rect 67 38 75 39
rect 77 50 85 51
rect 77 46 79 50
rect 83 46 85 50
rect 77 38 85 46
rect 87 59 95 66
rect 87 55 89 59
rect 93 55 95 59
rect 87 43 95 55
rect 87 39 89 43
rect 93 39 95 43
rect 87 38 95 39
rect 97 58 105 66
rect 97 54 99 58
rect 103 54 105 58
rect 97 51 105 54
rect 97 47 99 51
rect 103 47 105 51
rect 97 38 105 47
rect 107 50 115 66
rect 107 46 109 50
rect 113 46 115 50
rect 107 43 115 46
rect 107 39 109 43
rect 113 39 115 43
rect 107 38 115 39
rect 117 65 125 66
rect 117 61 119 65
rect 123 61 125 65
rect 117 58 125 61
rect 117 54 119 58
rect 123 54 125 58
rect 117 38 125 54
rect 127 51 132 66
rect 127 50 134 51
rect 127 46 129 50
rect 133 46 134 50
rect 127 43 134 46
rect 127 39 129 43
rect 133 39 134 43
rect 127 38 134 39
<< metal1 >>
rect -2 68 138 72
rect -2 64 4 68
rect 8 65 69 68
rect 8 64 14 65
rect 18 64 36 65
rect 14 58 18 61
rect 35 61 36 64
rect 40 64 69 65
rect 73 65 138 68
rect 73 64 119 65
rect 40 61 41 64
rect 35 58 41 61
rect 123 64 138 65
rect 35 54 36 58
rect 40 54 41 58
rect 49 58 72 59
rect 53 55 72 58
rect 76 55 89 59
rect 93 55 94 59
rect 98 58 103 59
rect 14 53 18 54
rect 49 51 53 54
rect 23 46 24 50
rect 28 47 49 50
rect 98 54 99 58
rect 98 51 103 54
rect 119 58 123 61
rect 119 53 123 54
rect 98 50 99 51
rect 28 46 53 47
rect 58 46 59 50
rect 63 46 79 50
rect 83 47 99 50
rect 83 46 103 47
rect 108 50 113 51
rect 108 46 109 50
rect 23 43 28 46
rect 2 35 6 43
rect 23 39 24 43
rect 58 43 63 46
rect 108 43 113 46
rect 129 50 134 51
rect 133 46 134 50
rect 129 43 134 46
rect 58 42 59 43
rect 23 38 28 39
rect 34 39 59 42
rect 34 38 63 39
rect 68 39 69 43
rect 73 39 74 43
rect 2 34 14 35
rect 2 30 10 34
rect 2 29 14 30
rect 23 25 27 38
rect 34 25 38 38
rect 68 34 74 39
rect 88 39 89 43
rect 93 42 94 43
rect 93 39 103 42
rect 108 39 109 43
rect 113 39 129 43
rect 133 39 134 43
rect 88 38 103 39
rect 99 34 103 38
rect 12 21 13 25
rect 17 21 27 25
rect 32 21 33 25
rect 37 21 38 25
rect 42 30 56 34
rect 60 30 86 34
rect 90 30 93 34
rect 99 30 102 34
rect 106 30 107 34
rect 42 25 48 30
rect 89 26 93 30
rect 112 26 116 39
rect 121 34 134 35
rect 121 30 122 34
rect 126 30 134 34
rect 42 21 43 25
rect 47 21 48 25
rect 53 25 57 26
rect 89 25 123 26
rect 89 22 119 25
rect 3 20 7 21
rect 3 8 7 16
rect 32 18 38 21
rect 53 18 57 21
rect 130 21 134 30
rect 119 18 123 21
rect 23 14 27 15
rect 32 14 33 18
rect 37 14 53 18
rect 57 14 89 18
rect 93 14 95 18
rect 109 17 113 18
rect 23 8 27 10
rect 119 13 123 14
rect 128 13 129 17
rect 133 13 134 17
rect 109 8 113 13
rect 128 8 134 13
rect -2 4 4 8
rect 8 4 71 8
rect 75 4 99 8
rect 103 4 138 8
rect -2 0 138 4
<< ntransistor >>
rect 9 15 11 26
rect 19 9 21 26
rect 39 12 41 26
rect 49 12 51 26
rect 59 7 61 26
rect 66 7 68 26
rect 78 7 80 26
rect 85 7 87 26
rect 115 12 117 26
rect 125 12 127 26
<< ptransistor >>
rect 20 38 22 66
rect 30 38 32 66
rect 45 38 47 66
rect 55 38 57 66
rect 65 38 67 51
rect 75 38 77 51
rect 85 38 87 66
rect 95 38 97 66
rect 105 38 107 66
rect 115 38 117 66
rect 125 38 127 66
<< polycontact >>
rect 72 55 76 59
rect 10 30 14 34
rect 56 30 60 34
rect 86 30 90 34
rect 102 30 106 34
rect 122 30 126 34
<< ndcontact >>
rect 3 16 7 20
rect 13 21 17 25
rect 23 10 27 14
rect 33 21 37 25
rect 33 14 37 18
rect 43 21 47 25
rect 53 21 57 25
rect 53 14 57 18
rect 71 4 75 8
rect 89 14 93 18
rect 109 13 113 17
rect 119 21 123 25
rect 119 14 123 18
rect 129 13 133 17
<< pdcontact >>
rect 14 61 18 65
rect 14 54 18 58
rect 24 46 28 50
rect 24 39 28 43
rect 36 61 40 65
rect 36 54 40 58
rect 49 54 53 58
rect 49 47 53 51
rect 59 46 63 50
rect 59 39 63 43
rect 69 39 73 43
rect 79 46 83 50
rect 89 55 93 59
rect 89 39 93 43
rect 99 54 103 58
rect 99 47 103 51
rect 109 46 113 50
rect 109 39 113 43
rect 119 61 123 65
rect 119 54 123 58
rect 129 46 133 50
rect 129 39 133 43
<< psubstratepcontact >>
rect 4 4 8 8
rect 99 4 103 8
<< nsubstratencontact >>
rect 4 64 8 68
rect 69 64 73 68
<< psubstratepdiff >>
rect 3 8 9 9
rect 3 4 4 8
rect 8 4 9 8
rect 3 3 9 4
rect 98 8 104 24
rect 98 4 99 8
rect 103 4 104 8
rect 98 3 104 4
<< nsubstratendiff >>
rect 3 68 9 69
rect 3 64 4 68
rect 8 64 9 68
rect 68 68 74 69
rect 3 40 9 64
rect 68 64 69 68
rect 73 64 74 68
rect 68 63 74 64
<< labels >>
rlabel polycontact 88 32 88 32 6 an
rlabel polycontact 74 57 74 57 6 bn
rlabel polycontact 104 32 104 32 6 bn
rlabel polycontact 12 32 12 32 6 b
rlabel metal1 4 36 4 36 6 b
rlabel metal1 44 16 44 16 6 z
rlabel metal1 19 23 19 23 6 bn
rlabel ndcontact 36 24 36 24 6 z
rlabel metal1 45 27 45 27 6 an
rlabel metal1 44 40 44 40 6 z
rlabel metal1 25 35 25 35 6 bn
rlabel metal1 51 52 51 52 6 bn
rlabel metal1 68 4 68 4 6 vss
rlabel metal1 76 16 76 16 6 z
rlabel metal1 68 16 68 16 6 z
rlabel metal1 60 16 60 16 6 z
rlabel metal1 52 16 52 16 6 z
rlabel metal1 52 40 52 40 6 z
rlabel pdcontact 60 40 60 40 6 z
rlabel metal1 71 36 71 36 6 an
rlabel metal1 76 48 76 48 6 z
rlabel metal1 68 48 68 48 6 z
rlabel metal1 68 68 68 68 6 vdd
rlabel ndcontact 92 16 92 16 6 z
rlabel metal1 84 16 84 16 6 z
rlabel metal1 101 36 101 36 6 bn
rlabel metal1 67 32 67 32 6 an
rlabel pdcontact 91 40 91 40 6 bn
rlabel metal1 84 48 84 48 6 z
rlabel metal1 100 52 100 52 6 z
rlabel metal1 92 48 92 48 6 z
rlabel metal1 71 57 71 57 6 bn
rlabel metal1 121 19 121 19 6 an
rlabel metal1 132 28 132 28 6 a
rlabel polycontact 124 32 124 32 6 a
rlabel metal1 131 45 131 45 6 an
rlabel metal1 121 41 121 41 6 an
rlabel metal1 110 45 110 45 6 an
<< end >>
