magic
tech scmos
timestamp 1179386589
<< checkpaint >>
rect -22 -25 86 105
<< ab >>
rect 0 0 64 80
<< pwell >>
rect -4 -7 68 36
<< nwell >>
rect -4 36 68 87
<< polysilicon >>
rect 37 70 39 74
rect 49 70 51 74
rect 15 63 17 67
rect 25 63 27 67
rect 15 46 17 49
rect 25 46 27 49
rect 15 45 27 46
rect 15 44 18 45
rect 17 41 18 44
rect 22 44 27 45
rect 22 41 23 44
rect 17 40 23 41
rect 7 38 13 39
rect 7 34 8 38
rect 12 35 13 38
rect 12 34 14 35
rect 7 33 14 34
rect 12 30 14 33
rect 19 30 21 40
rect 37 39 39 42
rect 33 38 39 39
rect 33 35 34 38
rect 26 34 34 35
rect 38 34 39 38
rect 49 39 51 42
rect 49 38 55 39
rect 26 33 39 34
rect 26 30 28 33
rect 36 30 38 33
rect 43 30 45 35
rect 49 34 50 38
rect 54 34 55 38
rect 49 33 55 34
rect 50 30 52 33
rect 12 11 14 16
rect 19 8 21 16
rect 26 12 28 16
rect 36 12 38 16
rect 43 8 45 16
rect 50 11 52 16
rect 19 6 45 8
<< ndiffusion >>
rect 2 28 12 30
rect 2 24 3 28
rect 7 24 12 28
rect 2 21 12 24
rect 2 17 3 21
rect 7 17 12 21
rect 2 16 12 17
rect 14 16 19 30
rect 21 16 26 30
rect 28 29 36 30
rect 28 25 30 29
rect 34 25 36 29
rect 28 16 36 25
rect 38 16 43 30
rect 45 16 50 30
rect 52 28 60 30
rect 52 24 54 28
rect 58 24 60 28
rect 52 21 60 24
rect 52 17 54 21
rect 58 17 60 21
rect 52 16 60 17
<< pdiffusion >>
rect 29 69 37 70
rect 29 65 30 69
rect 34 65 37 69
rect 29 63 37 65
rect 6 62 15 63
rect 6 58 8 62
rect 12 58 15 62
rect 6 49 15 58
rect 17 62 25 63
rect 17 58 19 62
rect 23 58 25 62
rect 17 54 25 58
rect 17 50 19 54
rect 23 50 25 54
rect 17 49 25 50
rect 27 62 37 63
rect 27 58 30 62
rect 34 58 37 62
rect 27 49 37 58
rect 29 42 37 49
rect 39 62 49 70
rect 39 58 42 62
rect 46 58 49 62
rect 39 54 49 58
rect 39 50 42 54
rect 46 50 49 54
rect 39 42 49 50
rect 51 69 59 70
rect 51 65 53 69
rect 57 65 59 69
rect 51 62 59 65
rect 51 58 53 62
rect 57 58 59 62
rect 51 42 59 58
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect -2 69 66 78
rect -2 68 30 69
rect 7 62 13 68
rect 29 65 30 68
rect 34 68 53 69
rect 34 65 35 68
rect 7 58 8 62
rect 12 58 13 62
rect 18 62 23 63
rect 18 58 19 62
rect 29 62 35 65
rect 52 65 53 68
rect 57 68 66 69
rect 57 65 58 68
rect 52 62 58 65
rect 29 58 30 62
rect 34 58 35 62
rect 41 58 42 62
rect 46 58 47 62
rect 52 58 53 62
rect 57 58 58 62
rect 9 46 14 55
rect 18 54 23 58
rect 41 54 47 58
rect 18 50 19 54
rect 23 50 42 54
rect 46 50 47 54
rect 9 45 22 46
rect 9 42 18 45
rect 7 34 8 38
rect 12 34 14 38
rect 3 28 7 29
rect 3 21 7 24
rect 10 22 14 34
rect 18 33 22 41
rect 26 25 30 50
rect 34 42 47 46
rect 34 38 38 42
rect 34 33 38 34
rect 42 34 50 38
rect 54 34 55 38
rect 34 25 35 29
rect 42 22 46 34
rect 10 18 46 22
rect 54 28 58 29
rect 54 21 58 24
rect 3 12 7 17
rect 54 12 58 17
rect -2 2 66 12
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
<< ntransistor >>
rect 12 16 14 30
rect 19 16 21 30
rect 26 16 28 30
rect 36 16 38 30
rect 43 16 45 30
rect 50 16 52 30
<< ptransistor >>
rect 15 49 17 63
rect 25 49 27 63
rect 37 42 39 70
rect 49 42 51 70
<< polycontact >>
rect 18 41 22 45
rect 8 34 12 38
rect 34 34 38 38
rect 50 34 54 38
<< ndcontact >>
rect 3 24 7 28
rect 3 17 7 21
rect 30 25 34 29
rect 54 24 58 28
rect 54 17 58 21
<< pdcontact >>
rect 30 65 34 69
rect 8 58 12 62
rect 19 58 23 62
rect 19 50 23 54
rect 30 58 34 62
rect 42 58 46 62
rect 42 50 46 54
rect 53 65 57 69
rect 53 58 57 62
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
<< psubstratepdiff >>
rect 0 2 64 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 64 2
rect 0 -3 64 -2
<< nsubstratendiff >>
rect 0 82 64 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 64 82
rect 0 77 64 78
<< labels >>
rlabel metal1 12 28 12 28 6 a
rlabel metal1 20 20 20 20 6 a
rlabel metal1 20 36 20 36 6 b
rlabel metal1 12 48 12 48 6 b
rlabel pdcontact 20 60 20 60 6 z
rlabel metal1 32 6 32 6 6 vss
rlabel metal1 28 20 28 20 6 a
rlabel metal1 36 20 36 20 6 a
rlabel metal1 28 44 28 44 6 z
rlabel polycontact 36 36 36 36 6 c
rlabel metal1 36 52 36 52 6 z
rlabel metal1 32 74 32 74 6 vdd
rlabel metal1 44 28 44 28 6 a
rlabel metal1 44 44 44 44 6 c
rlabel metal1 44 56 44 56 6 z
rlabel polycontact 52 36 52 36 6 a
<< end >>
