magic
tech scmos
timestamp 1179386090
<< checkpaint >>
rect -22 -25 118 105
<< ab >>
rect 0 0 96 80
<< pwell >>
rect -4 -7 100 36
<< nwell >>
rect -4 36 100 87
<< polysilicon >>
rect 13 70 15 74
rect 20 70 22 74
rect 30 70 32 74
rect 37 70 39 74
rect 49 70 51 74
rect 56 70 58 74
rect 66 70 68 74
rect 73 70 75 74
rect 85 60 87 65
rect 13 42 15 45
rect 2 41 15 42
rect 2 37 3 41
rect 7 40 15 41
rect 20 42 22 45
rect 30 42 32 45
rect 20 41 33 42
rect 20 40 28 41
rect 7 37 13 40
rect 2 36 13 37
rect 27 37 28 40
rect 32 37 33 41
rect 27 36 33 37
rect 11 27 13 36
rect 17 35 23 36
rect 17 31 18 35
rect 22 32 23 35
rect 37 32 39 45
rect 49 42 51 45
rect 47 40 51 42
rect 56 42 58 45
rect 66 42 68 45
rect 56 41 69 42
rect 56 40 64 41
rect 47 36 49 40
rect 63 37 64 40
rect 68 37 69 41
rect 63 36 69 37
rect 73 39 75 45
rect 73 38 79 39
rect 22 31 30 32
rect 17 30 30 31
rect 18 27 20 30
rect 28 27 30 30
rect 35 30 39 32
rect 43 35 49 36
rect 43 31 44 35
rect 48 31 49 35
rect 43 30 49 31
rect 53 35 59 36
rect 53 31 54 35
rect 58 32 59 35
rect 73 34 74 38
rect 78 34 79 38
rect 85 36 87 42
rect 73 33 79 34
rect 83 33 87 36
rect 73 32 75 33
rect 58 31 66 32
rect 53 30 66 31
rect 35 27 37 30
rect 47 27 49 30
rect 54 27 56 30
rect 64 27 66 30
rect 71 30 75 32
rect 83 30 85 33
rect 71 27 73 30
rect 11 8 13 16
rect 18 12 20 16
rect 28 12 30 16
rect 35 8 37 16
rect 11 6 37 8
rect 47 11 49 16
rect 54 11 56 16
rect 64 8 66 16
rect 71 12 73 16
rect 83 8 85 21
rect 64 6 85 8
<< ndiffusion >>
rect 78 27 83 30
rect 2 21 11 27
rect 2 17 3 21
rect 7 17 11 21
rect 2 16 11 17
rect 13 16 18 27
rect 20 22 28 27
rect 20 18 22 22
rect 26 18 28 22
rect 20 16 28 18
rect 30 16 35 27
rect 37 16 47 27
rect 49 16 54 27
rect 56 21 64 27
rect 56 17 58 21
rect 62 17 64 21
rect 56 16 64 17
rect 66 16 71 27
rect 73 26 83 27
rect 73 22 77 26
rect 81 22 83 26
rect 73 21 83 22
rect 85 29 92 30
rect 85 25 87 29
rect 91 25 92 29
rect 85 24 92 25
rect 85 21 90 24
rect 73 16 81 21
rect 39 12 45 16
rect 39 8 40 12
rect 44 8 45 12
rect 39 7 45 8
<< pdiffusion >>
rect 5 69 13 70
rect 5 65 7 69
rect 11 65 13 69
rect 5 45 13 65
rect 15 45 20 70
rect 22 62 30 70
rect 22 58 24 62
rect 28 58 30 62
rect 22 45 30 58
rect 32 45 37 70
rect 39 69 49 70
rect 39 65 42 69
rect 46 65 49 69
rect 39 45 49 65
rect 51 45 56 70
rect 58 62 66 70
rect 58 58 60 62
rect 64 58 66 62
rect 58 45 66 58
rect 68 45 73 70
rect 75 62 83 70
rect 75 58 78 62
rect 82 60 83 62
rect 82 58 85 60
rect 75 55 85 58
rect 75 51 78 55
rect 82 51 85 55
rect 75 45 85 51
rect 77 42 85 45
rect 87 55 92 60
rect 87 54 94 55
rect 87 50 89 54
rect 93 50 94 54
rect 87 47 94 50
rect 87 43 89 47
rect 93 43 94 47
rect 87 42 94 43
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect -2 69 98 78
rect -2 68 7 69
rect 6 65 7 68
rect 11 68 42 69
rect 11 65 12 68
rect 41 65 42 68
rect 46 68 98 69
rect 46 65 47 68
rect 78 62 82 68
rect 2 58 15 62
rect 19 58 24 62
rect 28 58 60 62
rect 64 58 65 62
rect 2 42 6 58
rect 19 55 23 58
rect 11 51 23 55
rect 78 55 82 58
rect 11 47 15 51
rect 26 50 68 54
rect 78 50 82 51
rect 89 54 93 55
rect 26 48 30 50
rect 10 43 15 47
rect 20 44 30 48
rect 64 46 68 50
rect 89 47 93 50
rect 2 41 7 42
rect 2 37 3 41
rect 2 36 7 37
rect 2 33 6 36
rect 10 22 14 43
rect 20 35 24 44
rect 33 42 56 46
rect 33 41 39 42
rect 27 37 28 41
rect 32 37 39 41
rect 17 31 18 35
rect 22 31 24 35
rect 33 34 39 37
rect 44 35 48 36
rect 52 35 56 42
rect 64 43 89 46
rect 93 43 94 46
rect 64 42 94 43
rect 64 41 68 42
rect 64 36 68 37
rect 52 31 54 35
rect 58 31 59 35
rect 73 34 74 38
rect 78 34 79 38
rect 73 33 79 34
rect 44 30 48 31
rect 41 28 48 30
rect 65 29 79 33
rect 90 29 94 42
rect 65 28 71 29
rect 41 26 71 28
rect 44 24 69 26
rect 76 22 77 26
rect 81 22 82 26
rect 86 25 87 29
rect 91 25 94 29
rect 3 21 7 22
rect 10 18 22 22
rect 26 21 31 22
rect 26 18 58 21
rect 27 17 58 18
rect 62 17 64 21
rect 3 12 7 17
rect 76 12 82 22
rect -2 8 40 12
rect 44 8 98 12
rect -2 2 98 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
<< ntransistor >>
rect 11 16 13 27
rect 18 16 20 27
rect 28 16 30 27
rect 35 16 37 27
rect 47 16 49 27
rect 54 16 56 27
rect 64 16 66 27
rect 71 16 73 27
rect 83 21 85 30
<< ptransistor >>
rect 13 45 15 70
rect 20 45 22 70
rect 30 45 32 70
rect 37 45 39 70
rect 49 45 51 70
rect 56 45 58 70
rect 66 45 68 70
rect 73 45 75 70
rect 85 42 87 60
<< polycontact >>
rect 3 37 7 41
rect 28 37 32 41
rect 18 31 22 35
rect 64 37 68 41
rect 44 31 48 35
rect 54 31 58 35
rect 74 34 78 38
<< ndcontact >>
rect 3 17 7 21
rect 22 18 26 22
rect 58 17 62 21
rect 77 22 81 26
rect 87 25 91 29
rect 40 8 44 12
<< pdcontact >>
rect 7 65 11 69
rect 24 58 28 62
rect 42 65 46 69
rect 60 58 64 62
rect 78 58 82 62
rect 78 51 82 55
rect 89 50 93 54
rect 89 43 93 47
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
rect 90 -2 94 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
rect 90 78 94 82
<< psubstratepdiff >>
rect 0 2 96 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 96 2
rect 0 -3 96 -2
<< nsubstratendiff >>
rect 0 82 96 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 96 82
rect 0 77 96 78
<< labels >>
rlabel ntransistor 19 24 19 24 6 sn
rlabel ptransistor 67 55 67 55 6 sn
rlabel metal1 4 44 4 44 6 a0
rlabel metal1 12 36 12 36 6 z
rlabel metal1 12 60 12 60 6 a0
rlabel metal1 20 20 20 20 6 z
rlabel metal1 28 20 28 20 6 z
rlabel metal1 22 39 22 39 6 sn
rlabel metal1 28 60 28 60 6 z
rlabel metal1 48 6 48 6 6 vss
rlabel metal1 44 28 44 28 6 a1
rlabel metal1 36 40 36 40 6 s
rlabel metal1 52 44 52 44 6 s
rlabel metal1 44 44 44 44 6 s
rlabel metal1 36 60 36 60 6 z
rlabel metal1 52 60 52 60 6 z
rlabel metal1 44 60 44 60 6 z
rlabel metal1 48 74 48 74 6 vdd
rlabel metal1 68 28 68 28 6 a1
rlabel polycontact 76 36 76 36 6 a1
rlabel metal1 60 60 60 60 6 z
rlabel metal1 92 35 92 35 6 sn
rlabel metal1 79 44 79 44 6 sn
rlabel metal1 91 48 91 48 6 sn
<< end >>
