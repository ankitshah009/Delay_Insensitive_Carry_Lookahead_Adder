magic
tech scmos
timestamp 1170759849
<< checkpaint >>
rect -22 -26 118 114
<< ab >>
rect 0 0 96 88
<< pwell >>
rect -4 -8 100 40
<< nwell >>
rect -4 40 100 96
<< polysilicon >>
rect 2 82 11 83
rect 2 78 6 82
rect 10 78 11 82
rect 2 77 11 78
rect 9 74 11 77
rect 21 82 30 83
rect 21 78 25 82
rect 29 78 30 82
rect 21 77 30 78
rect 34 77 43 83
rect 21 74 23 77
rect 41 74 43 77
rect 53 77 62 83
rect 66 82 75 83
rect 66 78 67 82
rect 71 78 75 82
rect 66 77 75 78
rect 53 74 55 77
rect 73 74 75 77
rect 85 77 94 83
rect 85 74 87 77
rect 9 43 11 46
rect 21 43 23 46
rect 41 43 43 46
rect 53 43 55 46
rect 73 43 75 46
rect 85 43 87 46
rect 2 37 14 43
rect 18 42 30 43
rect 18 38 19 42
rect 23 38 30 42
rect 18 37 30 38
rect 34 42 46 43
rect 34 38 35 42
rect 39 38 46 42
rect 34 37 46 38
rect 50 42 62 43
rect 50 38 55 42
rect 59 38 62 42
rect 50 37 62 38
rect 66 37 78 43
rect 82 42 94 43
rect 82 38 86 42
rect 90 38 94 42
rect 82 37 94 38
rect 9 34 11 37
rect 21 34 23 37
rect 41 34 43 37
rect 53 34 55 37
rect 73 34 75 37
rect 85 34 87 37
rect 9 11 11 14
rect 2 5 11 11
rect 21 11 23 14
rect 41 11 43 14
rect 21 5 30 11
rect 34 5 43 11
rect 53 11 55 14
rect 73 11 75 14
rect 53 5 62 11
rect 66 5 75 11
rect 85 11 87 14
rect 85 5 94 11
<< ndiffusion >>
rect 2 14 9 34
rect 11 26 21 34
rect 11 22 14 26
rect 18 22 21 26
rect 11 19 21 22
rect 11 15 14 19
rect 18 15 21 19
rect 11 14 21 15
rect 23 33 30 34
rect 23 29 25 33
rect 29 29 30 33
rect 23 26 30 29
rect 23 22 25 26
rect 29 22 30 26
rect 23 14 30 22
rect 34 27 41 34
rect 34 23 35 27
rect 39 23 41 27
rect 34 19 41 23
rect 34 15 35 19
rect 39 15 41 19
rect 34 14 41 15
rect 43 14 53 34
rect 55 19 62 34
rect 55 15 57 19
rect 61 15 62 19
rect 55 14 62 15
rect 66 29 73 34
rect 66 25 67 29
rect 71 25 73 29
rect 66 22 73 25
rect 66 18 67 22
rect 71 18 73 22
rect 66 14 73 18
rect 75 33 85 34
rect 75 29 78 33
rect 82 29 85 33
rect 75 26 85 29
rect 75 22 78 26
rect 82 22 85 26
rect 75 14 85 22
rect 87 26 94 34
rect 87 22 89 26
rect 93 22 94 26
rect 87 19 94 22
rect 87 15 89 19
rect 93 15 94 19
rect 87 14 94 15
rect 13 2 19 14
rect 45 2 51 14
rect 77 2 83 14
<< pdiffusion >>
rect 13 74 19 86
rect 45 74 51 86
rect 77 77 83 86
rect 77 74 78 77
rect 2 46 9 74
rect 11 73 21 74
rect 11 69 14 73
rect 18 69 21 73
rect 11 66 21 69
rect 11 62 14 66
rect 18 62 21 66
rect 11 46 21 62
rect 23 62 30 74
rect 23 58 25 62
rect 29 58 30 62
rect 23 55 30 58
rect 23 51 25 55
rect 29 51 30 55
rect 23 46 30 51
rect 34 62 41 74
rect 34 58 35 62
rect 39 58 41 62
rect 34 46 41 58
rect 43 51 53 74
rect 43 47 46 51
rect 50 47 53 51
rect 43 46 53 47
rect 55 70 62 74
rect 55 66 57 70
rect 61 66 62 70
rect 55 46 62 66
rect 66 69 73 74
rect 66 65 67 69
rect 71 65 73 69
rect 66 62 73 65
rect 66 58 67 62
rect 71 58 73 62
rect 66 46 73 58
rect 75 73 78 74
rect 82 74 83 77
rect 82 73 85 74
rect 75 70 85 73
rect 75 66 78 70
rect 82 66 85 70
rect 75 46 85 66
rect 87 70 94 74
rect 87 66 89 70
rect 93 66 94 70
rect 87 63 94 66
rect 87 59 89 63
rect 93 59 94 63
rect 87 46 94 59
<< metal1 >>
rect -2 86 2 90
rect 10 86 22 90
rect 30 86 34 90
rect 42 86 54 90
rect 62 86 66 90
rect 74 86 86 90
rect 94 86 98 90
rect 6 82 10 86
rect 6 77 10 78
rect 14 82 18 86
rect 78 82 82 86
rect 24 78 25 82
rect 29 78 67 82
rect 71 78 72 82
rect 14 73 18 78
rect 78 77 82 78
rect 78 70 82 73
rect 14 66 18 69
rect 14 61 18 62
rect 25 66 57 70
rect 61 69 71 70
rect 61 66 67 69
rect 25 62 29 66
rect 78 65 82 66
rect 89 70 93 71
rect 67 62 71 65
rect 89 63 93 66
rect 34 58 35 62
rect 39 58 58 62
rect 25 55 29 58
rect 14 42 18 55
rect 29 51 39 54
rect 25 50 39 51
rect 35 42 39 50
rect 14 38 19 42
rect 23 38 24 42
rect 14 33 18 38
rect 35 35 39 38
rect 25 33 39 35
rect 29 31 39 33
rect 46 51 50 55
rect 14 26 18 27
rect 14 19 18 22
rect 25 26 29 29
rect 46 30 50 47
rect 54 42 58 58
rect 67 57 71 58
rect 78 59 89 62
rect 78 58 93 59
rect 78 42 82 58
rect 54 38 55 42
rect 59 38 82 42
rect 78 33 82 38
rect 86 42 90 55
rect 86 33 90 38
rect 46 29 71 30
rect 46 27 67 29
rect 34 23 35 27
rect 39 26 67 27
rect 39 23 50 26
rect 25 21 29 22
rect 38 19 42 23
rect 67 22 71 25
rect 34 15 35 19
rect 39 15 42 19
rect 57 19 61 20
rect 78 26 82 29
rect 78 21 82 22
rect 89 26 93 27
rect 67 17 71 18
rect 89 19 93 22
rect 14 10 18 15
rect 14 2 18 6
rect 57 10 61 15
rect 57 2 61 6
rect 89 10 93 15
rect 89 2 93 6
rect -2 -2 2 2
rect 10 -2 22 2
rect 30 -2 34 2
rect 42 -2 54 2
rect 62 -2 66 2
rect 74 -2 86 2
rect 94 -2 98 2
<< metal2 >>
rect -2 86 6 90
rect 10 86 22 90
rect 26 86 38 90
rect 42 86 54 90
rect 58 86 70 90
rect 74 86 86 90
rect 90 86 98 90
rect -2 82 98 86
rect -2 78 14 82
rect 18 78 78 82
rect 82 78 98 82
rect -2 76 98 78
rect -2 10 98 12
rect -2 6 14 10
rect 18 6 57 10
rect 61 6 89 10
rect 93 6 98 10
rect -2 2 98 6
rect -2 -2 6 2
rect 10 -2 22 2
rect 26 -2 38 2
rect 42 -2 54 2
rect 58 -2 70 2
rect 74 -2 86 2
rect 90 -2 98 2
<< ntransistor >>
rect 9 14 11 34
rect 21 14 23 34
rect 41 14 43 34
rect 53 14 55 34
rect 73 14 75 34
rect 85 14 87 34
<< ptransistor >>
rect 9 46 11 74
rect 21 46 23 74
rect 41 46 43 74
rect 53 46 55 74
rect 73 46 75 74
rect 85 46 87 74
<< polycontact >>
rect 6 78 10 82
rect 25 78 29 82
rect 67 78 71 82
rect 19 38 23 42
rect 35 38 39 42
rect 55 38 59 42
rect 86 38 90 42
<< ndcontact >>
rect 14 22 18 26
rect 14 15 18 19
rect 25 29 29 33
rect 25 22 29 26
rect 35 23 39 27
rect 35 15 39 19
rect 57 15 61 19
rect 67 25 71 29
rect 67 18 71 22
rect 78 29 82 33
rect 78 22 82 26
rect 89 22 93 26
rect 89 15 93 19
<< pdcontact >>
rect 14 69 18 73
rect 14 62 18 66
rect 25 58 29 62
rect 25 51 29 55
rect 35 58 39 62
rect 46 47 50 51
rect 57 66 61 70
rect 67 65 71 69
rect 67 58 71 62
rect 78 73 82 77
rect 78 66 82 70
rect 89 66 93 70
rect 89 59 93 63
<< m2contact >>
rect 6 86 10 90
rect 22 86 26 90
rect 38 86 42 90
rect 54 86 58 90
rect 70 86 74 90
rect 86 86 90 90
rect 14 78 18 82
rect 78 78 82 82
rect 14 6 18 10
rect 57 6 61 10
rect 89 6 93 10
rect 6 -2 10 2
rect 22 -2 26 2
rect 38 -2 42 2
rect 54 -2 58 2
rect 70 -2 74 2
rect 86 -2 90 2
<< psubstratepcontact >>
rect 2 -2 6 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 90 -2 94 2
<< nsubstratencontact >>
rect 2 86 6 90
rect 26 86 30 90
rect 34 86 38 90
rect 58 86 62 90
rect 66 86 70 90
rect 90 86 94 90
<< psubstratepdiff >>
rect 0 2 7 3
rect 25 2 39 3
rect 57 2 71 3
rect 89 2 96 3
rect 0 -2 2 2
rect 6 -2 7 2
rect 0 -3 7 -2
rect 25 -2 26 2
rect 30 -2 34 2
rect 38 -2 39 2
rect 25 -3 39 -2
rect 57 -2 58 2
rect 62 -2 66 2
rect 70 -2 71 2
rect 57 -3 71 -2
rect 89 -2 90 2
rect 94 -2 96 2
rect 89 -3 96 -2
<< nsubstratendiff >>
rect 0 90 7 91
rect 0 86 2 90
rect 6 86 7 90
rect 25 90 39 91
rect 25 86 26 90
rect 30 86 34 90
rect 38 86 39 90
rect 57 90 71 91
rect 57 86 58 90
rect 62 86 66 90
rect 70 86 71 90
rect 89 90 96 91
rect 89 86 90 90
rect 94 86 96 90
rect 0 85 7 86
rect 25 85 39 86
rect 57 85 71 86
rect 89 85 96 86
<< labels >>
rlabel metal1 16 44 16 44 6 b
rlabel metal1 40 20 40 20 6 z
rlabel metal1 56 28 56 28 6 z
rlabel metal1 48 40 48 40 6 z
rlabel metal1 64 28 64 28 6 z
rlabel metal1 88 44 88 44 6 a
rlabel metal2 48 6 48 6 6 vss
rlabel metal2 48 82 48 82 6 vdd
<< end >>
