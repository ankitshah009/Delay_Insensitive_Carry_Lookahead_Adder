magic
tech scmos
timestamp 1179386363
<< checkpaint >>
rect -22 -22 70 94
<< ab >>
rect 0 0 48 72
<< pwell >>
rect -4 -4 52 32
<< nwell >>
rect -4 32 52 76
<< polysilicon >>
rect 9 62 11 67
rect 19 62 21 67
rect 9 35 11 38
rect 19 35 21 38
rect 9 34 15 35
rect 9 30 10 34
rect 14 30 15 34
rect 9 29 15 30
rect 19 34 32 35
rect 19 30 26 34
rect 30 30 32 34
rect 40 34 46 35
rect 40 31 41 34
rect 19 29 32 30
rect 13 26 15 29
rect 20 26 22 29
rect 30 26 32 29
rect 37 30 41 31
rect 45 30 46 34
rect 37 29 46 30
rect 37 26 39 29
rect 13 2 15 6
rect 20 2 22 6
rect 30 2 32 6
rect 37 2 39 6
<< ndiffusion >>
rect 5 11 13 26
rect 5 7 7 11
rect 11 7 13 11
rect 5 6 13 7
rect 15 6 20 26
rect 22 18 30 26
rect 22 14 24 18
rect 28 14 30 18
rect 22 6 30 14
rect 32 6 37 26
rect 39 18 46 26
rect 39 14 41 18
rect 45 14 46 18
rect 39 11 46 14
rect 39 7 41 11
rect 45 7 46 11
rect 39 6 46 7
<< pdiffusion >>
rect 2 61 9 62
rect 2 57 3 61
rect 7 57 9 61
rect 2 53 9 57
rect 2 49 3 53
rect 7 49 9 53
rect 2 38 9 49
rect 11 50 19 62
rect 11 46 13 50
rect 17 46 19 50
rect 11 43 19 46
rect 11 39 13 43
rect 17 39 19 43
rect 11 38 19 39
rect 21 61 29 62
rect 21 57 23 61
rect 27 57 29 61
rect 21 53 29 57
rect 21 49 23 53
rect 27 49 29 53
rect 21 38 29 49
<< metal1 >>
rect -2 68 50 72
rect -2 64 40 68
rect 44 64 50 68
rect 3 61 7 64
rect 3 53 7 57
rect 23 61 27 64
rect 23 53 27 57
rect 3 48 7 49
rect 12 46 13 50
rect 17 46 18 50
rect 23 48 27 49
rect 12 43 18 46
rect 2 39 13 43
rect 17 39 18 43
rect 2 18 6 39
rect 25 38 39 42
rect 10 34 19 35
rect 14 30 19 34
rect 25 34 31 38
rect 25 30 26 34
rect 30 30 31 34
rect 40 30 41 34
rect 45 30 46 34
rect 10 29 19 30
rect 15 26 19 29
rect 40 26 46 30
rect 15 22 46 26
rect 2 14 24 18
rect 28 14 31 18
rect 40 14 41 18
rect 45 14 46 18
rect 40 11 46 14
rect 6 8 7 11
rect -2 7 7 8
rect 11 8 12 11
rect 40 8 41 11
rect 11 7 41 8
rect 45 8 46 11
rect 45 7 50 8
rect -2 0 50 7
<< ntransistor >>
rect 13 6 15 26
rect 20 6 22 26
rect 30 6 32 26
rect 37 6 39 26
<< ptransistor >>
rect 9 38 11 62
rect 19 38 21 62
<< polycontact >>
rect 10 30 14 34
rect 26 30 30 34
rect 41 30 45 34
<< ndcontact >>
rect 7 7 11 11
rect 24 14 28 18
rect 41 14 45 18
rect 41 7 45 11
<< pdcontact >>
rect 3 57 7 61
rect 3 49 7 53
rect 13 46 17 50
rect 13 39 17 43
rect 23 57 27 61
rect 23 49 27 53
<< nsubstratencontact >>
rect 40 64 44 68
<< nsubstratendiff >>
rect 39 68 45 69
rect 39 64 40 68
rect 44 64 45 68
rect 39 40 45 64
<< labels >>
rlabel metal1 4 32 4 32 6 z
rlabel metal1 20 16 20 16 6 z
rlabel metal1 12 16 12 16 6 z
rlabel polycontact 12 32 12 32 6 a
rlabel metal1 20 24 20 24 6 a
rlabel metal1 24 4 24 4 6 vss
rlabel metal1 28 16 28 16 6 z
rlabel metal1 28 24 28 24 6 a
rlabel metal1 28 36 28 36 6 b
rlabel metal1 24 68 24 68 6 vdd
rlabel metal1 36 24 36 24 6 a
rlabel metal1 36 40 36 40 6 b
<< end >>
