magic
tech scmos
timestamp 1179387166
<< checkpaint >>
rect -22 -25 62 105
<< ab >>
rect 0 0 40 80
<< pwell >>
rect -4 -7 44 36
<< nwell >>
rect -4 36 44 87
<< polysilicon >>
rect 9 70 11 74
rect 22 70 24 74
rect 29 70 31 74
rect 9 39 11 42
rect 22 39 24 42
rect 29 39 31 42
rect 9 38 15 39
rect 9 34 10 38
rect 14 34 15 38
rect 9 33 15 34
rect 19 38 25 39
rect 19 34 20 38
rect 24 34 25 38
rect 19 33 25 34
rect 29 38 38 39
rect 29 34 33 38
rect 37 34 38 38
rect 29 33 38 34
rect 9 30 11 33
rect 19 25 21 33
rect 29 27 31 33
rect 9 11 11 16
rect 19 12 21 17
rect 29 15 31 19
<< ndiffusion >>
rect 2 29 9 30
rect 2 25 3 29
rect 7 25 9 29
rect 2 22 9 25
rect 2 18 3 22
rect 7 18 9 22
rect 2 16 9 18
rect 11 25 16 30
rect 24 25 29 27
rect 11 22 19 25
rect 11 18 13 22
rect 17 18 19 22
rect 11 17 19 18
rect 21 24 29 25
rect 21 20 23 24
rect 27 20 29 24
rect 21 19 29 20
rect 31 24 38 27
rect 31 20 33 24
rect 37 20 38 24
rect 31 19 38 20
rect 21 17 26 19
rect 11 16 16 17
<< pdiffusion >>
rect 13 72 20 73
rect 13 70 14 72
rect 4 64 9 70
rect 2 63 9 64
rect 2 59 3 63
rect 7 59 9 63
rect 2 56 9 59
rect 2 52 3 56
rect 7 52 9 56
rect 2 51 9 52
rect 4 42 9 51
rect 11 68 14 70
rect 18 70 20 72
rect 18 68 22 70
rect 11 42 22 68
rect 24 42 29 70
rect 31 64 36 70
rect 31 63 38 64
rect 31 59 33 63
rect 37 59 38 63
rect 31 58 38 59
rect 31 42 36 58
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect -2 72 42 78
rect -2 68 14 72
rect 18 68 42 72
rect 2 59 3 63
rect 7 59 14 63
rect 2 57 14 59
rect 18 59 33 63
rect 37 59 38 63
rect 2 56 7 57
rect 2 52 3 56
rect 18 54 22 59
rect 2 51 7 52
rect 2 30 6 51
rect 10 50 22 54
rect 10 38 14 50
rect 26 49 38 55
rect 2 29 7 30
rect 2 25 3 29
rect 10 29 14 34
rect 18 39 22 47
rect 18 38 30 39
rect 18 34 20 38
rect 24 34 30 38
rect 18 33 30 34
rect 33 38 38 49
rect 37 34 38 38
rect 33 33 38 34
rect 10 25 27 29
rect 2 22 7 25
rect 23 24 27 25
rect 2 18 3 22
rect 2 17 7 18
rect 12 18 13 22
rect 17 18 18 22
rect 23 19 27 20
rect 32 20 33 24
rect 37 20 38 24
rect 12 12 18 18
rect 32 12 38 20
rect -2 2 42 12
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
<< ntransistor >>
rect 9 16 11 30
rect 19 17 21 25
rect 29 19 31 27
<< ptransistor >>
rect 9 42 11 70
rect 22 42 24 70
rect 29 42 31 70
<< polycontact >>
rect 10 34 14 38
rect 20 34 24 38
rect 33 34 37 38
<< ndcontact >>
rect 3 25 7 29
rect 3 18 7 22
rect 13 18 17 22
rect 23 20 27 24
rect 33 20 37 24
<< pdcontact >>
rect 3 59 7 63
rect 3 52 7 56
rect 14 68 18 72
rect 33 59 37 63
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
<< psubstratepdiff >>
rect 0 2 40 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 40 2
rect 0 -3 40 -2
<< nsubstratendiff >>
rect 0 82 40 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 40 82
rect 0 77 40 78
<< labels >>
rlabel polycontact 12 36 12 36 6 zn
rlabel metal1 4 40 4 40 6 z
rlabel metal1 12 39 12 39 6 zn
rlabel metal1 12 60 12 60 6 z
rlabel metal1 20 6 20 6 6 vss
rlabel metal1 25 24 25 24 6 zn
rlabel metal1 28 36 28 36 6 a
rlabel metal1 20 40 20 40 6 a
rlabel metal1 28 52 28 52 6 b
rlabel metal1 20 74 20 74 6 vdd
rlabel metal1 36 44 36 44 6 b
rlabel metal1 28 61 28 61 6 zn
<< end >>
