magic
tech scmos
timestamp 1179387355
<< checkpaint >>
rect -22 -22 46 94
<< ab >>
rect 0 0 24 72
<< pwell >>
rect -4 -4 28 32
<< nwell >>
rect -4 32 28 76
<< metal1 >>
rect -2 68 26 72
rect -2 64 10 68
rect 14 64 26 68
rect -2 4 10 8
rect 14 4 26 8
rect -2 0 26 4
<< psubstratepcontact >>
rect 10 4 14 8
<< nsubstratencontact >>
rect 10 64 14 68
<< psubstratepdiff >>
rect 6 8 18 26
rect 6 4 10 8
rect 14 4 18 8
rect 6 3 18 4
<< nsubstratendiff >>
rect 6 68 18 69
rect 6 64 10 68
rect 14 64 18 68
rect 6 38 18 64
<< labels >>
rlabel metal1 12 4 12 4 6 vss
rlabel metal1 12 68 12 68 6 vdd
<< end >>
