magic
tech scmos
timestamp 1179387679
<< checkpaint >>
rect -22 -22 94 94
<< ab >>
rect 0 0 72 72
<< pwell >>
rect -4 -4 76 32
<< nwell >>
rect -4 32 76 76
<< polysilicon >>
rect 38 63 63 65
rect 28 59 34 60
rect 28 55 29 59
rect 33 55 34 59
rect 18 50 20 55
rect 28 54 34 55
rect 28 50 30 54
rect 38 50 40 63
rect 61 59 63 63
rect 48 50 50 55
rect 18 35 20 38
rect 9 34 20 35
rect 9 30 10 34
rect 14 33 20 34
rect 14 30 15 33
rect 9 29 15 30
rect 28 30 30 38
rect 38 34 40 38
rect 48 34 50 38
rect 61 35 63 47
rect 57 34 63 35
rect 47 33 53 34
rect 47 30 48 33
rect 12 25 14 29
rect 22 25 24 29
rect 28 28 34 30
rect 32 25 34 28
rect 42 29 48 30
rect 52 29 53 33
rect 57 30 58 34
rect 62 30 63 34
rect 57 29 63 30
rect 42 28 53 29
rect 42 25 44 28
rect 61 25 63 29
rect 12 14 14 19
rect 22 11 24 19
rect 32 15 34 19
rect 42 15 44 19
rect 61 11 63 19
rect 22 9 63 11
<< ndiffusion >>
rect 4 19 12 25
rect 14 24 22 25
rect 14 20 16 24
rect 20 20 22 24
rect 14 19 22 20
rect 24 24 32 25
rect 24 20 26 24
rect 30 20 32 24
rect 24 19 32 20
rect 34 24 42 25
rect 34 20 36 24
rect 40 20 42 24
rect 34 19 42 20
rect 44 24 61 25
rect 44 20 55 24
rect 59 20 61 24
rect 44 19 61 20
rect 63 24 70 25
rect 63 20 65 24
rect 69 20 70 24
rect 63 19 70 20
rect 4 17 10 19
rect 4 13 5 17
rect 9 13 10 17
rect 4 12 10 13
<< pdiffusion >>
rect 52 60 59 61
rect 52 56 54 60
rect 58 59 59 60
rect 58 56 61 59
rect 52 50 61 56
rect 8 49 18 50
rect 8 45 10 49
rect 14 45 18 49
rect 8 38 18 45
rect 20 43 28 50
rect 20 39 22 43
rect 26 39 28 43
rect 20 38 28 39
rect 30 43 38 50
rect 30 39 32 43
rect 36 39 38 43
rect 30 38 38 39
rect 40 43 48 50
rect 40 39 42 43
rect 46 39 48 43
rect 40 38 48 39
rect 50 47 61 50
rect 63 53 68 59
rect 63 52 70 53
rect 63 48 65 52
rect 69 48 70 52
rect 63 47 70 48
rect 50 38 59 47
<< metal1 >>
rect -2 68 74 72
rect -2 64 4 68
rect 8 64 12 68
rect 16 64 74 68
rect 10 49 14 64
rect 53 60 59 64
rect 28 55 29 59
rect 33 55 49 59
rect 53 56 54 60
rect 58 56 59 60
rect 45 52 49 55
rect 10 44 14 45
rect 34 44 38 51
rect 45 48 65 52
rect 69 48 70 52
rect 32 43 38 44
rect 17 39 22 43
rect 26 39 27 43
rect 36 39 38 43
rect 2 34 14 35
rect 2 30 10 34
rect 2 29 14 30
rect 2 21 6 29
rect 17 25 21 39
rect 32 37 38 39
rect 41 43 46 44
rect 41 39 42 43
rect 41 38 46 39
rect 32 34 36 37
rect 16 24 21 25
rect 20 20 21 24
rect 25 30 36 34
rect 25 24 31 30
rect 41 24 45 38
rect 50 37 62 43
rect 58 34 62 37
rect 25 20 26 24
rect 30 20 31 24
rect 35 20 36 24
rect 40 20 45 24
rect 48 33 52 34
rect 58 29 62 30
rect 16 19 21 20
rect 17 17 21 19
rect 48 17 52 29
rect 66 25 70 48
rect 4 13 5 17
rect 9 13 10 17
rect 17 13 52 17
rect 55 24 59 25
rect 4 8 10 13
rect 55 8 59 20
rect 65 24 70 25
rect 69 20 70 24
rect 65 19 70 20
rect -2 4 15 8
rect 19 4 74 8
rect -2 0 74 4
<< ntransistor >>
rect 12 19 14 25
rect 22 19 24 25
rect 32 19 34 25
rect 42 19 44 25
rect 61 19 63 25
<< ptransistor >>
rect 18 38 20 50
rect 28 38 30 50
rect 38 38 40 50
rect 48 38 50 50
rect 61 47 63 59
<< polycontact >>
rect 29 55 33 59
rect 10 30 14 34
rect 48 29 52 33
rect 58 30 62 34
<< ndcontact >>
rect 16 20 20 24
rect 26 20 30 24
rect 36 20 40 24
rect 55 20 59 24
rect 65 20 69 24
rect 5 13 9 17
<< pdcontact >>
rect 54 56 58 60
rect 10 45 14 49
rect 22 39 26 43
rect 32 39 36 43
rect 42 39 46 43
rect 65 48 69 52
<< psubstratepcontact >>
rect 15 4 19 8
<< nsubstratencontact >>
rect 4 64 8 68
rect 12 64 16 68
<< psubstratepdiff >>
rect 14 8 20 9
rect 14 4 15 8
rect 19 4 20 8
rect 14 3 20 4
<< nsubstratendiff >>
rect 3 68 17 69
rect 3 64 4 68
rect 8 64 12 68
rect 16 64 17 68
rect 3 63 17 64
<< labels >>
rlabel polycontact 31 57 31 57 6 bn
rlabel ptransistor 49 41 49 41 6 an
rlabel metal1 4 28 4 28 6 a
rlabel polycontact 12 32 12 32 6 a
rlabel metal1 28 28 28 28 6 z
rlabel metal1 19 28 19 28 6 an
rlabel metal1 22 41 22 41 6 an
rlabel metal1 36 4 36 4 6 vss
rlabel metal1 50 23 50 23 6 an
rlabel metal1 40 22 40 22 6 ai
rlabel metal1 52 40 52 40 6 b
rlabel metal1 43 32 43 32 6 ai
rlabel metal1 36 44 36 44 6 z
rlabel metal1 38 57 38 57 6 bn
rlabel metal1 36 68 36 68 6 vdd
rlabel metal1 60 36 60 36 6 b
rlabel metal1 68 35 68 35 6 bn
rlabel metal1 57 50 57 50 6 bn
<< end >>
