magic
tech scmos
timestamp 1179385672
<< checkpaint >>
rect -22 -25 150 105
<< ab >>
rect 0 0 128 80
<< pwell >>
rect -4 -7 132 36
<< nwell >>
rect -4 36 132 87
<< polysilicon >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 39 70 41 74
rect 51 70 53 74
rect 58 70 60 74
rect 68 70 70 74
rect 75 70 77 74
rect 87 70 89 74
rect 97 70 99 74
rect 107 70 109 74
rect 117 58 119 63
rect 9 39 11 42
rect 2 38 11 39
rect 2 34 3 38
rect 7 34 11 38
rect 2 33 11 34
rect 9 30 11 33
rect 19 39 21 42
rect 29 39 31 42
rect 19 38 31 39
rect 19 34 26 38
rect 30 34 31 38
rect 19 33 31 34
rect 19 30 21 33
rect 29 30 31 33
rect 39 39 41 42
rect 51 39 53 42
rect 39 38 53 39
rect 39 34 42 38
rect 46 34 53 38
rect 39 33 53 34
rect 39 30 41 33
rect 51 30 53 33
rect 58 39 60 42
rect 68 39 70 42
rect 58 38 70 39
rect 58 34 65 38
rect 69 34 70 38
rect 58 33 70 34
rect 58 30 60 33
rect 68 30 70 33
rect 75 39 77 42
rect 75 38 83 39
rect 75 34 78 38
rect 82 34 83 38
rect 75 33 83 34
rect 87 35 89 42
rect 97 35 99 42
rect 87 34 99 35
rect 75 30 77 33
rect 87 30 91 34
rect 95 30 99 34
rect 9 11 11 16
rect 19 11 21 16
rect 29 11 31 16
rect 39 11 41 16
rect 87 29 99 30
rect 87 26 89 29
rect 97 26 99 29
rect 107 39 109 42
rect 117 39 119 42
rect 107 38 119 39
rect 107 34 114 38
rect 118 34 119 38
rect 107 33 119 34
rect 107 26 109 33
rect 117 26 119 33
rect 68 15 70 19
rect 75 15 77 19
rect 51 8 53 13
rect 58 8 60 13
rect 87 7 89 12
rect 97 7 99 12
rect 107 10 109 15
rect 117 10 119 15
<< ndiffusion >>
rect 2 28 9 30
rect 2 24 3 28
rect 7 24 9 28
rect 2 21 9 24
rect 2 17 3 21
rect 7 17 9 21
rect 2 16 9 17
rect 11 21 19 30
rect 11 17 13 21
rect 17 17 19 21
rect 11 16 19 17
rect 21 29 29 30
rect 21 25 23 29
rect 27 25 29 29
rect 21 16 29 25
rect 31 21 39 30
rect 31 17 33 21
rect 37 17 39 21
rect 31 16 39 17
rect 41 16 51 30
rect 43 13 51 16
rect 53 13 58 30
rect 60 29 68 30
rect 60 25 62 29
rect 66 25 68 29
rect 60 19 68 25
rect 70 19 75 30
rect 77 26 85 30
rect 77 19 87 26
rect 60 13 65 19
rect 43 12 49 13
rect 43 8 44 12
rect 48 8 49 12
rect 79 12 87 19
rect 89 21 97 26
rect 89 17 91 21
rect 95 17 97 21
rect 89 12 97 17
rect 99 20 107 26
rect 99 16 101 20
rect 105 16 107 20
rect 99 15 107 16
rect 109 25 117 26
rect 109 21 111 25
rect 115 21 117 25
rect 109 15 117 21
rect 119 20 126 26
rect 119 16 121 20
rect 125 16 126 20
rect 119 15 126 16
rect 99 12 105 15
rect 79 8 80 12
rect 84 8 85 12
rect 43 7 49 8
rect 79 7 85 8
<< pdiffusion >>
rect 2 69 9 70
rect 2 65 3 69
rect 7 65 9 69
rect 2 62 9 65
rect 2 58 3 62
rect 7 58 9 62
rect 2 42 9 58
rect 11 62 19 70
rect 11 58 13 62
rect 17 58 19 62
rect 11 42 19 58
rect 21 47 29 70
rect 21 43 23 47
rect 27 43 29 47
rect 21 42 29 43
rect 31 62 39 70
rect 31 58 33 62
rect 37 58 39 62
rect 31 42 39 58
rect 41 69 51 70
rect 41 65 44 69
rect 48 65 51 69
rect 41 42 51 65
rect 53 42 58 70
rect 60 47 68 70
rect 60 43 62 47
rect 66 43 68 47
rect 60 42 68 43
rect 70 42 75 70
rect 77 69 87 70
rect 77 65 80 69
rect 84 65 87 69
rect 77 42 87 65
rect 89 61 97 70
rect 89 57 91 61
rect 95 57 97 61
rect 89 54 97 57
rect 89 50 91 54
rect 95 50 97 54
rect 89 42 97 50
rect 99 69 107 70
rect 99 65 101 69
rect 105 65 107 69
rect 99 61 107 65
rect 99 57 101 61
rect 105 57 107 61
rect 99 42 107 57
rect 109 58 114 70
rect 109 54 117 58
rect 109 50 111 54
rect 115 50 117 54
rect 109 47 117 50
rect 109 43 111 47
rect 115 43 117 47
rect 109 42 117 43
rect 119 57 126 58
rect 119 53 121 57
rect 125 53 126 57
rect 119 49 126 53
rect 119 45 121 49
rect 125 45 126 49
rect 119 42 126 45
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect 118 78 122 82
rect 126 78 130 82
rect -2 69 130 78
rect -2 68 3 69
rect 7 68 44 69
rect 43 65 44 68
rect 48 68 80 69
rect 48 65 49 68
rect 79 65 80 68
rect 84 68 101 69
rect 84 65 85 68
rect 105 68 130 69
rect 3 62 7 65
rect 12 58 13 62
rect 17 58 33 62
rect 37 61 95 62
rect 37 58 91 61
rect 3 57 7 58
rect 91 54 95 57
rect 101 61 105 65
rect 101 56 105 57
rect 121 57 125 68
rect 2 50 79 54
rect 2 38 7 50
rect 22 46 23 47
rect 2 34 3 38
rect 2 33 7 34
rect 17 43 23 46
rect 27 43 28 47
rect 17 42 28 43
rect 17 30 21 42
rect 33 38 39 46
rect 25 34 26 38
rect 30 34 39 38
rect 42 38 46 50
rect 61 46 62 47
rect 42 33 46 34
rect 50 43 62 46
rect 66 43 67 47
rect 50 42 67 43
rect 73 46 79 50
rect 91 49 95 50
rect 111 54 115 56
rect 111 47 115 50
rect 73 42 87 46
rect 106 43 111 47
rect 121 49 125 53
rect 121 44 125 45
rect 50 30 54 42
rect 78 38 82 42
rect 64 34 65 38
rect 69 34 75 38
rect 17 29 67 30
rect 3 28 7 29
rect 17 26 23 29
rect 22 25 23 26
rect 27 26 62 29
rect 27 25 28 26
rect 61 25 62 26
rect 66 25 67 29
rect 71 29 75 34
rect 78 33 82 34
rect 91 34 95 35
rect 91 29 95 30
rect 106 29 110 43
rect 114 38 126 39
rect 118 34 126 38
rect 114 33 126 34
rect 71 25 115 29
rect 122 25 126 33
rect 3 21 7 24
rect 12 17 13 21
rect 17 17 33 21
rect 37 17 91 21
rect 95 17 96 21
rect 101 20 105 21
rect 111 20 115 21
rect 121 20 125 21
rect 3 12 7 17
rect 101 12 105 16
rect 121 12 125 16
rect -2 8 44 12
rect 48 8 80 12
rect 84 8 130 12
rect -2 2 130 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 122 2
rect 126 -2 130 2
<< ntransistor >>
rect 9 16 11 30
rect 19 16 21 30
rect 29 16 31 30
rect 39 16 41 30
rect 51 13 53 30
rect 58 13 60 30
rect 68 19 70 30
rect 75 19 77 30
rect 87 12 89 26
rect 97 12 99 26
rect 107 15 109 26
rect 117 15 119 26
<< ptransistor >>
rect 9 42 11 70
rect 19 42 21 70
rect 29 42 31 70
rect 39 42 41 70
rect 51 42 53 70
rect 58 42 60 70
rect 68 42 70 70
rect 75 42 77 70
rect 87 42 89 70
rect 97 42 99 70
rect 107 42 109 70
rect 117 42 119 58
<< polycontact >>
rect 3 34 7 38
rect 26 34 30 38
rect 42 34 46 38
rect 65 34 69 38
rect 78 34 82 38
rect 91 30 95 34
rect 114 34 118 38
<< ndcontact >>
rect 3 24 7 28
rect 3 17 7 21
rect 13 17 17 21
rect 23 25 27 29
rect 33 17 37 21
rect 62 25 66 29
rect 44 8 48 12
rect 91 17 95 21
rect 101 16 105 20
rect 111 21 115 25
rect 121 16 125 20
rect 80 8 84 12
<< pdcontact >>
rect 3 65 7 69
rect 3 58 7 62
rect 13 58 17 62
rect 23 43 27 47
rect 33 58 37 62
rect 44 65 48 69
rect 62 43 66 47
rect 80 65 84 69
rect 91 57 95 61
rect 91 50 95 54
rect 101 65 105 69
rect 101 57 105 61
rect 111 50 115 54
rect 111 43 115 47
rect 121 53 125 57
rect 121 45 125 49
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
rect 90 -2 94 2
rect 98 -2 102 2
rect 106 -2 110 2
rect 114 -2 118 2
rect 122 -2 126 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
rect 90 78 94 82
rect 98 78 102 82
rect 106 78 110 82
rect 114 78 118 82
rect 122 78 126 82
<< psubstratepdiff >>
rect 0 2 128 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 122 2
rect 126 -2 128 2
rect 0 -3 128 -2
<< nsubstratendiff >>
rect 0 82 128 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect 118 78 122 82
rect 126 78 128 82
rect 0 77 128 78
<< labels >>
rlabel polysilicon 64 36 64 36 6 bn
rlabel metal1 20 28 20 28 6 z
rlabel metal1 20 44 20 44 6 z
rlabel metal1 4 40 4 40 6 a
rlabel metal1 12 52 12 52 6 a
rlabel metal1 20 52 20 52 6 a
rlabel metal1 28 28 28 28 6 z
rlabel metal1 36 28 36 28 6 z
rlabel metal1 44 28 44 28 6 z
rlabel polycontact 28 36 28 36 6 c
rlabel metal1 36 40 36 40 6 c
rlabel metal1 28 52 28 52 6 a
rlabel metal1 36 52 36 52 6 a
rlabel metal1 44 52 44 52 6 a
rlabel metal1 64 6 64 6 6 vss
rlabel metal1 60 28 60 28 6 z
rlabel metal1 52 36 52 36 6 z
rlabel metal1 69 36 69 36 6 bn
rlabel metal1 60 44 60 44 6 z
rlabel metal1 60 52 60 52 6 a
rlabel metal1 68 52 68 52 6 a
rlabel metal1 52 52 52 52 6 a
rlabel metal1 64 74 64 74 6 vdd
rlabel metal1 54 19 54 19 6 n3
rlabel metal1 93 30 93 30 6 bn
rlabel metal1 84 44 84 44 6 a
rlabel metal1 93 55 93 55 6 n1
rlabel metal1 76 48 76 48 6 a
rlabel metal1 53 60 53 60 6 n1
rlabel ndcontact 113 24 113 24 6 bn
rlabel metal1 124 32 124 32 6 b
rlabel polycontact 116 36 116 36 6 b
rlabel metal1 113 49 113 49 6 bn
<< end >>
