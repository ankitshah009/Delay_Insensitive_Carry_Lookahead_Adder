magic
tech scmos
timestamp 1180600834
<< checkpaint >>
rect -22 -22 302 122
<< ab >>
rect 0 0 280 100
<< pwell >>
rect -4 -4 284 48
<< nwell >>
rect -4 48 284 104
<< polysilicon >>
rect 27 94 29 98
rect 39 94 41 98
rect 51 94 53 98
rect 59 94 61 98
rect 71 94 73 98
rect 83 94 85 98
rect 91 94 93 98
rect 15 70 17 74
rect 15 53 17 56
rect 7 52 17 53
rect 7 48 8 52
rect 12 48 17 52
rect 7 47 17 48
rect 15 37 17 47
rect 27 53 29 75
rect 39 73 41 76
rect 33 72 41 73
rect 33 68 34 72
rect 38 68 41 72
rect 33 67 41 68
rect 195 94 197 98
rect 207 94 209 98
rect 219 94 221 98
rect 231 94 233 98
rect 243 94 245 98
rect 255 94 257 98
rect 267 94 269 98
rect 121 85 123 89
rect 147 85 149 89
rect 159 85 161 89
rect 171 85 173 89
rect 183 85 185 89
rect 27 52 33 53
rect 27 48 28 52
rect 32 48 33 52
rect 27 47 33 48
rect 15 25 17 29
rect 27 23 29 47
rect 39 41 41 67
rect 51 63 53 75
rect 47 62 53 63
rect 47 58 48 62
rect 52 58 53 62
rect 47 57 53 58
rect 47 52 53 53
rect 47 48 48 52
rect 52 51 53 52
rect 59 51 61 75
rect 71 73 73 76
rect 83 73 85 76
rect 52 49 61 51
rect 52 48 53 49
rect 47 47 53 48
rect 39 39 53 41
rect 33 32 41 33
rect 33 28 34 32
rect 38 28 41 32
rect 33 27 41 28
rect 39 23 41 27
rect 51 23 53 39
rect 59 23 61 49
rect 69 71 73 73
rect 79 71 85 73
rect 69 33 71 71
rect 79 53 81 71
rect 91 63 93 76
rect 103 69 105 73
rect 85 62 93 63
rect 85 58 86 62
rect 90 58 93 62
rect 85 57 93 58
rect 75 52 81 53
rect 75 48 76 52
rect 80 51 81 52
rect 103 51 105 55
rect 121 53 123 65
rect 147 63 149 66
rect 159 63 161 66
rect 171 63 173 66
rect 195 73 197 76
rect 195 72 203 73
rect 195 68 198 72
rect 202 68 203 72
rect 195 67 203 68
rect 141 61 149 63
rect 157 62 163 63
rect 80 49 105 51
rect 80 48 81 49
rect 75 47 81 48
rect 79 39 81 47
rect 65 32 71 33
rect 65 28 66 32
rect 70 28 71 32
rect 65 27 71 28
rect 75 37 81 39
rect 85 42 93 43
rect 85 38 86 42
rect 90 38 93 42
rect 85 37 93 38
rect 103 37 105 49
rect 117 52 123 53
rect 117 48 118 52
rect 122 48 123 52
rect 117 47 123 48
rect 129 52 135 53
rect 129 48 130 52
rect 134 51 135 52
rect 141 51 143 61
rect 157 58 158 62
rect 162 58 163 62
rect 157 57 163 58
rect 169 62 175 63
rect 169 58 170 62
rect 174 58 175 62
rect 169 57 175 58
rect 167 52 173 53
rect 167 51 168 52
rect 134 49 168 51
rect 134 48 135 49
rect 129 47 135 48
rect 75 23 77 37
rect 81 32 87 33
rect 81 28 82 32
rect 86 28 87 32
rect 81 27 87 28
rect 71 21 77 23
rect 71 18 73 21
rect 83 19 85 27
rect 91 19 93 37
rect 103 25 105 29
rect 121 25 123 47
rect 141 29 143 49
rect 167 48 168 49
rect 172 51 173 52
rect 183 51 185 65
rect 207 63 209 75
rect 201 62 209 63
rect 201 58 202 62
rect 206 58 209 62
rect 201 57 209 58
rect 219 51 221 75
rect 231 73 233 76
rect 225 72 233 73
rect 225 68 226 72
rect 230 68 233 72
rect 225 67 233 68
rect 243 53 245 75
rect 243 52 251 53
rect 172 49 233 51
rect 172 48 173 49
rect 167 47 173 48
rect 147 42 153 43
rect 147 38 148 42
rect 152 41 153 42
rect 177 42 185 43
rect 177 41 178 42
rect 152 39 178 41
rect 152 38 153 39
rect 147 37 153 38
rect 177 38 178 39
rect 182 41 185 42
rect 219 42 227 43
rect 219 41 222 42
rect 182 39 222 41
rect 182 38 185 39
rect 177 37 185 38
rect 157 32 163 33
rect 141 27 149 29
rect 157 28 158 32
rect 162 28 163 32
rect 157 27 163 28
rect 169 32 175 33
rect 169 28 170 32
rect 174 28 175 32
rect 169 27 175 28
rect 27 7 29 11
rect 39 7 41 11
rect 51 7 53 11
rect 59 7 61 11
rect 147 24 149 27
rect 159 24 161 27
rect 171 24 173 27
rect 183 25 185 37
rect 219 38 222 39
rect 226 38 227 42
rect 219 37 227 38
rect 201 32 209 33
rect 201 28 202 32
rect 206 28 209 32
rect 201 27 209 28
rect 121 11 123 15
rect 147 11 149 15
rect 71 2 73 6
rect 83 3 85 7
rect 91 3 93 7
rect 159 11 161 15
rect 171 11 173 15
rect 183 11 185 15
rect 195 22 203 23
rect 195 18 198 22
rect 202 18 203 22
rect 195 17 203 18
rect 195 14 197 17
rect 207 15 209 27
rect 219 25 221 37
rect 231 25 233 49
rect 243 48 246 52
rect 250 48 251 52
rect 243 47 251 48
rect 255 43 257 55
rect 267 43 269 55
rect 245 42 269 43
rect 245 38 246 42
rect 250 38 269 42
rect 245 37 269 38
rect 243 32 251 33
rect 243 28 246 32
rect 250 28 251 32
rect 243 27 251 28
rect 243 24 245 27
rect 255 25 257 37
rect 267 25 269 37
rect 219 11 221 15
rect 231 11 233 15
rect 243 11 245 15
rect 195 2 197 6
rect 207 2 209 6
rect 255 2 257 6
rect 267 2 269 6
<< ndiffusion >>
rect 7 29 15 37
rect 17 34 25 37
rect 17 30 20 34
rect 24 30 25 34
rect 17 29 25 30
rect 7 22 13 29
rect 43 32 49 33
rect 43 28 44 32
rect 48 28 49 32
rect 43 23 49 28
rect 7 18 8 22
rect 12 18 13 22
rect 7 17 13 18
rect 19 22 27 23
rect 19 18 20 22
rect 24 18 27 22
rect 19 11 27 18
rect 29 11 39 23
rect 41 11 51 23
rect 53 11 59 23
rect 61 22 69 23
rect 61 18 64 22
rect 68 18 69 22
rect 95 36 103 37
rect 95 32 96 36
rect 100 32 103 36
rect 95 29 103 32
rect 105 29 117 37
rect 107 25 117 29
rect 95 22 101 23
rect 95 19 96 22
rect 78 18 83 19
rect 61 11 71 18
rect 63 6 71 11
rect 73 12 83 18
rect 73 8 76 12
rect 80 8 83 12
rect 73 7 83 8
rect 85 7 91 19
rect 93 18 96 19
rect 100 18 101 22
rect 93 9 101 18
rect 107 15 121 25
rect 123 22 133 25
rect 178 24 183 25
rect 123 18 128 22
rect 132 18 133 22
rect 123 15 133 18
rect 139 22 147 24
rect 139 18 140 22
rect 144 18 147 22
rect 139 15 147 18
rect 149 15 159 24
rect 161 15 171 24
rect 173 22 183 24
rect 173 18 176 22
rect 180 18 183 22
rect 173 15 183 18
rect 185 15 193 25
rect 107 12 117 15
rect 93 7 98 9
rect 107 8 108 12
rect 112 8 117 12
rect 151 12 157 15
rect 107 7 117 8
rect 73 6 80 7
rect 151 8 152 12
rect 156 8 157 12
rect 187 14 193 15
rect 211 22 219 25
rect 211 18 212 22
rect 216 18 219 22
rect 211 15 219 18
rect 221 22 231 25
rect 221 18 224 22
rect 228 18 231 22
rect 221 15 231 18
rect 233 24 238 25
rect 250 24 255 25
rect 233 15 243 24
rect 245 22 255 24
rect 245 18 248 22
rect 252 18 255 22
rect 245 15 255 18
rect 202 14 207 15
rect 151 7 157 8
rect 187 6 195 14
rect 197 12 207 14
rect 197 8 200 12
rect 204 8 207 12
rect 197 6 207 8
rect 209 6 217 15
rect 247 12 255 15
rect 247 8 248 12
rect 252 8 255 12
rect 247 6 255 8
rect 257 22 267 25
rect 257 18 260 22
rect 264 18 267 22
rect 257 6 267 18
rect 269 22 277 25
rect 269 18 272 22
rect 276 18 277 22
rect 269 12 277 18
rect 269 8 272 12
rect 276 8 277 12
rect 269 6 277 8
<< pdiffusion >>
rect 7 82 13 83
rect 7 78 8 82
rect 12 78 13 82
rect 7 70 13 78
rect 19 82 27 94
rect 19 78 20 82
rect 24 78 27 82
rect 19 75 27 78
rect 29 76 39 94
rect 41 76 51 94
rect 29 75 34 76
rect 7 56 15 70
rect 17 62 25 70
rect 17 58 20 62
rect 24 58 25 62
rect 17 56 25 58
rect 43 75 51 76
rect 53 75 59 94
rect 61 82 71 94
rect 61 78 64 82
rect 68 78 71 82
rect 61 76 71 78
rect 73 92 83 94
rect 73 88 76 92
rect 80 88 83 92
rect 73 76 83 88
rect 85 76 91 94
rect 93 82 101 94
rect 93 78 96 82
rect 100 78 101 82
rect 93 76 101 78
rect 107 92 117 93
rect 107 88 108 92
rect 112 88 117 92
rect 151 94 157 95
rect 151 90 152 94
rect 156 90 157 94
rect 107 85 117 88
rect 151 85 157 90
rect 187 85 195 94
rect 61 75 66 76
rect 43 72 49 75
rect 43 68 44 72
rect 48 68 49 72
rect 43 67 49 68
rect 107 69 121 85
rect 95 62 103 69
rect 95 58 96 62
rect 100 58 103 62
rect 95 55 103 58
rect 105 65 121 69
rect 123 72 133 85
rect 123 68 128 72
rect 132 68 133 72
rect 123 65 133 68
rect 139 72 147 85
rect 139 68 140 72
rect 144 68 147 72
rect 139 66 147 68
rect 149 66 159 85
rect 161 66 171 85
rect 173 72 183 85
rect 173 68 176 72
rect 180 68 183 72
rect 173 66 183 68
rect 105 55 117 65
rect 178 65 183 66
rect 185 76 195 85
rect 197 92 207 94
rect 197 88 200 92
rect 204 88 207 92
rect 197 76 207 88
rect 185 65 193 76
rect 202 75 207 76
rect 209 82 219 94
rect 209 78 212 82
rect 216 78 219 82
rect 209 75 219 78
rect 221 82 231 94
rect 221 78 224 82
rect 228 78 231 82
rect 221 76 231 78
rect 233 76 243 94
rect 221 75 226 76
rect 238 75 243 76
rect 245 92 255 94
rect 245 88 248 92
rect 252 88 255 92
rect 245 82 255 88
rect 245 78 248 82
rect 252 78 255 82
rect 245 75 255 78
rect 247 72 255 75
rect 247 68 248 72
rect 252 68 255 72
rect 247 62 255 68
rect 247 58 248 62
rect 252 58 255 62
rect 247 55 255 58
rect 257 82 267 94
rect 257 78 260 82
rect 264 78 267 82
rect 257 72 267 78
rect 257 68 260 72
rect 264 68 267 72
rect 257 62 267 68
rect 257 58 260 62
rect 264 58 267 62
rect 257 55 267 58
rect 269 92 277 94
rect 269 88 272 92
rect 276 88 277 92
rect 269 82 277 88
rect 269 78 272 82
rect 276 78 277 82
rect 269 72 277 78
rect 269 68 272 72
rect 276 68 277 72
rect 269 62 277 68
rect 269 58 272 62
rect 276 58 277 62
rect 269 55 277 58
<< metal1 >>
rect -2 96 282 100
rect -2 92 126 96
rect 130 92 140 96
rect 144 94 164 96
rect 144 92 152 94
rect -2 88 76 92
rect 80 88 108 92
rect 112 90 152 92
rect 156 92 164 94
rect 168 92 176 96
rect 180 92 282 96
rect 156 90 200 92
rect 112 88 200 90
rect 204 88 248 92
rect 252 88 272 92
rect 276 88 282 92
rect 8 82 12 88
rect 96 82 100 83
rect 212 82 216 83
rect 248 82 252 88
rect 19 78 20 82
rect 24 78 64 82
rect 68 78 69 82
rect 100 78 162 82
rect 8 77 12 78
rect 8 72 12 73
rect 96 72 100 78
rect 8 68 34 72
rect 38 68 39 72
rect 43 68 44 72
rect 48 68 112 72
rect 8 52 12 68
rect 8 27 12 48
rect 18 58 20 62
rect 24 58 48 62
rect 52 58 53 62
rect 18 34 22 58
rect 28 52 32 53
rect 39 48 48 52
rect 52 48 53 52
rect 28 41 32 48
rect 58 42 62 68
rect 54 38 62 42
rect 68 52 72 63
rect 86 62 90 63
rect 77 58 86 62
rect 95 58 96 62
rect 100 58 102 62
rect 86 52 90 58
rect 68 48 76 52
rect 80 48 81 52
rect 86 48 93 52
rect 18 30 20 34
rect 24 32 25 34
rect 54 32 58 38
rect 68 37 72 48
rect 86 42 90 48
rect 77 38 86 42
rect 86 37 90 38
rect 98 37 102 58
rect 96 36 102 37
rect 100 32 102 36
rect 24 30 34 32
rect 20 28 34 30
rect 38 28 39 32
rect 43 28 44 32
rect 48 28 58 32
rect 65 28 66 32
rect 70 28 82 32
rect 86 28 100 32
rect 8 22 12 23
rect 108 22 112 68
rect 19 18 20 22
rect 24 18 64 22
rect 68 18 69 22
rect 95 18 96 22
rect 100 18 112 22
rect 118 52 122 73
rect 8 12 12 18
rect 118 17 122 48
rect 128 72 132 73
rect 139 68 140 72
rect 144 71 145 72
rect 144 68 152 71
rect 128 52 132 68
rect 140 67 152 68
rect 128 48 130 52
rect 134 48 135 52
rect 128 22 132 48
rect 148 42 152 67
rect 148 23 152 38
rect 158 62 162 78
rect 223 78 224 82
rect 228 78 240 82
rect 212 72 216 78
rect 175 68 176 72
rect 180 68 192 72
rect 197 68 198 72
rect 202 68 216 72
rect 188 62 192 68
rect 169 58 170 62
rect 174 58 182 62
rect 158 32 162 58
rect 168 52 172 53
rect 168 32 172 48
rect 178 42 182 58
rect 178 37 182 38
rect 188 58 202 62
rect 206 58 207 62
rect 188 32 192 58
rect 168 28 170 32
rect 174 28 175 32
rect 188 28 202 32
rect 206 28 207 32
rect 158 27 162 28
rect 140 22 152 23
rect 188 22 192 28
rect 212 22 216 68
rect 224 68 226 72
rect 230 68 231 72
rect 224 42 228 68
rect 221 38 222 42
rect 226 38 228 42
rect 236 42 240 78
rect 248 72 252 78
rect 248 62 252 68
rect 248 57 252 58
rect 258 82 262 83
rect 272 82 276 88
rect 258 78 260 82
rect 264 78 265 82
rect 258 72 262 78
rect 272 72 276 78
rect 258 68 260 72
rect 264 68 265 72
rect 258 62 262 68
rect 272 62 276 68
rect 258 58 260 62
rect 264 58 265 62
rect 258 52 262 58
rect 272 57 276 58
rect 245 48 246 52
rect 250 48 263 52
rect 236 38 246 42
rect 250 38 251 42
rect 236 22 240 38
rect 258 32 262 48
rect 245 28 246 32
rect 250 28 263 32
rect 139 18 140 22
rect 144 19 152 22
rect 144 18 145 19
rect 175 18 176 22
rect 180 18 192 22
rect 197 18 198 22
rect 202 18 212 22
rect 223 18 224 22
rect 228 18 240 22
rect 248 22 252 23
rect 128 17 132 18
rect 212 17 216 18
rect 248 12 252 18
rect 258 22 262 28
rect 272 22 276 23
rect 258 18 260 22
rect 264 18 265 22
rect 258 17 262 18
rect 272 12 276 18
rect -2 8 76 12
rect 80 8 108 12
rect 112 8 152 12
rect 156 8 200 12
rect 204 8 248 12
rect 252 8 272 12
rect 276 8 282 12
rect -2 4 126 8
rect 130 4 140 8
rect 144 4 164 8
rect 168 4 176 8
rect 180 4 224 8
rect 228 4 236 8
rect 240 4 282 8
rect -2 0 282 4
<< ntransistor >>
rect 15 29 17 37
rect 27 11 29 23
rect 39 11 41 23
rect 51 11 53 23
rect 59 11 61 23
rect 103 29 105 37
rect 71 6 73 18
rect 83 7 85 19
rect 91 7 93 19
rect 121 15 123 25
rect 147 15 149 24
rect 159 15 161 24
rect 171 15 173 24
rect 183 15 185 25
rect 219 15 221 25
rect 231 15 233 25
rect 243 15 245 24
rect 195 6 197 14
rect 207 6 209 15
rect 255 6 257 25
rect 267 6 269 25
<< ptransistor >>
rect 27 75 29 94
rect 39 76 41 94
rect 15 56 17 70
rect 51 75 53 94
rect 59 75 61 94
rect 71 76 73 94
rect 83 76 85 94
rect 91 76 93 94
rect 103 55 105 69
rect 121 65 123 85
rect 147 66 149 85
rect 159 66 161 85
rect 171 66 173 85
rect 183 65 185 85
rect 195 76 197 94
rect 207 75 209 94
rect 219 75 221 94
rect 231 76 233 94
rect 243 75 245 94
rect 255 55 257 94
rect 267 55 269 94
<< polycontact >>
rect 8 48 12 52
rect 34 68 38 72
rect 28 48 32 52
rect 48 58 52 62
rect 48 48 52 52
rect 34 28 38 32
rect 86 58 90 62
rect 76 48 80 52
rect 198 68 202 72
rect 66 28 70 32
rect 86 38 90 42
rect 118 48 122 52
rect 130 48 134 52
rect 158 58 162 62
rect 170 58 174 62
rect 82 28 86 32
rect 168 48 172 52
rect 202 58 206 62
rect 226 68 230 72
rect 148 38 152 42
rect 178 38 182 42
rect 158 28 162 32
rect 170 28 174 32
rect 222 38 226 42
rect 202 28 206 32
rect 198 18 202 22
rect 246 48 250 52
rect 246 38 250 42
rect 246 28 250 32
<< ndcontact >>
rect 20 30 24 34
rect 44 28 48 32
rect 8 18 12 22
rect 20 18 24 22
rect 64 18 68 22
rect 96 32 100 36
rect 76 8 80 12
rect 96 18 100 22
rect 128 18 132 22
rect 140 18 144 22
rect 176 18 180 22
rect 108 8 112 12
rect 152 8 156 12
rect 212 18 216 22
rect 224 18 228 22
rect 248 18 252 22
rect 200 8 204 12
rect 248 8 252 12
rect 260 18 264 22
rect 272 18 276 22
rect 272 8 276 12
<< pdcontact >>
rect 8 78 12 82
rect 20 78 24 82
rect 20 58 24 62
rect 64 78 68 82
rect 76 88 80 92
rect 96 78 100 82
rect 108 88 112 92
rect 152 90 156 94
rect 44 68 48 72
rect 96 58 100 62
rect 128 68 132 72
rect 140 68 144 72
rect 176 68 180 72
rect 200 88 204 92
rect 212 78 216 82
rect 224 78 228 82
rect 248 88 252 92
rect 248 78 252 82
rect 248 68 252 72
rect 248 58 252 62
rect 260 78 264 82
rect 260 68 264 72
rect 260 58 264 62
rect 272 88 276 92
rect 272 78 276 82
rect 272 68 276 72
rect 272 58 276 62
<< psubstratepcontact >>
rect 126 4 130 8
rect 140 4 144 8
rect 164 4 168 8
rect 176 4 180 8
rect 224 4 228 8
rect 236 4 240 8
<< nsubstratencontact >>
rect 126 92 130 96
rect 140 92 144 96
rect 164 92 168 96
rect 176 92 180 96
<< psubstratepdiff >>
rect 125 8 145 9
rect 125 4 126 8
rect 130 4 140 8
rect 144 4 145 8
rect 163 8 181 9
rect 125 3 145 4
rect 163 4 164 8
rect 168 4 176 8
rect 180 4 181 8
rect 223 8 241 9
rect 163 3 181 4
rect 223 4 224 8
rect 228 4 236 8
rect 240 4 241 8
rect 223 3 241 4
<< nsubstratendiff >>
rect 125 96 145 97
rect 125 92 126 96
rect 130 92 140 96
rect 144 92 145 96
rect 163 96 181 97
rect 125 91 145 92
rect 163 92 164 96
rect 168 92 176 96
rect 180 92 181 96
rect 163 91 181 92
<< labels >>
rlabel polycontact 30 50 30 50 6 i2
rlabel polycontact 10 50 10 50 6 cmd1
rlabel metal1 80 40 80 40 6 i0
rlabel polycontact 50 50 50 50 6 i1
rlabel metal1 70 50 70 50 6 cmd0
rlabel metal1 80 60 80 60 6 i0
rlabel metal1 120 45 120 45 6 ck
rlabel metal1 90 50 90 50 6 i0
rlabel metal1 140 6 140 6 6 vss
rlabel metal1 140 94 140 94 6 vdd
rlabel metal1 250 30 250 30 6 q
rlabel metal1 250 50 250 50 6 q
rlabel metal1 260 50 260 50 6 q
<< end >>
