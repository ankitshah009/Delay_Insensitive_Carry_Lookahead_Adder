magic
tech scmos
timestamp 1179386529
<< checkpaint >>
rect -22 -22 62 94
<< ab >>
rect 0 0 40 72
<< pwell >>
rect -4 -4 44 32
<< nwell >>
rect -4 32 44 76
<< polysilicon >>
rect 9 59 11 64
rect 19 59 21 64
rect 29 59 31 64
rect 9 32 11 49
rect 19 43 21 49
rect 19 42 25 43
rect 19 38 20 42
rect 24 38 25 42
rect 19 37 25 38
rect 9 31 17 32
rect 9 27 10 31
rect 14 27 17 31
rect 9 26 17 27
rect 15 23 17 26
rect 22 23 24 37
rect 29 35 31 49
rect 29 34 35 35
rect 29 30 30 34
rect 34 30 35 34
rect 29 29 35 30
rect 29 23 31 29
rect 15 8 17 13
rect 22 8 24 13
rect 29 8 31 13
<< ndiffusion >>
rect 10 19 15 23
rect 8 18 15 19
rect 8 14 9 18
rect 13 14 15 18
rect 8 13 15 14
rect 17 13 22 23
rect 24 13 29 23
rect 31 18 38 23
rect 31 14 33 18
rect 37 14 38 18
rect 31 13 38 14
<< pdiffusion >>
rect 4 55 9 59
rect 2 54 9 55
rect 2 50 3 54
rect 7 50 9 54
rect 2 49 9 50
rect 11 58 19 59
rect 11 54 13 58
rect 17 54 19 58
rect 11 49 19 54
rect 21 54 29 59
rect 21 50 23 54
rect 27 50 29 54
rect 21 49 29 50
rect 31 58 38 59
rect 31 54 33 58
rect 37 54 38 58
rect 31 49 38 54
<< metal1 >>
rect -2 64 42 72
rect 2 54 7 59
rect 12 58 18 64
rect 12 54 13 58
rect 17 54 18 58
rect 32 58 38 64
rect 23 54 27 55
rect 32 54 33 58
rect 37 54 38 58
rect 2 50 3 54
rect 2 46 27 50
rect 2 18 6 46
rect 34 42 38 51
rect 17 38 20 42
rect 24 38 38 42
rect 10 31 14 32
rect 25 30 30 34
rect 10 26 14 27
rect 10 21 23 26
rect 34 21 38 34
rect 2 14 9 18
rect 13 14 14 18
rect 2 13 6 14
rect 18 13 23 21
rect 32 14 33 18
rect 37 14 38 18
rect 32 8 38 14
rect -2 4 4 8
rect 8 4 42 8
rect -2 0 42 4
<< ntransistor >>
rect 15 13 17 23
rect 22 13 24 23
rect 29 13 31 23
<< ptransistor >>
rect 9 49 11 59
rect 19 49 21 59
rect 29 49 31 59
<< polycontact >>
rect 20 38 24 42
rect 10 27 14 31
rect 30 30 34 34
<< ndcontact >>
rect 9 14 13 18
rect 33 14 37 18
<< pdcontact >>
rect 3 50 7 54
rect 13 54 17 58
rect 23 50 27 54
rect 33 54 37 58
<< psubstratepcontact >>
rect 4 4 8 8
<< psubstratepdiff >>
rect 3 8 9 9
rect 3 4 4 8
rect 8 4 9 8
rect 3 3 9 4
<< labels >>
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 24 12 24 6 c
rlabel metal1 12 48 12 48 6 z
rlabel metal1 20 4 20 4 6 vss
rlabel metal1 20 20 20 20 6 c
rlabel metal1 28 32 28 32 6 a
rlabel metal1 28 40 28 40 6 b
rlabel metal1 20 40 20 40 6 b
rlabel metal1 20 48 20 48 6 z
rlabel metal1 20 68 20 68 6 vdd
rlabel metal1 36 24 36 24 6 a
rlabel metal1 36 48 36 48 6 b
<< end >>
