magic
tech scmos
timestamp 1179387360
<< checkpaint >>
rect -22 -22 54 94
<< ab >>
rect 0 0 32 72
<< pwell >>
rect -4 -4 36 32
<< nwell >>
rect -4 32 36 76
<< metal1 >>
rect -2 68 34 72
rect -2 64 7 68
rect 11 64 14 68
rect 18 64 21 68
rect 25 64 34 68
rect -2 4 7 8
rect 11 4 14 8
rect 18 4 21 8
rect 25 4 34 8
rect -2 0 34 4
<< psubstratepcontact >>
rect 7 4 11 8
rect 14 4 18 8
rect 21 4 25 8
<< nsubstratencontact >>
rect 7 64 11 68
rect 14 64 18 68
rect 21 64 25 68
<< psubstratepdiff >>
rect 6 8 26 26
rect 6 4 7 8
rect 11 4 14 8
rect 18 4 21 8
rect 25 4 26 8
rect 6 3 26 4
<< nsubstratendiff >>
rect 6 68 26 69
rect 6 64 7 68
rect 11 64 14 68
rect 18 64 21 68
rect 25 64 26 68
rect 6 38 26 64
<< labels >>
rlabel metal1 16 4 16 4 6 vss
rlabel metal1 16 68 16 68 6 vdd
<< end >>
