magic
tech scmos
timestamp 1180600691
<< checkpaint >>
rect -22 -22 82 122
<< ab >>
rect 0 0 60 100
<< pwell >>
rect -4 -4 64 48
<< nwell >>
rect -4 48 64 104
<< polysilicon >>
rect 11 94 13 98
rect 23 94 25 98
rect 35 94 37 98
rect 11 43 13 55
rect 23 43 25 55
rect 7 42 13 43
rect 7 38 8 42
rect 12 38 13 42
rect 7 37 13 38
rect 17 42 25 43
rect 17 38 18 42
rect 22 38 25 42
rect 17 37 25 38
rect 11 25 13 37
rect 23 25 25 37
rect 35 43 37 55
rect 35 42 43 43
rect 35 38 38 42
rect 42 38 43 42
rect 35 37 43 38
rect 35 25 37 37
rect 11 2 13 6
rect 23 2 25 6
rect 35 2 37 6
<< ndiffusion >>
rect 15 32 21 33
rect 15 28 16 32
rect 20 28 21 32
rect 15 25 21 28
rect 3 22 11 25
rect 3 18 4 22
rect 8 18 11 22
rect 3 6 11 18
rect 13 6 23 25
rect 25 22 35 25
rect 25 18 28 22
rect 32 18 35 22
rect 25 6 35 18
rect 37 12 45 25
rect 37 8 40 12
rect 44 8 45 12
rect 37 6 45 8
<< pdiffusion >>
rect 3 92 11 94
rect 3 88 4 92
rect 8 88 11 92
rect 3 55 11 88
rect 13 55 23 94
rect 25 82 35 94
rect 25 78 28 82
rect 32 78 35 82
rect 25 72 35 78
rect 25 68 28 72
rect 32 68 35 72
rect 25 62 35 68
rect 25 58 28 62
rect 32 58 35 62
rect 25 55 35 58
rect 37 92 45 94
rect 37 88 40 92
rect 44 88 45 92
rect 37 55 45 88
<< metal1 >>
rect -2 96 62 100
rect -2 92 52 96
rect 56 92 62 96
rect -2 88 4 92
rect 8 88 40 92
rect 44 88 62 92
rect 8 42 12 83
rect 8 37 12 38
rect 18 42 22 83
rect 18 37 22 38
rect 28 82 32 83
rect 28 72 32 78
rect 28 62 32 68
rect 28 32 32 58
rect 15 28 16 32
rect 20 28 32 32
rect 28 27 32 28
rect 38 42 42 83
rect 52 60 56 88
rect 52 55 56 56
rect 3 18 4 22
rect 8 18 28 22
rect 32 18 33 22
rect 38 17 42 38
rect 52 36 56 37
rect 52 12 56 32
rect -2 8 40 12
rect 44 8 62 12
rect -2 4 52 8
rect 56 4 62 8
rect -2 0 62 4
<< ntransistor >>
rect 11 6 13 25
rect 23 6 25 25
rect 35 6 37 25
<< ptransistor >>
rect 11 55 13 94
rect 23 55 25 94
rect 35 55 37 94
<< polycontact >>
rect 8 38 12 42
rect 18 38 22 42
rect 38 38 42 42
<< ndcontact >>
rect 16 28 20 32
rect 4 18 8 22
rect 28 18 32 22
rect 40 8 44 12
<< pdcontact >>
rect 4 88 8 92
rect 28 78 32 82
rect 28 68 32 72
rect 28 58 32 62
rect 40 88 44 92
<< psubstratepcontact >>
rect 52 32 56 36
rect 52 4 56 8
<< nsubstratencontact >>
rect 52 92 56 96
rect 52 56 56 60
<< psubstratepdiff >>
rect 51 36 57 37
rect 51 32 52 36
rect 56 32 57 36
rect 51 26 57 32
rect 51 8 57 14
rect 51 4 52 8
rect 56 4 57 8
rect 51 3 57 4
<< nsubstratendiff >>
rect 51 96 57 97
rect 51 92 52 96
rect 56 92 57 96
rect 51 86 57 92
rect 51 60 57 66
rect 51 56 52 60
rect 56 56 57 60
rect 51 55 57 56
<< labels >>
rlabel metal1 10 60 10 60 6 i0
rlabel metal1 20 30 20 30 6 nq
rlabel metal1 20 60 20 60 6 i1
rlabel metal1 30 6 30 6 6 vss
rlabel metal1 40 50 40 50 6 i2
rlabel metal1 30 55 30 55 6 nq
rlabel metal1 30 94 30 94 6 vdd
<< end >>
