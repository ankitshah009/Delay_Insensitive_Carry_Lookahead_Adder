magic
tech scmos
timestamp 1179387681
<< checkpaint >>
rect -22 -25 94 105
<< ab >>
rect 0 0 72 80
<< pwell >>
rect -4 -7 76 36
<< nwell >>
rect -4 36 76 87
<< polysilicon >>
rect 38 67 63 69
rect 28 63 34 64
rect 28 59 29 63
rect 33 59 34 63
rect 18 54 20 59
rect 28 58 34 59
rect 28 54 30 58
rect 38 54 40 67
rect 61 63 63 67
rect 48 54 50 59
rect 18 39 20 42
rect 9 38 20 39
rect 9 34 10 38
rect 14 37 20 38
rect 14 34 15 37
rect 9 33 15 34
rect 28 34 30 42
rect 38 38 40 42
rect 48 38 50 42
rect 61 39 63 51
rect 57 38 63 39
rect 47 37 53 38
rect 47 34 48 37
rect 12 29 14 33
rect 22 29 24 33
rect 28 32 34 34
rect 32 29 34 32
rect 42 33 48 34
rect 52 33 53 37
rect 57 34 58 38
rect 62 34 63 38
rect 57 33 63 34
rect 42 32 53 33
rect 42 29 44 32
rect 61 29 63 33
rect 12 18 14 23
rect 22 15 24 23
rect 32 19 34 23
rect 42 19 44 23
rect 61 15 63 23
rect 22 13 63 15
<< ndiffusion >>
rect 4 23 12 29
rect 14 28 22 29
rect 14 24 16 28
rect 20 24 22 28
rect 14 23 22 24
rect 24 28 32 29
rect 24 24 26 28
rect 30 24 32 28
rect 24 23 32 24
rect 34 28 42 29
rect 34 24 36 28
rect 40 24 42 28
rect 34 23 42 24
rect 44 28 61 29
rect 44 24 55 28
rect 59 24 61 28
rect 44 23 61 24
rect 63 28 70 29
rect 63 24 65 28
rect 69 24 70 28
rect 63 23 70 24
rect 4 21 10 23
rect 4 17 5 21
rect 9 17 10 21
rect 4 16 10 17
<< pdiffusion >>
rect 52 64 59 65
rect 52 60 54 64
rect 58 63 59 64
rect 58 60 61 63
rect 52 54 61 60
rect 8 53 18 54
rect 8 49 10 53
rect 14 49 18 53
rect 8 42 18 49
rect 20 47 28 54
rect 20 43 22 47
rect 26 43 28 47
rect 20 42 28 43
rect 30 47 38 54
rect 30 43 32 47
rect 36 43 38 47
rect 30 42 38 43
rect 40 47 48 54
rect 40 43 42 47
rect 46 43 48 47
rect 40 42 48 43
rect 50 51 61 54
rect 63 57 68 63
rect 63 56 70 57
rect 63 52 65 56
rect 69 52 70 56
rect 63 51 70 52
rect 50 42 59 51
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect -2 68 74 78
rect 10 53 14 68
rect 53 64 59 68
rect 28 59 29 63
rect 33 59 49 63
rect 53 60 54 64
rect 58 60 59 64
rect 45 56 49 59
rect 10 48 14 49
rect 34 48 38 55
rect 45 52 65 56
rect 69 52 70 56
rect 32 47 38 48
rect 17 43 22 47
rect 26 43 27 47
rect 36 43 38 47
rect 2 38 14 39
rect 2 34 10 38
rect 2 33 14 34
rect 2 25 6 33
rect 17 29 21 43
rect 32 41 38 43
rect 41 47 46 48
rect 41 43 42 47
rect 41 42 46 43
rect 32 38 36 41
rect 16 28 21 29
rect 20 24 21 28
rect 25 34 36 38
rect 25 28 31 34
rect 41 28 45 42
rect 50 41 62 47
rect 58 38 62 41
rect 25 24 26 28
rect 30 24 31 28
rect 35 24 36 28
rect 40 24 45 28
rect 48 37 52 38
rect 58 33 62 34
rect 16 23 21 24
rect 17 21 21 23
rect 48 21 52 33
rect 66 29 70 52
rect 4 17 5 21
rect 9 17 10 21
rect 17 17 52 21
rect 55 28 59 29
rect 4 12 10 17
rect 55 12 59 24
rect 65 28 70 29
rect 69 24 70 28
rect 65 23 70 24
rect -2 2 74 12
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
<< ntransistor >>
rect 12 23 14 29
rect 22 23 24 29
rect 32 23 34 29
rect 42 23 44 29
rect 61 23 63 29
<< ptransistor >>
rect 18 42 20 54
rect 28 42 30 54
rect 38 42 40 54
rect 48 42 50 54
rect 61 51 63 63
<< polycontact >>
rect 29 59 33 63
rect 10 34 14 38
rect 48 33 52 37
rect 58 34 62 38
<< ndcontact >>
rect 16 24 20 28
rect 26 24 30 28
rect 36 24 40 28
rect 55 24 59 28
rect 65 24 69 28
rect 5 17 9 21
<< pdcontact >>
rect 54 60 58 64
rect 10 49 14 53
rect 22 43 26 47
rect 32 43 36 47
rect 42 43 46 47
rect 65 52 69 56
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
<< psubstratepdiff >>
rect 0 2 72 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 72 2
rect 0 -3 72 -2
<< nsubstratendiff >>
rect 0 82 72 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 72 82
rect 0 77 72 78
<< labels >>
rlabel polycontact 31 61 31 61 6 bn
rlabel ptransistor 49 45 49 45 6 an
rlabel metal1 4 32 4 32 6 a
rlabel metal1 19 32 19 32 6 an
rlabel polycontact 12 36 12 36 6 a
rlabel metal1 22 45 22 45 6 an
rlabel metal1 36 6 36 6 6 vss
rlabel metal1 28 32 28 32 6 z
rlabel metal1 36 48 36 48 6 z
rlabel metal1 36 74 36 74 6 vdd
rlabel metal1 40 26 40 26 6 ai
rlabel metal1 50 27 50 27 6 an
rlabel metal1 52 44 52 44 6 b
rlabel metal1 43 36 43 36 6 ai
rlabel metal1 38 61 38 61 6 bn
rlabel metal1 60 40 60 40 6 b
rlabel metal1 68 39 68 39 6 bn
rlabel metal1 57 54 57 54 6 bn
<< end >>
