magic
tech scmos
timestamp 1180600627
<< checkpaint >>
rect -22 -22 102 122
<< ab >>
rect 0 0 80 100
<< pwell >>
rect -4 -4 84 48
<< nwell >>
rect -4 48 84 104
<< polysilicon >>
rect 53 94 55 98
rect 65 94 67 98
rect 11 85 13 89
rect 23 85 25 89
rect 35 85 37 89
rect 11 43 13 65
rect 23 63 25 66
rect 17 62 25 63
rect 17 58 18 62
rect 22 61 25 62
rect 22 58 23 61
rect 17 57 23 58
rect 35 53 37 65
rect 35 52 43 53
rect 35 51 38 52
rect 37 48 38 51
rect 42 48 43 52
rect 37 47 43 48
rect 27 46 33 47
rect 7 42 13 43
rect 7 38 8 42
rect 12 38 13 42
rect 7 37 13 38
rect 11 25 13 37
rect 17 42 23 43
rect 17 38 18 42
rect 22 38 23 42
rect 27 42 28 46
rect 32 43 33 46
rect 53 43 55 55
rect 65 43 67 55
rect 32 42 67 43
rect 27 41 67 42
rect 17 37 23 38
rect 17 35 25 37
rect 23 25 25 35
rect 37 32 43 33
rect 37 29 38 32
rect 35 28 38 29
rect 42 28 43 32
rect 35 27 43 28
rect 35 24 37 27
rect 53 25 55 41
rect 65 25 67 41
rect 11 11 13 15
rect 23 11 25 15
rect 35 11 37 15
rect 53 2 55 6
rect 65 2 67 6
<< ndiffusion >>
rect 15 32 21 33
rect 15 28 16 32
rect 20 28 21 32
rect 15 25 21 28
rect 3 22 11 25
rect 3 18 4 22
rect 8 18 11 22
rect 3 15 11 18
rect 13 15 23 25
rect 25 24 30 25
rect 44 24 53 25
rect 25 22 35 24
rect 25 18 28 22
rect 32 18 35 22
rect 25 15 35 18
rect 37 15 53 24
rect 39 12 53 15
rect 39 8 44 12
rect 48 8 53 12
rect 39 6 53 8
rect 55 22 65 25
rect 55 18 58 22
rect 62 18 65 22
rect 55 6 65 18
rect 67 22 75 25
rect 67 18 70 22
rect 74 18 75 22
rect 67 12 75 18
rect 67 8 70 12
rect 74 8 75 12
rect 67 6 75 8
<< pdiffusion >>
rect 3 92 9 93
rect 3 88 4 92
rect 8 88 9 92
rect 39 92 53 94
rect 3 85 9 88
rect 39 88 44 92
rect 48 88 53 92
rect 39 85 53 88
rect 3 65 11 85
rect 13 66 23 85
rect 25 82 35 85
rect 25 78 28 82
rect 32 78 35 82
rect 25 72 35 78
rect 25 68 28 72
rect 32 68 35 72
rect 25 66 35 68
rect 13 65 18 66
rect 30 65 35 66
rect 37 65 53 85
rect 39 55 53 65
rect 55 82 65 94
rect 55 78 58 82
rect 62 78 65 82
rect 55 72 65 78
rect 55 68 58 72
rect 62 68 65 72
rect 55 62 65 68
rect 55 58 58 62
rect 62 58 65 62
rect 55 55 65 58
rect 67 92 75 94
rect 67 88 70 92
rect 74 88 75 92
rect 67 82 75 88
rect 67 78 70 82
rect 74 78 75 82
rect 67 72 75 78
rect 67 68 70 72
rect 74 68 75 72
rect 67 62 75 68
rect 67 58 70 62
rect 74 58 75 62
rect 67 55 75 58
<< metal1 >>
rect -2 96 82 100
rect -2 92 16 96
rect 20 92 28 96
rect 32 92 82 96
rect -2 88 4 92
rect 8 88 44 92
rect 48 88 70 92
rect 74 88 82 92
rect 8 42 12 83
rect 8 37 12 38
rect 18 62 22 83
rect 18 42 22 58
rect 18 37 22 38
rect 28 82 32 83
rect 28 72 32 78
rect 28 46 32 68
rect 28 32 32 42
rect 15 28 16 32
rect 20 28 32 32
rect 38 52 42 83
rect 38 32 42 48
rect 3 18 4 22
rect 8 18 28 22
rect 32 18 33 22
rect 38 17 42 28
rect 58 82 62 83
rect 58 72 62 78
rect 58 62 62 68
rect 58 22 62 58
rect 70 82 74 88
rect 70 72 74 78
rect 70 62 74 68
rect 70 57 74 58
rect 58 17 62 18
rect 70 22 74 23
rect 70 12 74 18
rect -2 8 44 12
rect 48 8 70 12
rect 74 8 82 12
rect -2 4 4 8
rect 8 4 16 8
rect 20 4 28 8
rect 32 4 82 8
rect -2 0 82 4
<< ntransistor >>
rect 11 15 13 25
rect 23 15 25 25
rect 35 15 37 24
rect 53 6 55 25
rect 65 6 67 25
<< ptransistor >>
rect 11 65 13 85
rect 23 66 25 85
rect 35 65 37 85
rect 53 55 55 94
rect 65 55 67 94
<< polycontact >>
rect 18 58 22 62
rect 38 48 42 52
rect 8 38 12 42
rect 18 38 22 42
rect 28 42 32 46
rect 38 28 42 32
<< ndcontact >>
rect 16 28 20 32
rect 4 18 8 22
rect 28 18 32 22
rect 44 8 48 12
rect 58 18 62 22
rect 70 18 74 22
rect 70 8 74 12
<< pdcontact >>
rect 4 88 8 92
rect 44 88 48 92
rect 28 78 32 82
rect 28 68 32 72
rect 58 78 62 82
rect 58 68 62 72
rect 58 58 62 62
rect 70 88 74 92
rect 70 78 74 82
rect 70 68 74 72
rect 70 58 74 62
<< psubstratepcontact >>
rect 4 4 8 8
rect 16 4 20 8
rect 28 4 32 8
<< nsubstratencontact >>
rect 16 92 20 96
rect 28 92 32 96
<< psubstratepdiff >>
rect 3 8 33 9
rect 3 4 4 8
rect 8 4 16 8
rect 20 4 28 8
rect 32 4 33 8
rect 3 3 33 4
<< nsubstratendiff >>
rect 15 96 33 97
rect 15 92 16 96
rect 20 92 28 96
rect 32 92 33 96
rect 15 91 33 92
<< labels >>
rlabel metal1 10 60 10 60 6 i0
rlabel polycontact 20 60 20 60 6 i1
rlabel metal1 40 6 40 6 6 vss
rlabel polycontact 40 50 40 50 6 i2
rlabel metal1 40 94 40 94 6 vdd
rlabel metal1 60 50 60 50 6 q
<< end >>
