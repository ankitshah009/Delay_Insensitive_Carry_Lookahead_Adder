magic
tech scmos
timestamp 1185039039
<< checkpaint >>
rect -22 -24 82 124
<< ab >>
rect 0 0 60 100
<< pwell >>
rect -2 -4 62 49
<< nwell >>
rect -2 49 62 104
<< polysilicon >>
rect 19 95 21 98
rect 27 95 29 98
rect 35 95 37 98
rect 43 95 45 98
rect 19 53 21 55
rect 17 52 23 53
rect 17 49 18 52
rect 11 48 18 49
rect 22 48 23 52
rect 11 47 23 48
rect 11 25 13 47
rect 27 43 29 55
rect 35 53 37 55
rect 43 53 45 55
rect 35 51 39 53
rect 43 51 49 53
rect 27 42 33 43
rect 27 39 28 42
rect 23 38 28 39
rect 32 38 33 42
rect 23 37 33 38
rect 23 25 25 37
rect 37 33 39 51
rect 47 43 49 51
rect 47 42 53 43
rect 47 38 48 42
rect 52 38 53 42
rect 47 37 53 38
rect 37 32 43 33
rect 37 29 38 32
rect 35 28 38 29
rect 42 28 43 32
rect 35 27 43 28
rect 35 25 37 27
rect 47 25 49 37
rect 11 12 13 15
rect 23 12 25 15
rect 35 12 37 15
rect 47 12 49 15
<< ndiffusion >>
rect 3 15 11 25
rect 13 22 23 25
rect 13 18 16 22
rect 20 18 23 22
rect 13 15 23 18
rect 25 15 35 25
rect 37 22 47 25
rect 37 18 40 22
rect 44 18 47 22
rect 37 15 47 18
rect 49 15 57 25
rect 3 12 9 15
rect 27 12 33 15
rect 51 12 57 15
rect 3 8 4 12
rect 8 8 9 12
rect 3 7 9 8
rect 27 8 28 12
rect 32 8 33 12
rect 27 7 33 8
rect 51 8 52 12
rect 56 8 57 12
rect 51 5 57 8
<< pdiffusion >>
rect 15 85 19 95
rect 7 82 19 85
rect 7 78 8 82
rect 12 78 19 82
rect 7 72 19 78
rect 7 68 8 72
rect 12 68 19 72
rect 7 62 19 68
rect 7 58 8 62
rect 12 58 19 62
rect 7 55 19 58
rect 21 55 27 95
rect 29 55 35 95
rect 37 55 43 95
rect 45 92 53 95
rect 45 88 48 92
rect 52 88 53 92
rect 45 55 53 88
<< metal1 >>
rect -2 92 62 101
rect -2 88 48 92
rect 52 88 62 92
rect -2 87 62 88
rect 7 82 13 83
rect 7 78 8 82
rect 12 78 13 82
rect 7 72 13 78
rect 7 68 8 72
rect 12 68 13 72
rect 7 62 13 68
rect 7 58 8 62
rect 12 58 13 62
rect 7 23 13 58
rect 17 52 23 82
rect 17 48 18 52
rect 22 48 23 52
rect 17 28 23 48
rect 27 42 33 82
rect 27 38 28 42
rect 32 38 33 42
rect 27 28 33 38
rect 37 32 43 82
rect 37 28 38 32
rect 42 28 43 32
rect 47 42 53 82
rect 47 38 48 42
rect 52 38 53 42
rect 47 28 53 38
rect 37 27 43 28
rect 7 22 45 23
rect 7 18 16 22
rect 20 18 40 22
rect 44 18 45 22
rect 7 17 45 18
rect -2 12 62 13
rect -2 8 4 12
rect 8 8 28 12
rect 32 8 52 12
rect 56 8 62 12
rect -2 -1 62 8
<< ntransistor >>
rect 11 15 13 25
rect 23 15 25 25
rect 35 15 37 25
rect 47 15 49 25
<< ptransistor >>
rect 19 55 21 95
rect 27 55 29 95
rect 35 55 37 95
rect 43 55 45 95
<< polycontact >>
rect 18 48 22 52
rect 28 38 32 42
rect 48 38 52 42
rect 38 28 42 32
<< ndcontact >>
rect 16 18 20 22
rect 40 18 44 22
rect 4 8 8 12
rect 28 8 32 12
rect 52 8 56 12
<< pdcontact >>
rect 8 78 12 82
rect 8 68 12 72
rect 8 58 12 62
rect 48 88 52 92
<< labels >>
rlabel metal1 10 50 10 50 6 nq
rlabel metal1 10 50 10 50 6 nq
rlabel metal1 20 55 20 55 6 i1
rlabel metal1 20 55 20 55 6 i1
rlabel metal1 30 6 30 6 6 vss
rlabel metal1 30 6 30 6 6 vss
rlabel metal1 30 55 30 55 6 i0
rlabel metal1 30 55 30 55 6 i0
rlabel metal1 40 55 40 55 6 i2
rlabel metal1 40 55 40 55 6 i2
rlabel metal1 30 94 30 94 6 vdd
rlabel metal1 30 94 30 94 6 vdd
rlabel metal1 50 55 50 55 6 i3
rlabel metal1 50 55 50 55 6 i3
<< end >>
