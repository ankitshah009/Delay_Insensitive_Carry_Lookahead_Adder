magic
tech scmos
timestamp 1179386483
<< checkpaint >>
rect -22 -22 94 94
<< ab >>
rect 0 0 72 72
<< pwell >>
rect -4 -4 76 32
<< nwell >>
rect -4 32 76 76
<< polysilicon >>
rect 9 65 11 70
rect 19 65 21 70
rect 29 65 31 70
rect 39 65 41 70
rect 49 65 51 70
rect 59 65 61 70
rect 9 35 11 38
rect 19 35 21 38
rect 29 35 31 38
rect 39 35 41 38
rect 49 35 51 38
rect 59 35 61 38
rect 9 34 15 35
rect 9 30 10 34
rect 14 30 15 34
rect 9 29 15 30
rect 19 34 33 35
rect 19 30 26 34
rect 30 30 33 34
rect 19 29 33 30
rect 12 26 14 29
rect 19 26 21 29
rect 31 26 33 29
rect 38 34 51 35
rect 38 30 42 34
rect 46 30 51 34
rect 38 29 51 30
rect 55 34 61 35
rect 55 30 56 34
rect 60 30 61 34
rect 55 29 61 30
rect 38 26 40 29
rect 48 26 50 29
rect 55 26 57 29
rect 12 11 14 15
rect 19 10 21 15
rect 31 2 33 6
rect 38 2 40 6
rect 48 2 50 6
rect 55 2 57 6
<< ndiffusion >>
rect 5 25 12 26
rect 5 21 6 25
rect 10 21 12 25
rect 5 20 12 21
rect 7 15 12 20
rect 14 15 19 26
rect 21 15 31 26
rect 23 11 31 15
rect 23 7 24 11
rect 28 7 31 11
rect 23 6 31 7
rect 33 6 38 26
rect 40 18 48 26
rect 40 14 42 18
rect 46 14 48 18
rect 40 6 48 14
rect 50 6 55 26
rect 57 8 66 26
rect 57 6 60 8
rect 59 4 60 6
rect 64 4 66 8
rect 59 3 66 4
<< pdiffusion >>
rect 2 64 9 65
rect 2 60 3 64
rect 7 60 9 64
rect 2 57 9 60
rect 2 53 3 57
rect 7 53 9 57
rect 2 38 9 53
rect 11 58 19 65
rect 11 54 13 58
rect 17 54 19 58
rect 11 50 19 54
rect 11 46 13 50
rect 17 46 19 50
rect 11 38 19 46
rect 21 64 29 65
rect 21 60 23 64
rect 27 60 29 64
rect 21 57 29 60
rect 21 53 23 57
rect 27 53 29 57
rect 21 38 29 53
rect 31 58 39 65
rect 31 54 33 58
rect 37 54 39 58
rect 31 50 39 54
rect 31 46 33 50
rect 37 46 39 50
rect 31 38 39 46
rect 41 64 49 65
rect 41 60 43 64
rect 47 60 49 64
rect 41 57 49 60
rect 41 53 43 57
rect 47 53 49 57
rect 41 38 49 53
rect 51 58 59 65
rect 51 54 53 58
rect 57 54 59 58
rect 51 51 59 54
rect 51 47 53 51
rect 57 47 59 51
rect 51 38 59 47
rect 61 64 68 65
rect 61 60 63 64
rect 67 60 68 64
rect 61 57 68 60
rect 61 53 63 57
rect 67 53 68 57
rect 61 38 68 53
<< metal1 >>
rect -2 64 74 72
rect 2 60 3 64
rect 7 60 8 64
rect 2 57 8 60
rect 22 60 23 64
rect 27 60 28 64
rect 2 53 3 57
rect 7 53 8 57
rect 13 58 17 59
rect 13 50 17 54
rect 22 57 28 60
rect 42 60 43 64
rect 47 60 48 64
rect 22 53 23 57
rect 27 53 28 57
rect 33 58 38 59
rect 37 54 38 58
rect 33 50 38 54
rect 42 57 48 60
rect 62 60 63 64
rect 67 60 68 64
rect 42 53 43 57
rect 47 53 48 57
rect 53 58 57 59
rect 53 51 57 54
rect 62 57 68 60
rect 62 53 63 57
rect 67 53 68 57
rect 2 46 13 50
rect 17 46 33 50
rect 37 47 53 50
rect 57 47 63 50
rect 37 46 63 47
rect 2 21 6 46
rect 25 38 63 42
rect 10 34 21 35
rect 14 30 21 34
rect 25 34 31 38
rect 55 34 61 38
rect 25 30 26 34
rect 30 30 31 34
rect 41 30 42 34
rect 46 30 47 34
rect 55 30 56 34
rect 60 30 61 34
rect 10 29 21 30
rect 17 26 21 29
rect 41 26 47 30
rect 10 21 11 25
rect 17 22 55 26
rect 7 18 11 21
rect 7 14 42 18
rect 46 14 47 18
rect 23 8 24 11
rect -2 4 4 8
rect 8 4 12 8
rect 16 7 24 8
rect 28 8 29 11
rect 28 7 60 8
rect 16 4 60 7
rect 64 4 74 8
rect -2 0 74 4
<< ntransistor >>
rect 12 15 14 26
rect 19 15 21 26
rect 31 6 33 26
rect 38 6 40 26
rect 48 6 50 26
rect 55 6 57 26
<< ptransistor >>
rect 9 38 11 65
rect 19 38 21 65
rect 29 38 31 65
rect 39 38 41 65
rect 49 38 51 65
rect 59 38 61 65
<< polycontact >>
rect 10 30 14 34
rect 26 30 30 34
rect 42 30 46 34
rect 56 30 60 34
<< ndcontact >>
rect 6 21 10 25
rect 24 7 28 11
rect 42 14 46 18
rect 60 4 64 8
<< pdcontact >>
rect 3 60 7 64
rect 3 53 7 57
rect 13 54 17 58
rect 13 46 17 50
rect 23 60 27 64
rect 23 53 27 57
rect 33 54 37 58
rect 33 46 37 50
rect 43 60 47 64
rect 43 53 47 57
rect 53 54 57 58
rect 53 47 57 51
rect 63 60 67 64
rect 63 53 67 57
<< psubstratepcontact >>
rect 4 4 8 8
rect 12 4 16 8
<< psubstratepdiff >>
rect 3 8 17 9
rect 3 4 4 8
rect 8 4 12 8
rect 16 4 17 8
rect 3 3 17 4
<< labels >>
rlabel metal1 4 32 4 32 6 z
rlabel metal1 20 16 20 16 6 z
rlabel metal1 12 16 12 16 6 z
rlabel metal1 20 24 20 24 6 b
rlabel polycontact 12 32 12 32 6 b
rlabel metal1 12 48 12 48 6 z
rlabel metal1 20 48 20 48 6 z
rlabel metal1 36 4 36 4 6 vss
rlabel metal1 36 16 36 16 6 z
rlabel metal1 28 16 28 16 6 z
rlabel metal1 28 24 28 24 6 b
rlabel metal1 36 24 36 24 6 b
rlabel metal1 28 36 28 36 6 a
rlabel metal1 36 40 36 40 6 a
rlabel metal1 28 48 28 48 6 z
rlabel metal1 36 52 36 52 6 z
rlabel metal1 36 68 36 68 6 vdd
rlabel ndcontact 44 16 44 16 6 z
rlabel metal1 52 24 52 24 6 b
rlabel metal1 44 28 44 28 6 b
rlabel metal1 44 40 44 40 6 a
rlabel metal1 52 40 52 40 6 a
rlabel metal1 44 48 44 48 6 z
rlabel metal1 52 48 52 48 6 z
rlabel metal1 60 40 60 40 6 a
rlabel metal1 60 48 60 48 6 z
<< end >>
