magic
tech scmos
timestamp 1179387809
<< checkpaint >>
rect -22 -22 150 94
<< ab >>
rect 0 0 128 72
<< pwell >>
rect -4 -4 132 32
<< nwell >>
rect -4 32 132 76
<< polysilicon >>
rect 9 66 11 70
rect 19 66 21 70
rect 29 66 31 70
rect 39 66 41 70
rect 49 66 51 70
rect 69 66 71 70
rect 79 66 81 70
rect 89 66 91 70
rect 39 49 41 52
rect 49 49 51 52
rect 39 48 51 49
rect 39 47 46 48
rect 45 44 46 47
rect 50 44 51 48
rect 45 43 51 44
rect 100 60 116 61
rect 100 59 111 60
rect 100 56 102 59
rect 110 56 111 59
rect 115 56 116 60
rect 110 55 116 56
rect 110 52 112 55
rect 100 38 102 42
rect 9 35 11 38
rect 19 35 21 38
rect 29 35 31 38
rect 69 35 71 38
rect 79 35 81 38
rect 9 34 15 35
rect 9 30 10 34
rect 14 30 15 34
rect 9 29 15 30
rect 19 34 25 35
rect 19 30 20 34
rect 24 30 25 34
rect 29 34 65 35
rect 29 33 60 34
rect 19 29 25 30
rect 10 20 12 29
rect 19 25 21 29
rect 37 25 39 33
rect 59 30 60 33
rect 64 30 65 34
rect 59 29 65 30
rect 69 34 75 35
rect 69 30 70 34
rect 74 30 75 34
rect 69 29 75 30
rect 79 34 85 35
rect 79 30 80 34
rect 84 30 85 34
rect 89 34 91 38
rect 89 33 103 34
rect 89 32 98 33
rect 79 29 85 30
rect 97 29 98 32
rect 102 29 103 33
rect 49 28 55 29
rect 17 23 21 25
rect 17 20 19 23
rect 27 20 29 25
rect 49 24 50 28
rect 54 24 55 28
rect 49 23 55 24
rect 49 20 51 23
rect 72 20 74 29
rect 79 20 81 29
rect 97 28 103 29
rect 99 25 101 28
rect 110 26 112 38
rect 89 20 91 25
rect 37 8 39 12
rect 10 2 12 7
rect 17 2 19 7
rect 27 4 29 7
rect 49 4 51 9
rect 27 2 51 4
rect 99 8 101 12
rect 72 2 74 7
rect 79 2 81 7
rect 89 4 91 7
rect 110 4 112 15
rect 89 2 112 4
<< ndiffusion >>
rect 32 20 37 25
rect 2 8 10 20
rect 2 4 3 8
rect 7 7 10 8
rect 12 7 17 20
rect 19 18 27 20
rect 19 14 21 18
rect 25 14 27 18
rect 19 7 27 14
rect 29 19 37 20
rect 29 15 31 19
rect 35 15 37 19
rect 29 12 37 15
rect 39 20 47 25
rect 105 25 110 26
rect 94 20 99 25
rect 39 12 49 20
rect 29 7 34 12
rect 41 11 49 12
rect 41 7 42 11
rect 46 9 49 11
rect 51 19 58 20
rect 51 15 53 19
rect 57 15 58 19
rect 51 14 58 15
rect 51 9 56 14
rect 46 7 47 9
rect 7 4 8 7
rect 2 3 8 4
rect 41 6 47 7
rect 64 8 72 20
rect 64 4 65 8
rect 69 7 72 8
rect 74 7 79 20
rect 81 18 89 20
rect 81 14 83 18
rect 87 14 89 18
rect 81 7 89 14
rect 91 19 99 20
rect 91 15 93 19
rect 97 15 99 19
rect 91 12 99 15
rect 101 17 110 25
rect 101 13 103 17
rect 107 15 110 17
rect 112 25 119 26
rect 112 21 114 25
rect 118 21 119 25
rect 112 20 119 21
rect 112 15 117 20
rect 107 13 108 15
rect 101 12 108 13
rect 91 7 96 12
rect 69 4 70 7
rect 64 3 70 4
<< pdiffusion >>
rect 4 59 9 66
rect 2 58 9 59
rect 2 54 3 58
rect 7 54 9 58
rect 2 53 9 54
rect 4 38 9 53
rect 11 50 19 66
rect 11 46 13 50
rect 17 46 19 50
rect 11 38 19 46
rect 21 50 29 66
rect 21 46 23 50
rect 27 46 29 50
rect 21 43 29 46
rect 21 39 23 43
rect 27 39 29 43
rect 21 38 29 39
rect 31 65 39 66
rect 31 61 33 65
rect 37 61 39 65
rect 31 52 39 61
rect 41 58 49 66
rect 41 54 43 58
rect 47 54 49 58
rect 41 52 49 54
rect 51 65 58 66
rect 51 61 53 65
rect 57 61 58 65
rect 51 58 58 61
rect 64 59 69 66
rect 51 54 53 58
rect 57 54 58 58
rect 51 52 58 54
rect 62 58 69 59
rect 62 54 63 58
rect 67 54 69 58
rect 62 53 69 54
rect 31 38 37 52
rect 64 38 69 53
rect 71 50 79 66
rect 71 46 73 50
rect 77 46 79 50
rect 71 38 79 46
rect 81 50 89 66
rect 81 46 83 50
rect 87 46 89 50
rect 81 43 89 46
rect 81 39 83 43
rect 87 39 89 43
rect 81 38 89 39
rect 91 65 98 66
rect 91 61 93 65
rect 97 61 98 65
rect 116 68 122 69
rect 116 64 117 68
rect 121 64 122 68
rect 116 63 122 64
rect 91 56 98 61
rect 91 42 100 56
rect 102 52 107 56
rect 118 52 122 63
rect 102 47 110 52
rect 102 43 104 47
rect 108 43 110 47
rect 102 42 110 43
rect 91 38 98 42
rect 105 38 110 42
rect 112 38 122 52
<< metal1 >>
rect -2 68 130 72
rect -2 65 105 68
rect -2 64 33 65
rect 32 61 33 64
rect 37 64 53 65
rect 37 61 38 64
rect 52 61 53 64
rect 57 64 93 65
rect 57 61 58 64
rect 92 61 93 64
rect 97 64 105 65
rect 109 64 117 68
rect 121 64 130 68
rect 97 61 98 64
rect 52 58 58 61
rect 110 59 111 60
rect 2 54 3 58
rect 7 54 43 58
rect 47 54 48 58
rect 52 54 53 58
rect 57 54 58 58
rect 62 54 63 58
rect 67 54 94 58
rect 2 46 13 50
rect 17 46 18 50
rect 22 46 23 50
rect 27 46 28 50
rect 2 18 6 46
rect 22 43 28 46
rect 10 39 23 43
rect 27 39 28 43
rect 10 34 14 39
rect 32 34 36 54
rect 83 50 87 51
rect 41 48 54 50
rect 41 44 46 48
rect 19 30 20 34
rect 24 30 45 34
rect 10 26 14 30
rect 10 22 35 26
rect 31 19 35 22
rect 2 14 21 18
rect 25 14 26 18
rect 41 19 45 30
rect 50 28 54 48
rect 62 46 73 50
rect 77 46 78 50
rect 62 34 66 46
rect 83 43 87 46
rect 59 30 60 34
rect 64 30 66 34
rect 50 23 54 24
rect 41 15 53 19
rect 57 15 58 19
rect 62 18 66 30
rect 70 39 83 42
rect 70 38 87 39
rect 90 42 94 54
rect 106 56 111 59
rect 115 59 116 60
rect 115 56 118 59
rect 106 53 118 56
rect 104 47 108 48
rect 114 45 118 53
rect 104 42 108 43
rect 90 38 118 42
rect 70 34 74 38
rect 90 34 94 38
rect 79 30 80 34
rect 84 30 94 34
rect 98 33 111 35
rect 70 26 74 30
rect 102 29 111 33
rect 70 22 97 26
rect 105 22 111 29
rect 114 25 118 38
rect 93 19 97 22
rect 114 20 118 21
rect 31 14 35 15
rect 62 14 83 18
rect 87 14 88 18
rect 93 14 97 15
rect 103 17 107 18
rect 41 8 42 11
rect -2 4 3 8
rect 7 7 42 8
rect 46 8 47 11
rect 103 8 107 13
rect 46 7 65 8
rect 7 4 65 7
rect 69 4 116 8
rect 120 4 130 8
rect -2 0 130 4
<< ntransistor >>
rect 10 7 12 20
rect 17 7 19 20
rect 27 7 29 20
rect 37 12 39 25
rect 49 9 51 20
rect 72 7 74 20
rect 79 7 81 20
rect 89 7 91 20
rect 99 12 101 25
rect 110 15 112 26
<< ptransistor >>
rect 9 38 11 66
rect 19 38 21 66
rect 29 38 31 66
rect 39 52 41 66
rect 49 52 51 66
rect 69 38 71 66
rect 79 38 81 66
rect 89 38 91 66
rect 100 42 102 56
rect 110 38 112 52
<< polycontact >>
rect 46 44 50 48
rect 111 56 115 60
rect 10 30 14 34
rect 20 30 24 34
rect 60 30 64 34
rect 70 30 74 34
rect 80 30 84 34
rect 98 29 102 33
rect 50 24 54 28
<< ndcontact >>
rect 3 4 7 8
rect 21 14 25 18
rect 31 15 35 19
rect 42 7 46 11
rect 53 15 57 19
rect 65 4 69 8
rect 83 14 87 18
rect 93 15 97 19
rect 103 13 107 17
rect 114 21 118 25
<< pdcontact >>
rect 3 54 7 58
rect 13 46 17 50
rect 23 46 27 50
rect 23 39 27 43
rect 33 61 37 65
rect 43 54 47 58
rect 53 61 57 65
rect 53 54 57 58
rect 63 54 67 58
rect 73 46 77 50
rect 83 46 87 50
rect 83 39 87 43
rect 93 61 97 65
rect 117 64 121 68
rect 104 43 108 47
<< psubstratepcontact >>
rect 116 4 120 8
<< nsubstratencontact >>
rect 105 64 109 68
<< psubstratepdiff >>
rect 115 8 121 9
rect 115 4 116 8
rect 120 4 121 8
rect 115 3 121 4
<< nsubstratendiff >>
rect 102 68 112 69
rect 102 64 105 68
rect 109 64 112 68
rect 102 63 112 64
<< labels >>
rlabel polycontact 22 32 22 32 6 cn
rlabel ntransistor 73 18 73 18 6 an
rlabel polycontact 82 32 82 32 6 bn
rlabel metal1 12 16 12 16 6 z
rlabel metal1 20 16 20 16 6 z
rlabel metal1 4 32 4 32 6 z
rlabel metal1 12 48 12 48 6 z
rlabel metal1 44 48 44 48 6 c
rlabel metal1 25 56 25 56 6 cn
rlabel metal1 34 44 34 44 6 cn
rlabel metal1 64 4 64 4 6 vss
rlabel metal1 49 17 49 17 6 cn
rlabel polycontact 72 32 72 32 6 an
rlabel metal1 52 36 52 36 6 c
rlabel metal1 64 68 64 68 6 vdd
rlabel metal1 95 20 95 20 6 an
rlabel polycontact 100 32 100 32 6 a
rlabel metal1 86 32 86 32 6 bn
rlabel metal1 85 44 85 44 6 an
rlabel metal1 78 56 78 56 6 bn
rlabel metal1 108 28 108 28 6 a
rlabel metal1 116 31 116 31 6 bn
rlabel metal1 106 43 106 43 6 bn
rlabel metal1 116 52 116 52 6 b
rlabel metal1 108 56 108 56 6 b
<< end >>
