magic
tech scmos
timestamp 1179387016
<< checkpaint >>
rect -22 -22 62 94
<< ab >>
rect 0 0 40 72
<< pwell >>
rect -4 -4 44 32
<< nwell >>
rect -4 32 44 76
<< polysilicon >>
rect 12 66 14 70
rect 22 66 24 70
rect 29 66 31 70
rect 12 46 14 52
rect 9 45 15 46
rect 9 41 10 45
rect 14 41 15 45
rect 9 40 15 41
rect 9 18 11 40
rect 22 36 24 39
rect 17 35 24 36
rect 17 31 18 35
rect 22 31 24 35
rect 17 30 24 31
rect 29 35 31 39
rect 29 34 38 35
rect 29 30 33 34
rect 37 30 38 34
rect 19 18 21 30
rect 29 29 38 30
rect 29 18 31 29
rect 9 2 11 6
rect 19 2 21 6
rect 29 2 31 6
<< ndiffusion >>
rect 2 17 9 18
rect 2 13 3 17
rect 7 13 9 17
rect 2 12 9 13
rect 4 6 9 12
rect 11 17 19 18
rect 11 13 13 17
rect 17 13 19 17
rect 11 6 19 13
rect 21 11 29 18
rect 21 7 23 11
rect 27 7 29 11
rect 21 6 29 7
rect 31 17 38 18
rect 31 13 33 17
rect 37 13 38 17
rect 31 12 38 13
rect 31 6 36 12
<< pdiffusion >>
rect 4 65 12 66
rect 4 61 6 65
rect 10 61 12 65
rect 4 52 12 61
rect 14 58 22 66
rect 14 54 16 58
rect 20 54 22 58
rect 14 52 22 54
rect 17 39 22 52
rect 24 39 29 66
rect 31 65 38 66
rect 31 61 33 65
rect 37 61 38 65
rect 31 58 38 61
rect 31 54 33 58
rect 37 54 38 58
rect 31 39 38 54
<< metal1 >>
rect -2 65 42 72
rect -2 64 6 65
rect 5 61 6 64
rect 10 64 33 65
rect 10 61 11 64
rect 32 61 33 64
rect 37 64 42 65
rect 37 61 38 64
rect 32 58 38 61
rect 2 54 16 58
rect 20 54 23 58
rect 32 54 33 58
rect 37 54 38 58
rect 2 18 6 54
rect 10 45 14 46
rect 25 43 31 50
rect 10 26 14 41
rect 18 38 31 43
rect 18 35 22 38
rect 18 30 22 31
rect 25 30 33 34
rect 37 30 38 34
rect 10 22 23 26
rect 34 21 38 30
rect 2 17 8 18
rect 2 13 3 17
rect 7 13 8 17
rect 12 17 38 18
rect 12 13 13 17
rect 17 14 33 17
rect 17 13 18 14
rect 32 13 33 14
rect 37 13 38 17
rect 22 8 23 11
rect -2 7 23 8
rect 27 8 28 11
rect 27 7 42 8
rect -2 0 42 7
<< ntransistor >>
rect 9 6 11 18
rect 19 6 21 18
rect 29 6 31 18
<< ptransistor >>
rect 12 52 14 66
rect 22 39 24 66
rect 29 39 31 66
<< polycontact >>
rect 10 41 14 45
rect 18 31 22 35
rect 33 30 37 34
<< ndcontact >>
rect 3 13 7 17
rect 13 13 17 17
rect 23 7 27 11
rect 33 13 37 17
<< pdcontact >>
rect 6 61 10 65
rect 16 54 20 58
rect 33 61 37 65
rect 33 54 37 58
<< labels >>
rlabel metal1 4 32 4 32 6 z
rlabel metal1 12 36 12 36 6 b
rlabel metal1 12 56 12 56 6 z
rlabel metal1 20 4 20 4 6 vss
rlabel metal1 20 24 20 24 6 b
rlabel metal1 28 32 28 32 6 a1
rlabel metal1 20 40 20 40 6 a2
rlabel metal1 28 44 28 44 6 a2
rlabel metal1 20 56 20 56 6 z
rlabel metal1 20 68 20 68 6 vdd
rlabel ndcontact 35 15 35 15 6 n1
rlabel metal1 25 16 25 16 6 n1
rlabel metal1 36 24 36 24 6 a1
<< end >>
