magic
tech scmos
timestamp 1182081828
<< checkpaint >>
rect -25 -26 121 114
<< ab >>
rect 0 0 96 88
<< pwell >>
rect -7 -8 103 40
<< nwell >>
rect -7 40 103 96
<< polysilicon >>
rect 5 85 14 86
rect 5 81 6 85
rect 10 81 14 85
rect 5 80 14 81
rect 18 85 27 86
rect 18 81 22 85
rect 26 81 27 85
rect 18 80 27 81
rect 37 80 46 86
rect 50 80 59 86
rect 69 85 78 86
rect 69 81 70 85
rect 74 81 78 85
rect 69 80 78 81
rect 82 80 91 86
rect 9 77 11 80
rect 21 77 23 80
rect 41 77 43 80
rect 53 77 55 80
rect 73 77 75 80
rect 85 77 87 80
rect 9 48 11 51
rect 21 48 23 51
rect 41 48 43 51
rect 53 48 55 51
rect 73 48 75 51
rect 85 48 87 51
rect 2 42 11 48
rect 15 47 30 48
rect 15 43 22 47
rect 26 43 30 47
rect 15 42 30 43
rect 34 47 43 48
rect 34 43 38 47
rect 42 43 43 47
rect 34 42 43 43
rect 47 47 62 48
rect 47 43 54 47
rect 58 43 62 47
rect 47 42 62 43
rect 66 42 75 48
rect 79 47 94 48
rect 79 43 86 47
rect 90 43 94 47
rect 79 42 94 43
rect 2 32 17 38
rect 21 37 30 38
rect 21 33 22 37
rect 26 33 30 37
rect 21 32 30 33
rect 34 37 49 38
rect 34 33 38 37
rect 42 33 49 37
rect 34 32 49 33
rect 53 37 62 38
rect 53 33 54 37
rect 58 33 62 37
rect 53 32 62 33
rect 66 32 81 38
rect 85 37 94 38
rect 85 33 86 37
rect 90 33 94 37
rect 85 32 94 33
rect 9 29 11 32
rect 21 29 23 32
rect 41 29 43 32
rect 53 29 55 32
rect 73 29 75 32
rect 85 29 87 32
rect 9 8 11 11
rect 21 8 23 11
rect 41 8 43 11
rect 53 8 55 11
rect 73 8 75 11
rect 85 8 87 11
rect 5 7 14 8
rect 5 3 6 7
rect 10 3 14 7
rect 5 2 14 3
rect 18 2 27 8
rect 37 2 46 8
rect 50 7 59 8
rect 69 7 78 8
rect 50 3 51 7
rect 55 3 59 7
rect 50 2 59 3
rect 69 3 70 7
rect 74 3 78 7
rect 69 2 78 3
rect 82 2 91 8
<< ndiffusion >>
rect 2 11 9 29
rect 11 24 21 29
rect 11 20 14 24
rect 18 20 21 24
rect 11 17 21 20
rect 11 13 14 17
rect 18 13 21 17
rect 11 11 21 13
rect 23 26 30 29
rect 23 22 25 26
rect 29 22 30 26
rect 23 18 30 22
rect 23 14 25 18
rect 29 14 30 18
rect 23 11 30 14
rect 34 26 41 29
rect 34 22 35 26
rect 39 22 41 26
rect 34 18 41 22
rect 34 14 35 18
rect 39 14 41 18
rect 34 11 41 14
rect 43 26 53 29
rect 43 22 46 26
rect 50 22 53 26
rect 43 18 53 22
rect 43 14 46 18
rect 50 14 53 18
rect 43 11 53 14
rect 55 25 62 29
rect 55 21 57 25
rect 61 21 62 25
rect 55 18 62 21
rect 55 14 57 18
rect 61 14 62 18
rect 55 11 62 14
rect 66 11 73 29
rect 75 18 85 29
rect 75 14 78 18
rect 82 14 85 18
rect 75 11 85 14
rect 87 25 94 29
rect 87 21 89 25
rect 93 21 94 25
rect 87 18 94 21
rect 87 14 89 18
rect 93 14 94 18
rect 87 11 94 14
<< pdiffusion >>
rect 2 51 9 77
rect 11 75 21 77
rect 11 71 14 75
rect 18 71 21 75
rect 11 68 21 71
rect 11 64 14 68
rect 18 64 21 68
rect 11 51 21 64
rect 23 63 30 77
rect 23 59 25 63
rect 29 59 30 63
rect 23 56 30 59
rect 23 52 25 56
rect 29 52 30 56
rect 23 51 30 52
rect 34 71 41 77
rect 34 67 35 71
rect 39 67 41 71
rect 34 51 41 67
rect 43 51 53 77
rect 55 56 62 77
rect 55 52 57 56
rect 61 52 62 56
rect 55 51 62 52
rect 66 56 73 77
rect 66 52 67 56
rect 71 52 73 56
rect 66 51 73 52
rect 75 63 85 77
rect 75 59 78 63
rect 82 59 85 63
rect 75 56 85 59
rect 75 52 78 56
rect 82 52 85 56
rect 75 51 85 52
rect 87 74 94 77
rect 87 70 89 74
rect 93 70 94 74
rect 87 67 94 70
rect 87 63 89 67
rect 93 63 94 67
rect 87 51 94 63
<< metal1 >>
rect -2 86 2 90
rect 30 86 34 90
rect 2 82 6 85
rect -2 81 6 82
rect 10 81 18 85
rect 14 75 18 81
rect 21 81 22 85
rect 26 81 27 85
rect 30 81 34 82
rect 62 86 66 90
rect 94 86 98 90
rect 62 81 66 82
rect 69 81 70 85
rect 74 81 75 85
rect 21 78 27 81
rect 69 78 75 81
rect 21 74 75 78
rect 89 82 94 85
rect 89 81 98 82
rect 89 74 93 81
rect 14 68 35 71
rect 18 67 35 68
rect 39 67 40 71
rect 89 67 93 70
rect 14 63 18 64
rect 25 63 29 64
rect 14 48 18 59
rect 25 56 29 59
rect 38 63 82 64
rect 38 60 78 63
rect 29 52 34 55
rect 25 51 34 52
rect 14 47 26 48
rect 14 44 22 47
rect 22 37 26 43
rect 22 29 26 33
rect 30 26 34 51
rect 38 47 42 60
rect 89 62 93 63
rect 78 56 82 59
rect 38 37 42 43
rect 38 32 42 33
rect 46 52 57 56
rect 61 52 67 56
rect 71 52 72 56
rect 46 26 50 52
rect 54 47 58 48
rect 54 37 58 43
rect 54 32 58 33
rect 78 26 82 52
rect 86 47 90 51
rect 86 37 90 43
rect 86 29 90 33
rect 14 24 18 25
rect 24 22 25 26
rect 29 22 35 26
rect 39 22 40 26
rect 14 17 18 20
rect 30 18 34 22
rect 46 18 50 22
rect 24 14 25 18
rect 29 14 35 18
rect 39 14 42 18
rect 14 7 18 13
rect 38 7 42 14
rect 46 13 50 14
rect 57 25 93 26
rect 61 22 89 25
rect 57 18 61 21
rect 57 13 61 14
rect 78 18 82 19
rect 78 7 82 14
rect 89 18 93 21
rect 89 13 93 14
rect -2 6 6 7
rect 2 3 6 6
rect 10 6 34 7
rect 10 3 30 6
rect -2 -2 2 2
rect 38 3 51 7
rect 55 3 56 7
rect 62 6 70 7
rect 30 -2 34 2
rect 66 3 70 6
rect 74 6 98 7
rect 74 3 94 6
rect 62 -2 66 2
rect 94 -2 98 2
<< metal2 >>
rect -2 86 98 90
rect 2 82 30 86
rect 34 82 62 86
rect 66 82 94 86
rect -2 80 98 82
rect -2 6 98 8
rect 2 2 30 6
rect 34 2 62 6
rect 66 2 94 6
rect -2 -2 98 2
<< ntransistor >>
rect 9 11 11 29
rect 21 11 23 29
rect 41 11 43 29
rect 53 11 55 29
rect 73 11 75 29
rect 85 11 87 29
<< ptransistor >>
rect 9 51 11 77
rect 21 51 23 77
rect 41 51 43 77
rect 53 51 55 77
rect 73 51 75 77
rect 85 51 87 77
<< polycontact >>
rect 6 81 10 85
rect 22 81 26 85
rect 70 81 74 85
rect 22 43 26 47
rect 38 43 42 47
rect 54 43 58 47
rect 86 43 90 47
rect 22 33 26 37
rect 38 33 42 37
rect 54 33 58 37
rect 86 33 90 37
rect 6 3 10 7
rect 51 3 55 7
rect 70 3 74 7
<< ndcontact >>
rect 14 20 18 24
rect 14 13 18 17
rect 25 22 29 26
rect 25 14 29 18
rect 35 22 39 26
rect 35 14 39 18
rect 46 22 50 26
rect 46 14 50 18
rect 57 21 61 25
rect 57 14 61 18
rect 78 14 82 18
rect 89 21 93 25
rect 89 14 93 18
<< pdcontact >>
rect 14 71 18 75
rect 14 64 18 68
rect 25 59 29 63
rect 25 52 29 56
rect 35 67 39 71
rect 57 52 61 56
rect 67 52 71 56
rect 78 59 82 63
rect 78 52 82 56
rect 89 70 93 74
rect 89 63 93 67
<< m2contact >>
rect -2 82 2 86
rect 30 82 34 86
rect 62 82 66 86
rect 94 82 98 86
rect -2 2 2 6
rect 30 2 34 6
rect 62 2 66 6
rect 94 2 98 6
<< psubstratepcontact >>
rect -2 2 2 6
rect 30 2 34 6
rect 62 2 66 6
rect 94 2 98 6
<< nsubstratencontact >>
rect -2 82 2 86
rect 30 82 34 86
rect 62 82 66 86
rect 94 82 98 86
<< psubstratepdiff >>
rect -3 6 3 7
rect -3 2 -2 6
rect 2 2 3 6
rect 29 6 35 7
rect 29 2 30 6
rect 34 2 35 6
rect 61 6 67 7
rect 61 2 62 6
rect 66 2 67 6
rect 93 6 99 7
rect 93 2 94 6
rect 98 2 99 6
rect -3 0 3 2
rect 29 0 35 2
rect 61 0 67 2
rect 93 0 99 2
<< nsubstratendiff >>
rect -3 86 3 88
rect 29 86 35 88
rect 61 86 67 88
rect 93 86 99 88
rect -3 82 -2 86
rect 2 82 3 86
rect -3 81 3 82
rect 29 82 30 86
rect 34 82 35 86
rect 29 81 35 82
rect 61 82 62 86
rect 66 82 67 86
rect 61 81 67 82
rect 93 82 94 86
rect 98 82 99 86
rect 93 81 99 82
<< labels >>
rlabel polycontact 24 36 24 36 6 b
rlabel metal1 16 52 16 52 6 b
rlabel metal1 48 32 48 32 6 z
rlabel metal1 88 40 88 40 6 a
rlabel metal2 48 4 48 4 6 vss
rlabel metal2 48 84 48 84 6 vdd
<< end >>
