magic
tech scmos
timestamp 1179385318
<< checkpaint >>
rect -22 -25 166 105
<< ab >>
rect 0 0 144 80
<< pwell >>
rect -4 -7 148 36
<< nwell >>
rect -4 36 148 87
<< polysilicon >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 39 70 41 74
rect 49 70 51 74
rect 59 70 61 74
rect 69 70 71 74
rect 79 70 81 74
rect 89 70 91 74
rect 99 70 101 74
rect 109 70 111 74
rect 119 70 121 74
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 39 39 41 42
rect 49 39 51 42
rect 59 39 61 42
rect 69 39 71 42
rect 79 39 81 42
rect 89 39 91 42
rect 99 39 101 42
rect 109 39 111 42
rect 9 38 15 39
rect 9 34 10 38
rect 14 34 15 38
rect 19 38 34 39
rect 19 37 26 38
rect 9 33 15 34
rect 25 34 26 37
rect 30 34 34 38
rect 25 33 34 34
rect 32 30 34 33
rect 39 38 51 39
rect 39 34 42 38
rect 46 34 51 38
rect 39 33 51 34
rect 39 30 41 33
rect 49 30 51 33
rect 56 38 63 39
rect 56 34 58 38
rect 62 34 63 38
rect 56 33 63 34
rect 68 38 74 39
rect 68 34 69 38
rect 73 34 74 38
rect 68 33 74 34
rect 56 30 58 33
rect 72 30 74 33
rect 79 38 91 39
rect 79 34 82 38
rect 86 34 91 38
rect 79 33 91 34
rect 79 30 81 33
rect 89 30 91 33
rect 96 38 111 39
rect 96 34 98 38
rect 102 34 106 38
rect 110 34 111 38
rect 96 33 111 34
rect 119 39 121 42
rect 119 38 127 39
rect 119 34 122 38
rect 126 34 127 38
rect 119 33 127 34
rect 96 30 98 33
rect 32 6 34 11
rect 39 6 41 11
rect 49 6 51 11
rect 56 6 58 11
rect 72 6 74 11
rect 79 6 81 11
rect 89 6 91 11
rect 96 6 98 11
<< ndiffusion >>
rect 23 12 32 30
rect 23 8 25 12
rect 29 11 32 12
rect 34 11 39 30
rect 41 22 49 30
rect 41 18 43 22
rect 47 18 49 22
rect 41 11 49 18
rect 51 11 56 30
rect 58 14 72 30
rect 58 11 63 14
rect 29 8 30 11
rect 23 7 30 8
rect 60 10 63 11
rect 67 11 72 14
rect 74 11 79 30
rect 81 22 89 30
rect 81 18 83 22
rect 87 18 89 22
rect 81 11 89 18
rect 91 11 96 30
rect 98 23 106 30
rect 98 19 100 23
rect 104 19 106 23
rect 98 16 106 19
rect 98 12 100 16
rect 104 12 106 16
rect 98 11 106 12
rect 67 10 70 11
rect 60 9 70 10
<< pdiffusion >>
rect 4 64 9 70
rect 2 63 9 64
rect 2 59 3 63
rect 7 59 9 63
rect 2 56 9 59
rect 2 52 3 56
rect 7 52 9 56
rect 2 51 9 52
rect 4 42 9 51
rect 11 54 19 70
rect 11 50 13 54
rect 17 50 19 54
rect 11 47 19 50
rect 11 43 13 47
rect 17 43 19 47
rect 11 42 19 43
rect 21 63 29 70
rect 21 59 23 63
rect 27 59 29 63
rect 21 42 29 59
rect 31 54 39 70
rect 31 50 33 54
rect 37 50 39 54
rect 31 42 39 50
rect 41 63 49 70
rect 41 59 43 63
rect 47 59 49 63
rect 41 42 49 59
rect 51 54 59 70
rect 51 50 53 54
rect 57 50 59 54
rect 51 42 59 50
rect 61 62 69 70
rect 61 58 63 62
rect 67 58 69 62
rect 61 55 69 58
rect 61 51 63 55
rect 67 51 69 55
rect 61 42 69 51
rect 71 69 79 70
rect 71 65 73 69
rect 77 65 79 69
rect 71 62 79 65
rect 71 58 73 62
rect 77 58 79 62
rect 71 42 79 58
rect 81 61 89 70
rect 81 57 83 61
rect 87 57 89 61
rect 81 54 89 57
rect 81 50 83 54
rect 87 50 89 54
rect 81 42 89 50
rect 91 69 99 70
rect 91 65 93 69
rect 97 65 99 69
rect 91 62 99 65
rect 91 58 93 62
rect 97 58 99 62
rect 91 42 99 58
rect 101 61 109 70
rect 101 57 103 61
rect 107 57 109 61
rect 101 54 109 57
rect 101 50 103 54
rect 107 50 109 54
rect 101 42 109 50
rect 111 69 119 70
rect 111 65 113 69
rect 117 65 119 69
rect 111 62 119 65
rect 111 58 113 62
rect 117 58 119 62
rect 111 42 119 58
rect 121 55 126 70
rect 121 54 128 55
rect 121 50 123 54
rect 127 50 128 54
rect 121 47 128 50
rect 121 43 123 47
rect 127 43 128 47
rect 121 42 128 43
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect 118 78 122 82
rect 126 78 130 82
rect 134 78 138 82
rect 142 78 146 82
rect -2 69 146 78
rect -2 68 73 69
rect 72 65 73 68
rect 77 68 93 69
rect 77 65 78 68
rect 2 59 3 63
rect 7 59 23 63
rect 27 59 43 63
rect 47 62 67 63
rect 47 59 63 62
rect 2 56 7 59
rect 2 52 3 56
rect 72 62 78 65
rect 92 65 93 68
rect 97 68 113 69
rect 97 65 98 68
rect 92 62 98 65
rect 112 65 113 68
rect 117 68 146 69
rect 117 65 118 68
rect 112 62 118 65
rect 72 58 73 62
rect 77 58 78 62
rect 83 61 87 62
rect 63 55 67 58
rect 2 51 7 52
rect 12 50 13 54
rect 17 50 33 54
rect 37 50 53 54
rect 57 50 58 54
rect 92 58 93 62
rect 97 58 98 62
rect 103 61 107 62
rect 83 54 87 57
rect 112 58 113 62
rect 117 58 118 62
rect 103 54 107 57
rect 67 51 83 54
rect 63 50 83 51
rect 87 50 103 54
rect 107 50 123 54
rect 127 50 128 54
rect 12 47 18 50
rect 2 43 13 47
rect 17 43 18 47
rect 122 47 128 50
rect 2 22 6 43
rect 25 42 63 46
rect 10 38 14 39
rect 25 38 31 42
rect 57 38 63 42
rect 25 34 26 38
rect 30 34 31 38
rect 41 34 42 38
rect 46 34 47 38
rect 57 34 58 38
rect 62 34 63 38
rect 69 42 103 46
rect 122 43 123 47
rect 127 43 128 47
rect 69 38 73 42
rect 97 38 103 42
rect 122 38 126 39
rect 10 30 14 34
rect 41 30 47 34
rect 69 30 73 34
rect 10 26 47 30
rect 65 26 73 30
rect 81 34 82 38
rect 86 34 87 38
rect 97 34 98 38
rect 102 34 106 38
rect 110 34 111 38
rect 81 30 87 34
rect 122 30 126 34
rect 81 26 126 30
rect 2 18 43 22
rect 47 18 83 22
rect 87 18 88 22
rect 99 19 100 23
rect 104 19 105 23
rect 99 16 105 19
rect 122 17 126 26
rect 62 12 63 14
rect -2 8 25 12
rect 29 10 63 12
rect 67 12 68 14
rect 99 12 100 16
rect 104 12 105 16
rect 67 10 146 12
rect 29 8 146 10
rect -2 2 146 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 122 2
rect 126 -2 130 2
rect 134 -2 138 2
rect 142 -2 146 2
<< ntransistor >>
rect 32 11 34 30
rect 39 11 41 30
rect 49 11 51 30
rect 56 11 58 30
rect 72 11 74 30
rect 79 11 81 30
rect 89 11 91 30
rect 96 11 98 30
<< ptransistor >>
rect 9 42 11 70
rect 19 42 21 70
rect 29 42 31 70
rect 39 42 41 70
rect 49 42 51 70
rect 59 42 61 70
rect 69 42 71 70
rect 79 42 81 70
rect 89 42 91 70
rect 99 42 101 70
rect 109 42 111 70
rect 119 42 121 70
<< polycontact >>
rect 10 34 14 38
rect 26 34 30 38
rect 42 34 46 38
rect 58 34 62 38
rect 69 34 73 38
rect 82 34 86 38
rect 98 34 102 38
rect 106 34 110 38
rect 122 34 126 38
<< ndcontact >>
rect 25 8 29 12
rect 43 18 47 22
rect 63 10 67 14
rect 83 18 87 22
rect 100 19 104 23
rect 100 12 104 16
<< pdcontact >>
rect 3 59 7 63
rect 3 52 7 56
rect 13 50 17 54
rect 13 43 17 47
rect 23 59 27 63
rect 33 50 37 54
rect 43 59 47 63
rect 53 50 57 54
rect 63 58 67 62
rect 63 51 67 55
rect 73 65 77 69
rect 73 58 77 62
rect 83 57 87 61
rect 83 50 87 54
rect 93 65 97 69
rect 93 58 97 62
rect 103 57 107 61
rect 103 50 107 54
rect 113 65 117 69
rect 113 58 117 62
rect 123 50 127 54
rect 123 43 127 47
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
rect 90 -2 94 2
rect 98 -2 102 2
rect 106 -2 110 2
rect 114 -2 118 2
rect 122 -2 126 2
rect 130 -2 134 2
rect 138 -2 142 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
rect 90 78 94 82
rect 98 78 102 82
rect 106 78 110 82
rect 114 78 118 82
rect 122 78 126 82
rect 130 78 134 82
rect 138 78 142 82
<< psubstratepdiff >>
rect 0 2 144 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 122 2
rect 126 -2 130 2
rect 134 -2 138 2
rect 142 -2 144 2
rect 0 -3 144 -2
<< nsubstratendiff >>
rect 0 82 144 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect 118 78 122 82
rect 126 78 130 82
rect 134 78 138 82
rect 142 78 144 82
rect 0 77 144 78
<< labels >>
rlabel metal1 12 20 12 20 6 z
rlabel polycontact 12 36 12 36 6 b2
rlabel metal1 4 36 4 36 6 z
rlabel metal1 4 57 4 57 6 n3
rlabel metal1 20 20 20 20 6 z
rlabel metal1 36 20 36 20 6 z
rlabel ndcontact 44 20 44 20 6 z
rlabel metal1 28 20 28 20 6 z
rlabel metal1 28 28 28 28 6 b2
rlabel metal1 36 28 36 28 6 b2
rlabel metal1 20 28 20 28 6 b2
rlabel metal1 44 32 44 32 6 b2
rlabel metal1 28 40 28 40 6 b1
rlabel metal1 44 44 44 44 6 b1
rlabel metal1 36 44 36 44 6 b1
rlabel metal1 20 52 20 52 6 z
rlabel metal1 28 52 28 52 6 z
rlabel metal1 44 52 44 52 6 z
rlabel pdcontact 36 52 36 52 6 z
rlabel metal1 68 20 68 20 6 z
rlabel metal1 60 20 60 20 6 z
rlabel metal1 52 20 52 20 6 z
rlabel metal1 68 28 68 28 6 a1
rlabel metal1 52 44 52 44 6 b1
rlabel metal1 60 40 60 40 6 b1
rlabel metal1 52 52 52 52 6 z
rlabel metal1 65 56 65 56 6 n3
rlabel metal1 34 61 34 61 6 n3
rlabel metal1 72 6 72 6 6 vss
rlabel metal1 76 20 76 20 6 z
rlabel ndcontact 84 20 84 20 6 z
rlabel metal1 92 28 92 28 6 a2
rlabel metal1 84 32 84 32 6 a2
rlabel metal1 84 44 84 44 6 a1
rlabel metal1 92 44 92 44 6 a1
rlabel metal1 76 44 76 44 6 a1
rlabel metal1 85 56 85 56 6 n3
rlabel metal1 72 74 72 74 6 vdd
rlabel metal1 108 28 108 28 6 a2
rlabel metal1 116 28 116 28 6 a2
rlabel metal1 100 28 100 28 6 a2
rlabel polycontact 108 36 108 36 6 a1
rlabel metal1 100 40 100 40 6 a1
rlabel metal1 105 56 105 56 6 n3
rlabel metal1 124 28 124 28 6 a2
rlabel metal1 125 48 125 48 6 n3
rlabel metal1 95 52 95 52 6 n3
<< end >>
