magic
tech scmos
timestamp 1179386970
<< checkpaint >>
rect -22 -25 78 105
<< ab >>
rect 0 0 56 80
<< pwell >>
rect -4 -7 60 36
<< nwell >>
rect -4 36 60 87
<< polysilicon >>
rect 38 70 40 74
rect 45 70 47 74
rect 10 61 12 65
rect 20 61 22 65
rect 10 38 12 46
rect 20 39 22 46
rect 38 40 40 43
rect 34 39 40 40
rect 19 38 25 39
rect 9 37 15 38
rect 9 33 10 37
rect 14 33 15 37
rect 9 32 15 33
rect 19 34 20 38
rect 24 34 25 38
rect 34 36 35 39
rect 19 33 25 34
rect 29 35 35 36
rect 39 35 40 39
rect 29 34 40 35
rect 45 38 47 43
rect 45 37 54 38
rect 12 29 14 32
rect 19 29 21 33
rect 29 29 31 34
rect 45 33 49 37
rect 53 33 54 37
rect 45 32 54 33
rect 45 29 47 32
rect 12 7 14 12
rect 19 7 21 12
rect 29 7 31 12
rect 45 7 47 12
<< ndiffusion >>
rect 7 22 12 29
rect 5 21 12 22
rect 5 17 6 21
rect 10 17 12 21
rect 5 16 12 17
rect 7 12 12 16
rect 14 12 19 29
rect 21 21 29 29
rect 21 17 23 21
rect 27 17 29 21
rect 21 12 29 17
rect 31 12 45 29
rect 47 22 52 29
rect 47 21 54 22
rect 47 17 49 21
rect 53 17 54 21
rect 47 16 54 17
rect 47 12 52 16
rect 33 8 36 12
rect 40 8 43 12
rect 33 7 43 8
<< pdiffusion >>
rect 24 69 38 70
rect 24 65 28 69
rect 32 65 38 69
rect 2 64 8 65
rect 2 60 3 64
rect 7 61 8 64
rect 24 61 38 65
rect 7 60 10 61
rect 2 46 10 60
rect 12 60 20 61
rect 12 56 14 60
rect 18 56 20 60
rect 12 46 20 56
rect 22 46 38 61
rect 24 43 38 46
rect 40 43 45 70
rect 47 62 52 70
rect 47 61 54 62
rect 47 57 49 61
rect 53 57 54 61
rect 47 54 54 57
rect 47 50 49 54
rect 53 50 54 54
rect 47 49 54 50
rect 47 43 52 49
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect -2 69 58 78
rect -2 68 28 69
rect 3 64 7 68
rect 27 65 28 68
rect 32 68 58 69
rect 32 65 33 68
rect 3 59 7 60
rect 14 61 54 62
rect 14 60 49 61
rect 18 58 49 60
rect 14 55 18 56
rect 2 50 18 55
rect 53 57 54 61
rect 49 54 54 57
rect 25 50 39 54
rect 2 17 6 50
rect 10 42 23 46
rect 33 42 39 50
rect 53 50 54 54
rect 49 49 54 50
rect 10 37 14 42
rect 35 39 39 42
rect 10 25 14 33
rect 18 34 20 38
rect 24 34 31 38
rect 35 34 39 35
rect 49 37 54 39
rect 18 25 22 34
rect 53 33 54 37
rect 49 30 54 33
rect 41 25 54 30
rect 10 17 11 21
rect 22 17 23 21
rect 27 17 49 21
rect 53 17 54 21
rect -2 8 36 12
rect 40 8 58 12
rect -2 2 58 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
<< ntransistor >>
rect 12 12 14 29
rect 19 12 21 29
rect 29 12 31 29
rect 45 12 47 29
<< ptransistor >>
rect 10 46 12 61
rect 20 46 22 61
rect 38 43 40 70
rect 45 43 47 70
<< polycontact >>
rect 10 33 14 37
rect 20 34 24 38
rect 35 35 39 39
rect 49 33 53 37
<< ndcontact >>
rect 6 17 10 21
rect 23 17 27 21
rect 49 17 53 21
rect 36 8 40 12
<< pdcontact >>
rect 28 65 32 69
rect 3 60 7 64
rect 14 56 18 60
rect 49 57 53 61
rect 49 50 53 54
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
<< psubstratepdiff >>
rect 0 2 56 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 56 2
rect 0 -3 56 -2
<< nsubstratendiff >>
rect 0 82 56 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 56 82
rect 0 77 56 78
<< labels >>
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 32 12 32 6 c
rlabel metal1 12 52 12 52 6 z
rlabel metal1 28 6 28 6 6 vss
rlabel metal1 20 28 20 28 6 b
rlabel metal1 20 44 20 44 6 c
rlabel metal1 28 36 28 36 6 b
rlabel metal1 28 52 28 52 6 a1
rlabel metal1 20 60 20 60 6 z
rlabel metal1 28 60 28 60 6 z
rlabel metal1 28 74 28 74 6 vdd
rlabel metal1 44 28 44 28 6 a2
rlabel metal1 36 48 36 48 6 a1
rlabel metal1 36 60 36 60 6 z
rlabel metal1 44 60 44 60 6 z
rlabel metal1 38 19 38 19 6 n1
rlabel metal1 52 32 52 32 6 a2
rlabel pdcontact 52 52 52 52 6 z
<< end >>
