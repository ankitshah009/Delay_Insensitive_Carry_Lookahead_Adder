magic
tech scmos
timestamp 1180600766
<< checkpaint >>
rect -22 -22 142 122
<< ab >>
rect 0 0 120 100
<< pwell >>
rect -4 -4 124 48
<< nwell >>
rect -4 48 124 104
<< polysilicon >>
rect 23 94 25 98
rect 35 94 37 98
rect 47 94 49 98
rect 59 94 61 98
rect 11 76 13 80
rect 11 53 13 56
rect 23 53 25 56
rect 11 52 25 53
rect 11 51 18 52
rect 17 48 18 51
rect 22 51 25 52
rect 35 53 37 56
rect 95 94 97 98
rect 107 94 109 98
rect 71 76 73 80
rect 35 52 43 53
rect 35 51 38 52
rect 22 48 23 51
rect 17 47 23 48
rect 37 48 38 51
rect 42 48 43 52
rect 37 47 43 48
rect 3 42 9 43
rect 3 38 4 42
rect 8 41 9 42
rect 47 41 49 55
rect 59 53 61 56
rect 71 53 73 56
rect 59 52 73 53
rect 59 51 68 52
rect 67 48 68 51
rect 72 48 73 52
rect 67 47 73 48
rect 95 43 97 55
rect 107 43 109 55
rect 8 39 49 41
rect 8 38 9 39
rect 3 37 9 38
rect 17 32 23 33
rect 17 29 18 32
rect 11 28 18 29
rect 22 29 23 32
rect 37 32 43 33
rect 37 29 38 32
rect 22 28 25 29
rect 11 27 25 28
rect 11 24 13 27
rect 23 24 25 27
rect 35 28 38 29
rect 42 28 43 32
rect 35 27 43 28
rect 35 24 37 27
rect 47 25 49 39
rect 57 42 63 43
rect 57 38 58 42
rect 62 41 63 42
rect 77 42 83 43
rect 77 41 78 42
rect 62 39 78 41
rect 62 38 63 39
rect 57 37 63 38
rect 77 38 78 39
rect 82 38 83 42
rect 77 37 83 38
rect 87 42 109 43
rect 87 38 88 42
rect 92 38 109 42
rect 87 37 109 38
rect 59 25 61 37
rect 67 32 73 33
rect 67 28 68 32
rect 72 28 73 32
rect 67 27 73 28
rect 11 10 13 14
rect 71 24 73 27
rect 95 25 97 37
rect 107 25 109 37
rect 71 10 73 14
rect 23 2 25 6
rect 35 2 37 6
rect 47 2 49 6
rect 59 2 61 6
rect 95 2 97 6
rect 107 2 109 6
<< ndiffusion >>
rect 42 24 47 25
rect 3 22 11 24
rect 3 18 4 22
rect 8 18 11 22
rect 3 14 11 18
rect 13 14 23 24
rect 15 12 23 14
rect 15 8 16 12
rect 20 8 23 12
rect 15 6 23 8
rect 25 6 35 24
rect 37 22 47 24
rect 37 18 40 22
rect 44 18 47 22
rect 37 6 47 18
rect 49 6 59 25
rect 61 24 66 25
rect 75 32 83 33
rect 75 28 78 32
rect 82 28 83 32
rect 75 27 83 28
rect 75 24 81 27
rect 61 14 71 24
rect 73 14 81 24
rect 90 21 95 25
rect 61 12 69 14
rect 61 8 64 12
rect 68 8 69 12
rect 87 12 95 21
rect 61 6 69 8
rect 87 8 88 12
rect 92 8 95 12
rect 87 6 95 8
rect 97 22 107 25
rect 97 18 100 22
rect 104 18 107 22
rect 97 6 107 18
rect 109 22 117 25
rect 109 18 112 22
rect 116 18 117 22
rect 109 12 117 18
rect 109 8 112 12
rect 116 8 117 12
rect 109 6 117 8
<< pdiffusion >>
rect 15 92 23 94
rect 15 88 16 92
rect 20 88 23 92
rect 15 76 23 88
rect 3 62 11 76
rect 3 58 4 62
rect 8 58 11 62
rect 3 56 11 58
rect 13 56 23 76
rect 25 82 35 94
rect 25 78 28 82
rect 32 78 35 82
rect 25 56 35 78
rect 37 72 47 94
rect 37 68 40 72
rect 44 68 47 72
rect 37 56 47 68
rect 42 55 47 56
rect 49 82 59 94
rect 49 78 52 82
rect 56 78 59 82
rect 49 56 59 78
rect 61 92 69 94
rect 61 88 64 92
rect 68 88 69 92
rect 61 76 69 88
rect 87 92 95 94
rect 87 88 88 92
rect 92 88 95 92
rect 87 82 95 88
rect 87 78 88 82
rect 92 78 95 82
rect 61 56 71 76
rect 73 61 81 76
rect 87 72 95 78
rect 87 68 88 72
rect 92 68 95 72
rect 87 67 95 68
rect 73 60 83 61
rect 73 56 78 60
rect 82 56 83 60
rect 49 55 54 56
rect 77 55 83 56
rect 90 55 95 67
rect 97 82 107 94
rect 97 78 100 82
rect 104 78 107 82
rect 97 72 107 78
rect 97 68 100 72
rect 104 68 107 72
rect 97 62 107 68
rect 97 58 100 62
rect 104 58 107 62
rect 97 55 107 58
rect 109 92 117 94
rect 109 88 112 92
rect 116 88 117 92
rect 109 82 117 88
rect 109 78 112 82
rect 116 78 117 82
rect 109 72 117 78
rect 109 68 112 72
rect 116 68 117 72
rect 109 62 117 68
rect 109 58 112 62
rect 116 58 117 62
rect 109 55 117 58
<< metal1 >>
rect -2 96 122 100
rect -2 92 4 96
rect 8 92 76 96
rect 80 92 122 96
rect -2 88 16 92
rect 20 88 64 92
rect 68 88 88 92
rect 92 88 112 92
rect 116 88 122 92
rect 4 62 8 63
rect 4 42 8 58
rect 4 22 8 38
rect 4 17 8 18
rect 18 52 22 83
rect 27 78 28 82
rect 32 78 52 82
rect 56 78 57 82
rect 18 32 22 48
rect 18 17 22 28
rect 28 68 40 72
rect 44 68 45 72
rect 28 22 32 68
rect 68 52 72 83
rect 88 82 92 88
rect 88 72 92 78
rect 88 67 92 68
rect 98 82 102 83
rect 112 82 116 88
rect 98 78 100 82
rect 104 78 105 82
rect 98 72 102 78
rect 112 72 116 78
rect 98 68 100 72
rect 104 68 105 72
rect 98 62 102 68
rect 112 62 116 68
rect 37 48 38 52
rect 42 48 52 52
rect 48 42 52 48
rect 48 38 58 42
rect 62 38 63 42
rect 68 32 72 48
rect 37 28 38 32
rect 42 28 68 32
rect 68 27 72 28
rect 78 60 82 61
rect 78 42 82 56
rect 98 58 100 62
rect 104 58 105 62
rect 78 32 82 38
rect 78 27 82 28
rect 88 42 92 43
rect 88 22 92 38
rect 28 18 40 22
rect 44 18 92 22
rect 98 22 102 58
rect 112 57 116 58
rect 112 22 116 23
rect 98 18 100 22
rect 104 18 105 22
rect 98 17 102 18
rect 112 12 116 18
rect -2 8 16 12
rect 20 8 64 12
rect 68 8 88 12
rect 92 8 112 12
rect 116 8 122 12
rect -2 0 122 8
<< ntransistor >>
rect 11 14 13 24
rect 23 6 25 24
rect 35 6 37 24
rect 47 6 49 25
rect 59 6 61 25
rect 71 14 73 24
rect 95 6 97 25
rect 107 6 109 25
<< ptransistor >>
rect 11 56 13 76
rect 23 56 25 94
rect 35 56 37 94
rect 47 55 49 94
rect 59 56 61 94
rect 71 56 73 76
rect 95 55 97 94
rect 107 55 109 94
<< polycontact >>
rect 18 48 22 52
rect 38 48 42 52
rect 4 38 8 42
rect 68 48 72 52
rect 18 28 22 32
rect 38 28 42 32
rect 58 38 62 42
rect 78 38 82 42
rect 88 38 92 42
rect 68 28 72 32
<< ndcontact >>
rect 4 18 8 22
rect 16 8 20 12
rect 40 18 44 22
rect 78 28 82 32
rect 64 8 68 12
rect 88 8 92 12
rect 100 18 104 22
rect 112 18 116 22
rect 112 8 116 12
<< pdcontact >>
rect 16 88 20 92
rect 4 58 8 62
rect 28 78 32 82
rect 40 68 44 72
rect 52 78 56 82
rect 64 88 68 92
rect 88 88 92 92
rect 88 78 92 82
rect 88 68 92 72
rect 78 56 82 60
rect 100 78 104 82
rect 100 68 104 72
rect 100 58 104 62
rect 112 88 116 92
rect 112 78 116 82
rect 112 68 116 72
rect 112 58 116 62
<< nsubstratencontact >>
rect 4 92 8 96
rect 76 92 80 96
<< nsubstratendiff >>
rect 3 96 9 97
rect 3 92 4 96
rect 8 92 9 96
rect 75 96 81 97
rect 3 86 9 92
rect 75 92 76 96
rect 80 92 81 96
rect 75 86 81 92
<< labels >>
rlabel polycontact 40 30 40 30 6 i1
rlabel polycontact 20 50 20 50 6 i0
rlabel metal1 60 6 60 6 6 vss
rlabel metal1 50 30 50 30 6 i1
rlabel metal1 60 30 60 30 6 i1
rlabel metal1 60 94 60 94 6 vdd
rlabel metal1 70 55 70 55 6 i1
rlabel metal1 100 50 100 50 6 nq
<< end >>
