.subckt na2_x4 i0 i1 nq vdd vss
*   SPICE3 file   created from na2_x4.ext -      technology: scmos
m00 w1     i0     vdd    vdd p w=20u  l=2.3636u ad=100p     pd=30u      as=124p     ps=38.8571u
m01 vdd    i1     w1     vdd p w=20u  l=2.3636u ad=124p     pd=38.8571u as=100p     ps=30u
m02 nq     w2     vdd    vdd p w=40u  l=2.3636u ad=200p     pd=50u      as=248p     ps=77.7143u
m03 vdd    w2     nq     vdd p w=40u  l=2.3636u ad=248p     pd=77.7143u as=200p     ps=50u
m04 w2     w1     vdd    vdd p w=20u  l=2.3636u ad=160p     pd=56u      as=124p     ps=38.8571u
m05 w3     i0     w1     vss n w=20u  l=2.3636u ad=80p      pd=28u      as=160p     ps=56u
m06 vss    i1     w3     vss n w=20u  l=2.3636u ad=125.714p pd=40u      as=80p      ps=28u
m07 nq     w2     vss    vss n w=20u  l=2.3636u ad=100p     pd=30u      as=125.714p ps=40u
m08 vss    w2     nq     vss n w=20u  l=2.3636u ad=125.714p pd=40u      as=100p     ps=30u
m09 w2     w1     vss    vss n w=10u  l=2.3636u ad=80p      pd=36u      as=62.8571p ps=20u
C0  vdd    w2     0.026f
C1  vss    i1     0.019f
C2  w3     w1     0.016f
C3  nq     i1     0.095f
C4  w3     i0     0.004f
C5  w1     i0     0.142f
C6  nq     vdd    0.043f
C7  i1     vdd    0.015f
C8  w1     w2     0.199f
C9  i0     w2     0.028f
C10 vss    w1     0.232f
C11 nq     w1     0.408f
C12 vss    i0     0.015f
C13 w3     i1     0.012f
C14 vss    w2     0.074f
C15 w1     i1     0.370f
C16 nq     i0     0.056f
C17 w1     vdd    0.415f
C18 i1     i0     0.410f
C19 nq     w2     0.183f
C20 i1     w2     0.085f
C21 i0     vdd    0.035f
C22 vss    nq     0.069f
C24 nq     vss    0.018f
C25 w1     vss    0.034f
C26 i1     vss    0.040f
C27 i0     vss    0.032f
C29 w2     vss    0.069f
.ends
