magic
tech scmos
timestamp 1185094701
<< checkpaint >>
rect -22 -22 122 122
<< ab >>
rect 0 0 100 100
<< pwell >>
rect -4 -4 104 48
<< nwell >>
rect -4 48 104 104
<< polysilicon >>
rect 13 94 15 98
rect 37 90 39 95
rect 45 90 47 95
rect 59 94 61 98
rect 71 94 73 98
rect 83 94 85 98
rect 25 74 27 79
rect 13 43 15 56
rect 25 53 27 56
rect 19 52 27 53
rect 19 48 20 52
rect 24 48 27 52
rect 19 47 27 48
rect 11 42 21 43
rect 11 38 16 42
rect 20 38 21 42
rect 11 37 21 38
rect 11 34 13 37
rect 25 33 27 47
rect 37 43 39 56
rect 45 53 47 56
rect 59 53 61 56
rect 71 53 73 56
rect 83 53 85 56
rect 45 52 61 53
rect 45 48 48 52
rect 52 48 56 52
rect 60 48 61 52
rect 45 47 61 48
rect 67 52 75 53
rect 67 48 68 52
rect 72 48 75 52
rect 67 47 75 48
rect 79 52 85 53
rect 79 48 80 52
rect 84 49 85 52
rect 84 48 89 49
rect 79 47 89 48
rect 21 31 27 33
rect 33 42 41 43
rect 33 38 36 42
rect 40 38 41 42
rect 33 37 41 38
rect 21 28 23 31
rect 33 28 35 37
rect 45 31 47 47
rect 59 43 61 47
rect 73 43 75 47
rect 59 41 69 43
rect 73 41 77 43
rect 67 38 69 41
rect 75 38 77 41
rect 11 11 13 15
rect 21 8 23 13
rect 33 8 35 13
rect 45 11 47 16
rect 87 32 89 47
rect 87 8 89 13
rect 67 2 69 6
rect 75 2 77 6
<< ndiffusion >>
rect 3 33 11 34
rect 3 29 4 33
rect 8 29 11 33
rect 3 25 11 29
rect 3 21 4 25
rect 8 21 11 25
rect 3 20 11 21
rect 6 15 11 20
rect 13 28 19 34
rect 59 37 67 38
rect 59 33 60 37
rect 64 33 67 37
rect 59 32 67 33
rect 37 30 45 31
rect 37 28 38 30
rect 13 15 21 28
rect 15 13 21 15
rect 23 21 33 28
rect 23 17 26 21
rect 30 17 33 21
rect 23 13 33 17
rect 35 26 38 28
rect 42 26 45 30
rect 35 16 45 26
rect 47 22 52 31
rect 47 21 55 22
rect 47 17 50 21
rect 54 17 55 21
rect 47 16 55 17
rect 35 13 40 16
rect 15 9 19 13
rect 13 8 19 9
rect 13 4 14 8
rect 18 4 19 8
rect 13 3 19 4
rect 62 6 67 32
rect 69 6 75 38
rect 77 32 85 38
rect 77 22 87 32
rect 77 18 80 22
rect 84 18 87 22
rect 77 13 87 18
rect 89 31 97 32
rect 89 27 92 31
rect 96 27 97 31
rect 89 23 97 27
rect 89 19 92 23
rect 96 19 97 23
rect 89 18 97 19
rect 89 13 94 18
rect 77 12 85 13
rect 77 8 80 12
rect 84 8 85 12
rect 77 6 85 8
<< pdiffusion >>
rect 8 70 13 94
rect 5 69 13 70
rect 5 65 6 69
rect 10 65 13 69
rect 5 61 13 65
rect 5 57 6 61
rect 10 57 13 61
rect 5 56 13 57
rect 15 92 23 94
rect 15 88 18 92
rect 22 88 23 92
rect 49 92 59 94
rect 49 90 52 92
rect 15 82 23 88
rect 15 78 18 82
rect 22 78 23 82
rect 15 74 23 78
rect 32 74 37 90
rect 15 56 25 74
rect 27 62 37 74
rect 27 58 30 62
rect 34 58 37 62
rect 27 56 37 58
rect 39 56 45 90
rect 47 88 52 90
rect 56 88 59 92
rect 47 82 59 88
rect 47 78 52 82
rect 56 78 59 82
rect 47 56 59 78
rect 61 82 71 94
rect 61 78 64 82
rect 68 78 71 82
rect 61 72 71 78
rect 61 68 64 72
rect 68 68 71 72
rect 61 56 71 68
rect 73 92 83 94
rect 73 88 76 92
rect 80 88 83 92
rect 73 82 83 88
rect 73 78 76 82
rect 80 78 83 82
rect 73 56 83 78
rect 85 70 90 94
rect 85 69 93 70
rect 85 65 88 69
rect 92 65 93 69
rect 85 61 93 65
rect 85 57 88 61
rect 92 57 93 61
rect 85 56 93 57
<< metal1 >>
rect -2 92 102 100
rect -2 88 18 92
rect 22 88 52 92
rect 56 88 76 92
rect 80 88 102 92
rect 18 82 22 88
rect 18 77 22 78
rect 52 82 56 88
rect 52 77 56 78
rect 64 82 68 83
rect 6 69 12 73
rect 64 72 68 78
rect 76 82 80 88
rect 76 77 80 78
rect 10 65 12 69
rect 6 61 12 65
rect 10 57 12 61
rect 6 56 12 57
rect 8 34 12 56
rect 20 68 64 72
rect 68 68 84 72
rect 20 52 24 68
rect 20 47 24 48
rect 28 62 34 63
rect 28 58 30 62
rect 28 57 34 58
rect 38 58 72 63
rect 28 43 32 57
rect 38 43 42 58
rect 16 42 32 43
rect 20 38 32 42
rect 16 37 32 38
rect 36 42 42 43
rect 40 38 42 42
rect 36 37 42 38
rect 48 52 62 53
rect 52 48 56 52
rect 60 48 62 52
rect 48 47 62 48
rect 68 52 72 58
rect 68 47 72 48
rect 80 52 84 68
rect 4 33 12 34
rect 8 29 12 33
rect 4 27 12 29
rect 28 30 32 37
rect 4 25 8 27
rect 28 26 38 30
rect 42 26 43 30
rect 48 27 52 47
rect 80 37 84 48
rect 59 33 60 37
rect 64 33 84 37
rect 88 69 92 73
rect 88 61 92 65
rect 88 32 92 57
rect 88 31 96 32
rect 88 27 92 31
rect 92 23 96 27
rect 80 22 84 23
rect 4 20 8 21
rect 25 17 26 21
rect 30 17 50 21
rect 54 17 55 21
rect 92 18 96 19
rect 80 12 84 18
rect -2 8 80 12
rect 84 8 102 12
rect -2 4 14 8
rect 18 4 48 8
rect 52 4 102 8
rect -2 0 102 4
<< ntransistor >>
rect 11 15 13 34
rect 21 13 23 28
rect 33 13 35 28
rect 45 16 47 31
rect 67 6 69 38
rect 75 6 77 38
rect 87 13 89 32
<< ptransistor >>
rect 13 56 15 94
rect 25 56 27 74
rect 37 56 39 90
rect 45 56 47 90
rect 59 56 61 94
rect 71 56 73 94
rect 83 56 85 94
<< polycontact >>
rect 20 48 24 52
rect 16 38 20 42
rect 48 48 52 52
rect 56 48 60 52
rect 68 48 72 52
rect 80 48 84 52
rect 36 38 40 42
<< ndcontact >>
rect 4 29 8 33
rect 4 21 8 25
rect 60 33 64 37
rect 26 17 30 21
rect 38 26 42 30
rect 50 17 54 21
rect 14 4 18 8
rect 80 18 84 22
rect 92 27 96 31
rect 92 19 96 23
rect 80 8 84 12
<< pdcontact >>
rect 6 65 10 69
rect 6 57 10 61
rect 18 88 22 92
rect 18 78 22 82
rect 30 58 34 62
rect 52 88 56 92
rect 52 78 56 82
rect 64 78 68 82
rect 64 68 68 72
rect 76 88 80 92
rect 76 78 80 82
rect 88 65 92 69
rect 88 57 92 61
<< psubstratepcontact >>
rect 48 4 52 8
<< psubstratepdiff >>
rect 47 8 53 9
rect 47 4 48 8
rect 52 4 53 8
rect 47 3 53 4
<< labels >>
rlabel polysilicon 16 40 16 40 6 son
rlabel polycontact 23 50 23 50 6 con
rlabel polycontact 82 50 82 50 6 con
rlabel metal1 10 50 10 50 6 so
rlabel metal1 24 40 24 40 6 son
rlabel pdcontact 31 60 31 60 6 son
rlabel metal1 22 59 22 59 6 con
rlabel psubstratepcontact 50 6 50 6 6 vss
rlabel metal1 40 19 40 19 6 n2
rlabel metal1 35 28 35 28 6 son
rlabel metal1 50 40 50 40 6 a
rlabel metal1 40 50 40 50 6 b
rlabel metal1 50 60 50 60 6 b
rlabel metal1 50 94 50 94 6 vdd
rlabel metal1 60 50 60 50 6 a
rlabel metal1 70 55 70 55 6 b
rlabel metal1 60 60 60 60 6 b
rlabel metal1 66 75 66 75 6 con
rlabel metal1 71 35 71 35 6 con
rlabel metal1 90 50 90 50 6 co
rlabel metal1 82 52 82 52 6 con
rlabel metal1 52 70 52 70 6 con
<< end >>
