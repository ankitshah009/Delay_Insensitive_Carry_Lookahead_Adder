magic
tech scmos
timestamp 1179386477
<< checkpaint >>
rect -22 -25 78 105
<< ab >>
rect 0 0 56 80
<< pwell >>
rect -4 -7 60 36
<< nwell >>
rect -4 36 60 87
<< polysilicon >>
rect 9 70 11 74
rect 19 70 21 74
rect 30 70 32 74
rect 40 70 42 74
rect 9 39 11 42
rect 19 39 21 42
rect 30 39 32 42
rect 9 38 15 39
rect 9 34 10 38
rect 14 34 15 38
rect 9 33 15 34
rect 19 38 32 39
rect 19 34 26 38
rect 30 34 32 38
rect 40 39 42 42
rect 40 38 47 39
rect 40 35 42 38
rect 19 33 32 34
rect 13 29 15 33
rect 20 29 22 33
rect 30 29 32 33
rect 37 34 42 35
rect 46 34 47 38
rect 37 33 47 34
rect 37 29 39 33
rect 13 6 15 11
rect 20 6 22 11
rect 30 6 32 11
rect 37 6 39 11
<< ndiffusion >>
rect 4 15 13 29
rect 4 11 6 15
rect 10 11 13 15
rect 15 11 20 29
rect 22 22 30 29
rect 22 18 24 22
rect 28 18 30 22
rect 22 11 30 18
rect 32 11 37 29
rect 39 23 47 29
rect 39 19 41 23
rect 45 19 47 23
rect 39 16 47 19
rect 39 12 41 16
rect 45 12 47 16
rect 39 11 47 12
rect 4 9 11 11
<< pdiffusion >>
rect 2 69 9 70
rect 2 65 3 69
rect 7 65 9 69
rect 2 61 9 65
rect 2 57 3 61
rect 7 57 9 61
rect 2 42 9 57
rect 11 54 19 70
rect 11 50 13 54
rect 17 50 19 54
rect 11 47 19 50
rect 11 43 13 47
rect 17 43 19 47
rect 11 42 19 43
rect 21 69 30 70
rect 21 65 23 69
rect 27 65 30 69
rect 21 62 30 65
rect 21 58 23 62
rect 27 58 30 62
rect 21 42 30 58
rect 32 61 40 70
rect 32 57 34 61
rect 38 57 40 61
rect 32 54 40 57
rect 32 50 34 54
rect 38 50 40 54
rect 32 42 40 50
rect 42 69 50 70
rect 42 65 44 69
rect 48 65 50 69
rect 42 62 50 65
rect 42 58 44 62
rect 48 58 50 62
rect 42 42 50 58
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect -2 69 58 78
rect -2 68 3 69
rect 7 68 23 69
rect 3 61 7 65
rect 22 65 23 68
rect 27 68 44 69
rect 27 65 28 68
rect 22 62 28 65
rect 43 65 44 68
rect 48 68 58 69
rect 48 65 49 68
rect 22 58 23 62
rect 27 58 28 62
rect 34 61 39 63
rect 3 56 7 57
rect 38 57 39 61
rect 43 62 49 65
rect 43 58 44 62
rect 48 58 49 62
rect 34 54 39 57
rect 12 50 13 54
rect 17 50 34 54
rect 38 50 39 54
rect 12 47 18 50
rect 2 43 13 47
rect 17 43 18 47
rect 2 22 6 43
rect 25 42 39 46
rect 10 38 14 39
rect 25 38 31 42
rect 25 34 26 38
rect 30 34 31 38
rect 41 34 42 38
rect 46 34 47 38
rect 10 30 14 34
rect 41 30 47 34
rect 10 26 47 30
rect 2 18 24 22
rect 28 18 31 22
rect 40 19 41 23
rect 45 19 46 23
rect 40 16 46 19
rect 5 12 6 15
rect -2 11 6 12
rect 10 12 11 15
rect 40 12 41 16
rect 45 12 46 16
rect 10 11 58 12
rect -2 2 58 11
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
<< ntransistor >>
rect 13 11 15 29
rect 20 11 22 29
rect 30 11 32 29
rect 37 11 39 29
<< ptransistor >>
rect 9 42 11 70
rect 19 42 21 70
rect 30 42 32 70
rect 40 42 42 70
<< polycontact >>
rect 10 34 14 38
rect 26 34 30 38
rect 42 34 46 38
<< ndcontact >>
rect 6 11 10 15
rect 24 18 28 22
rect 41 19 45 23
rect 41 12 45 16
<< pdcontact >>
rect 3 65 7 69
rect 3 57 7 61
rect 13 50 17 54
rect 13 43 17 47
rect 23 65 27 69
rect 23 58 27 62
rect 34 57 38 61
rect 34 50 38 54
rect 44 65 48 69
rect 44 58 48 62
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
<< psubstratepdiff >>
rect 0 2 56 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 56 2
rect 0 -3 56 -2
<< nsubstratendiff >>
rect 0 82 56 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 56 82
rect 0 77 56 78
<< labels >>
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 20 12 20 6 z
rlabel polycontact 12 36 12 36 6 a
rlabel metal1 28 6 28 6 6 vss
rlabel metal1 20 20 20 20 6 z
rlabel metal1 20 28 20 28 6 a
rlabel metal1 28 28 28 28 6 a
rlabel metal1 28 20 28 20 6 z
rlabel metal1 28 40 28 40 6 b
rlabel metal1 28 52 28 52 6 z
rlabel metal1 20 52 20 52 6 z
rlabel metal1 28 74 28 74 6 vdd
rlabel metal1 36 28 36 28 6 a
rlabel metal1 44 32 44 32 6 a
rlabel metal1 36 44 36 44 6 b
rlabel metal1 36 56 36 56 6 z
<< end >>
