magic
tech scmos
timestamp 1180640054
<< checkpaint >>
rect -24 -26 94 126
<< ab >>
rect 0 0 70 100
<< pwell >>
rect -4 -6 74 49
<< nwell >>
rect -4 49 74 106
<< polysilicon >>
rect 33 94 35 98
rect 45 94 47 98
rect 57 94 59 98
rect 21 83 23 88
rect 57 63 59 66
rect 55 62 61 63
rect 55 58 56 62
rect 60 58 61 62
rect 55 57 61 58
rect 21 52 23 55
rect 33 52 35 55
rect 17 51 23 52
rect 17 48 18 51
rect 13 47 18 48
rect 22 47 23 51
rect 13 46 23 47
rect 27 51 35 52
rect 27 47 28 51
rect 32 48 35 51
rect 45 52 47 55
rect 45 51 53 52
rect 32 47 39 48
rect 27 46 39 47
rect 13 31 15 46
rect 37 39 39 46
rect 45 47 48 51
rect 52 47 53 51
rect 45 46 53 47
rect 45 39 47 46
rect 57 39 59 57
rect 13 12 15 17
rect 57 20 59 25
rect 37 2 39 6
rect 45 2 47 6
<< ndiffusion >>
rect 32 33 37 39
rect 29 32 37 33
rect 5 30 13 31
rect 5 26 6 30
rect 10 26 13 30
rect 5 22 13 26
rect 5 18 6 22
rect 10 18 13 22
rect 5 17 13 18
rect 15 22 23 31
rect 15 18 18 22
rect 22 18 23 22
rect 15 17 23 18
rect 29 28 30 32
rect 34 28 37 32
rect 29 22 37 28
rect 29 18 30 22
rect 34 18 37 22
rect 29 17 37 18
rect 32 6 37 17
rect 39 6 45 39
rect 47 32 57 39
rect 47 28 50 32
rect 54 28 57 32
rect 47 25 57 28
rect 59 38 67 39
rect 59 34 62 38
rect 66 34 67 38
rect 59 30 67 34
rect 59 26 62 30
rect 66 26 67 30
rect 59 25 67 26
rect 47 22 55 25
rect 47 18 50 22
rect 54 18 55 22
rect 47 12 55 18
rect 47 8 50 12
rect 54 8 55 12
rect 47 6 55 8
<< pdiffusion >>
rect 25 92 33 94
rect 25 88 26 92
rect 30 88 33 92
rect 25 83 33 88
rect 16 71 21 83
rect 13 70 21 71
rect 13 66 14 70
rect 18 66 21 70
rect 13 62 21 66
rect 13 58 14 62
rect 18 58 21 62
rect 13 57 21 58
rect 16 55 21 57
rect 23 82 33 83
rect 23 78 26 82
rect 30 78 33 82
rect 23 72 33 78
rect 23 68 26 72
rect 30 68 33 72
rect 23 55 33 68
rect 35 72 45 94
rect 35 68 38 72
rect 42 68 45 72
rect 35 62 45 68
rect 35 58 38 62
rect 42 58 45 62
rect 35 55 45 58
rect 47 92 57 94
rect 47 88 50 92
rect 54 88 57 92
rect 47 66 57 88
rect 59 73 64 94
rect 59 72 67 73
rect 59 68 62 72
rect 66 68 67 72
rect 59 66 67 68
rect 47 55 52 66
<< metal1 >>
rect -2 92 72 100
rect -2 88 26 92
rect 30 88 50 92
rect 54 88 72 92
rect 26 82 30 88
rect 26 72 30 78
rect 48 78 63 83
rect 14 70 18 71
rect 26 67 30 68
rect 38 72 42 73
rect 14 62 18 66
rect 38 62 42 68
rect 6 58 14 62
rect 18 58 32 62
rect 6 30 10 58
rect 18 51 22 53
rect 18 42 22 47
rect 28 51 32 58
rect 28 46 32 47
rect 18 38 33 42
rect 18 27 22 38
rect 38 33 42 58
rect 48 63 52 78
rect 61 72 68 73
rect 61 68 62 72
rect 66 68 68 72
rect 61 67 68 68
rect 48 62 60 63
rect 48 58 56 62
rect 48 57 60 58
rect 64 51 68 67
rect 47 47 48 51
rect 52 47 68 51
rect 62 38 66 47
rect 28 32 42 33
rect 28 28 30 32
rect 34 28 42 32
rect 28 27 42 28
rect 50 32 54 33
rect 6 22 10 26
rect 6 17 10 18
rect 18 22 22 23
rect 18 12 22 18
rect 28 22 34 27
rect 28 18 30 22
rect 28 17 34 18
rect 50 22 54 28
rect 62 30 66 34
rect 62 25 66 26
rect 50 12 54 18
rect -2 8 50 12
rect 54 8 72 12
rect -2 0 72 8
<< ntransistor >>
rect 13 17 15 31
rect 37 6 39 39
rect 45 6 47 39
rect 57 25 59 39
<< ptransistor >>
rect 21 55 23 83
rect 33 55 35 94
rect 45 55 47 94
rect 57 66 59 94
<< polycontact >>
rect 56 58 60 62
rect 18 47 22 51
rect 28 47 32 51
rect 48 47 52 51
<< ndcontact >>
rect 6 26 10 30
rect 6 18 10 22
rect 18 18 22 22
rect 30 28 34 32
rect 30 18 34 22
rect 50 28 54 32
rect 62 34 66 38
rect 62 26 66 30
rect 50 18 54 22
rect 50 8 54 12
<< pdcontact >>
rect 26 88 30 92
rect 14 66 18 70
rect 14 58 18 62
rect 26 78 30 82
rect 26 68 30 72
rect 38 68 42 72
rect 38 58 42 62
rect 50 88 54 92
rect 62 68 66 72
<< psubstratepcontact >>
rect 8 4 12 8
rect 18 4 22 8
<< nsubstratencontact >>
rect 4 92 8 96
rect 14 92 18 96
<< psubstratepdiff >>
rect 7 8 23 9
rect 7 4 8 8
rect 12 4 18 8
rect 22 4 23 8
rect 7 3 23 4
<< nsubstratendiff >>
rect 3 96 19 97
rect 3 92 4 96
rect 8 92 14 96
rect 18 92 19 96
rect 3 91 19 92
<< labels >>
rlabel metal1 8 39 8 39 6 bn
rlabel metal1 30 25 30 25 6 z
rlabel metal1 30 25 30 25 6 z
rlabel metal1 20 40 20 40 6 b
rlabel metal1 20 40 20 40 6 b
rlabel metal1 30 40 30 40 6 b
rlabel metal1 30 40 30 40 6 b
rlabel metal1 16 64 16 64 6 bn
rlabel metal1 35 6 35 6 6 vss
rlabel metal1 35 6 35 6 6 vss
rlabel metal1 40 50 40 50 6 z
rlabel metal1 40 50 40 50 6 z
rlabel metal1 50 70 50 70 6 a
rlabel metal1 50 70 50 70 6 a
rlabel metal1 35 94 35 94 6 vdd
rlabel metal1 35 94 35 94 6 vdd
rlabel metal1 57 49 57 49 6 an
rlabel metal1 64 38 64 38 6 an
rlabel pdcontact 64 70 64 70 6 an
rlabel metal1 60 80 60 80 6 a
rlabel metal1 60 80 60 80 6 a
<< end >>
