magic
tech scmos
timestamp 1185094854
<< checkpaint >>
rect -22 -22 92 122
<< ab >>
rect 0 0 70 100
<< pwell >>
rect -4 -4 74 48
<< nwell >>
rect -4 48 74 104
<< polysilicon >>
rect 11 94 13 98
rect 23 94 25 98
rect 35 94 37 98
rect 51 94 53 98
rect 61 72 67 73
rect 61 68 62 72
rect 66 68 67 72
rect 61 67 67 68
rect 11 47 13 56
rect 23 53 25 56
rect 35 53 37 56
rect 51 53 53 56
rect 65 53 67 67
rect 23 51 29 53
rect 35 51 43 53
rect 51 51 67 53
rect 27 47 29 51
rect 11 46 23 47
rect 11 44 18 46
rect 13 42 18 44
rect 22 42 23 46
rect 13 41 23 42
rect 27 46 33 47
rect 27 42 28 46
rect 32 42 33 46
rect 27 41 33 42
rect 41 43 43 51
rect 41 42 47 43
rect 13 32 15 41
rect 27 37 29 41
rect 41 38 42 42
rect 46 38 47 42
rect 41 37 47 38
rect 21 35 29 37
rect 21 32 23 35
rect 33 32 35 37
rect 45 32 47 37
rect 57 32 59 51
rect 13 11 15 15
rect 21 11 23 15
rect 33 5 35 15
rect 45 10 47 15
rect 57 5 59 15
rect 33 3 59 5
<< ndiffusion >>
rect 4 15 13 32
rect 15 15 21 32
rect 23 22 33 32
rect 23 18 26 22
rect 30 18 33 22
rect 23 15 33 18
rect 35 30 45 32
rect 35 26 38 30
rect 42 26 45 30
rect 35 22 45 26
rect 35 18 38 22
rect 42 18 45 22
rect 35 15 45 18
rect 47 15 57 32
rect 59 31 67 32
rect 59 27 62 31
rect 66 27 67 31
rect 59 23 67 27
rect 59 19 62 23
rect 66 19 67 23
rect 59 18 67 19
rect 59 15 64 18
rect 4 12 11 15
rect 4 8 6 12
rect 10 8 11 12
rect 4 7 11 8
rect 49 12 55 15
rect 49 8 50 12
rect 54 8 55 12
rect 49 7 55 8
<< pdiffusion >>
rect 6 83 11 94
rect 3 82 11 83
rect 3 78 4 82
rect 8 78 11 82
rect 3 77 11 78
rect 6 56 11 77
rect 13 72 23 94
rect 13 68 16 72
rect 20 68 23 72
rect 13 56 23 68
rect 25 72 35 94
rect 25 68 28 72
rect 32 68 35 72
rect 25 64 35 68
rect 25 60 28 64
rect 32 60 35 64
rect 25 56 35 60
rect 37 92 51 94
rect 37 88 44 92
rect 48 88 51 92
rect 37 82 51 88
rect 37 78 44 82
rect 48 78 51 82
rect 37 56 51 78
rect 53 62 58 94
rect 53 61 61 62
rect 53 57 56 61
rect 60 57 61 61
rect 53 56 61 57
<< metal1 >>
rect -2 92 72 100
rect -2 88 44 92
rect 48 88 72 92
rect 44 82 48 88
rect 3 78 4 82
rect 8 78 40 82
rect 8 72 23 73
rect 8 68 16 72
rect 20 68 23 72
rect 28 72 32 73
rect 8 23 12 68
rect 28 64 32 68
rect 18 60 28 62
rect 18 58 32 60
rect 18 46 22 58
rect 36 52 40 78
rect 44 77 48 78
rect 58 73 62 83
rect 48 72 67 73
rect 48 68 62 72
rect 66 68 67 72
rect 48 67 67 68
rect 48 57 52 67
rect 56 61 60 62
rect 56 52 60 57
rect 18 32 22 42
rect 28 48 66 52
rect 28 46 32 48
rect 28 41 32 42
rect 37 42 52 43
rect 37 38 42 42
rect 46 38 52 42
rect 18 30 42 32
rect 18 28 38 30
rect 8 22 32 23
rect 8 18 26 22
rect 30 18 32 22
rect 8 17 32 18
rect 38 22 42 26
rect 38 17 42 18
rect 48 17 52 38
rect 62 31 66 48
rect 62 23 66 27
rect 62 18 66 19
rect -2 8 6 12
rect 10 8 50 12
rect 54 8 72 12
rect -2 4 18 8
rect 22 4 72 8
rect -2 0 72 4
<< ntransistor >>
rect 13 15 15 32
rect 21 15 23 32
rect 33 15 35 32
rect 45 15 47 32
rect 57 15 59 32
<< ptransistor >>
rect 11 56 13 94
rect 23 56 25 94
rect 35 56 37 94
rect 51 56 53 94
<< polycontact >>
rect 62 68 66 72
rect 18 42 22 46
rect 28 42 32 46
rect 42 38 46 42
<< ndcontact >>
rect 26 18 30 22
rect 38 26 42 30
rect 38 18 42 22
rect 62 27 66 31
rect 62 19 66 23
rect 6 8 10 12
rect 50 8 54 12
<< pdcontact >>
rect 4 78 8 82
rect 16 68 20 72
rect 28 68 32 72
rect 28 60 32 64
rect 44 88 48 92
rect 44 78 48 82
rect 56 57 60 61
<< psubstratepcontact >>
rect 18 4 22 8
<< psubstratepdiff >>
rect 17 8 23 9
rect 17 4 18 8
rect 22 4 23 8
rect 17 3 23 4
<< labels >>
rlabel polysilicon 17 45 17 45 6 an
rlabel polycontact 30 44 30 44 6 bn
rlabel metal1 10 45 10 45 6 z
rlabel metal1 20 20 20 20 6 z
rlabel metal1 30 20 30 20 6 z
rlabel metal1 30 46 30 46 6 bn
rlabel polycontact 20 45 20 45 6 an
rlabel metal1 20 70 20 70 6 z
rlabel metal1 30 65 30 65 6 an
rlabel metal1 35 6 35 6 6 vss
rlabel metal1 40 24 40 24 6 an
rlabel metal1 50 30 50 30 6 a
rlabel metal1 40 40 40 40 6 a
rlabel metal1 50 65 50 65 6 b
rlabel metal1 35 94 35 94 6 vdd
rlabel metal1 21 80 21 80 6 bn
rlabel metal1 58 55 58 55 6 bn
rlabel metal1 64 35 64 35 6 bn
rlabel metal1 60 75 60 75 6 b
<< end >>
