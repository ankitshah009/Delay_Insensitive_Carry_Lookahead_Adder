.subckt aoi21v0x1 a1 a2 b vdd vss z
*   SPICE3 file   created from aoi21v0x1.ext -      technology: scmos
m00 vdd    vdd    w1     vdd p w=26u  l=2.3636u ad=147.333p pd=46u      as=182p     ps=66u
m01 w2     a1     vdd    vdd p w=26u  l=2.3636u ad=147.333p pd=46u      as=147.333p ps=46u
m02 w2     a2     vdd    vdd p w=26u  l=2.3636u ad=147.333p pd=46u      as=147.333p ps=46u
m03 z      b      w2     vdd p w=26u  l=2.3636u ad=182p     pd=66u      as=147.333p ps=46u
m04 vss    vss    w3     vss n w=18u  l=2.3636u ad=102p     pd=35.3333u as=126p     ps=50u
m05 w4     a1     vss    vss n w=18u  l=2.3636u ad=126p     pd=50u      as=102p     ps=35.3333u
m06 z      a2     w4     vss n w=18u  l=2.3636u ad=90p      pd=28u      as=126p     ps=50u
m07 vss    b      z      vss n w=18u  l=2.3636u ad=102p     pd=35.3333u as=90p      ps=28u
C0  b      a1     0.046f
C1  vss    z      0.069f
C2  a2     vdd    0.030f
C3  w4     a2     0.022f
C4  z      w2     0.110f
C5  z      b      0.224f
C6  vss    a2     0.020f
C7  z      a1     0.041f
C8  vss    vdd    0.047f
C9  w2     a2     0.016f
C10 w4     vss    0.136f
C11 w2     vdd    0.188f
C12 b      a2     0.183f
C13 w4     w2     0.012f
C14 b      vdd    0.014f
C15 a2     a1     0.129f
C16 a1     vdd    0.094f
C17 w4     a1     0.013f
C18 vss    b      0.032f
C19 z      a2     0.176f
C20 vss    a1     0.101f
C21 z      vdd    0.004f
C22 w2     a1     0.021f
C23 w4     z      0.040f
C24 w4     vss    0.004f
C26 z      vss    0.006f
C27 w2     vss    0.002f
C28 b      vss    0.062f
C29 a2     vss    0.062f
C30 a1     vss    0.061f
.ends
