.subckt nd2av0x2 a b vdd vss z
*   SPICE3 file   created from nd2av0x2.ext -      technology: scmos
m00 z      b      vdd    vdd p w=24u  l=2.3636u ad=96p      pd=32u      as=152.727p ps=48u
m01 vdd    an     z      vdd p w=24u  l=2.3636u ad=152.727p pd=48u      as=96p      ps=32u
m02 an     a      vdd    vdd p w=18u  l=2.3636u ad=102p     pd=50u      as=114.545p ps=36u
m03 w1     b      z      vss n w=19u  l=2.3636u ad=47.5p    pd=24u      as=107p     ps=52u
m04 vss    an     w1     vss n w=19u  l=2.3636u ad=141.143p pd=42.0714u as=47.5p    ps=24u
m05 an     a      vss    vss n w=9u   l=2.3636u ad=57p      pd=32u      as=66.8571p ps=19.9286u
C0  a      b      0.021f
C1  z      an     0.120f
C2  an     b      0.193f
C3  z      vdd    0.187f
C4  b      vdd    0.013f
C5  vss    a      0.017f
C6  vss    an     0.121f
C7  vss    vdd    0.003f
C8  a      an     0.292f
C9  w1     b      0.013f
C10 z      b      0.171f
C11 a      vdd    0.033f
C12 an     vdd    0.119f
C13 vss    w1     0.005f
C14 vss    z      0.076f
C15 a      z      0.018f
C16 vss    b      0.107f
C18 a      vss    0.018f
C19 z      vss    0.012f
C20 an     vss    0.020f
C21 b      vss    0.015f
.ends
