.subckt nr2v1x1 a b vdd vss z
*   SPICE3 file   created from nr2v1x1.ext -      technology: scmos
m00 w1     b      z      vdd p w=28u  l=2.3636u ad=70p      pd=33u      as=166p     ps=70u
m01 vdd    a      w1     vdd p w=28u  l=2.3636u ad=252p     pd=74u      as=70p      ps=33u
m02 z      b      vss    vss n w=14u  l=2.3636u ad=56p      pd=22u      as=130p     ps=50u
m03 vss    a      z      vss n w=14u  l=2.3636u ad=130p     pd=50u      as=56p      ps=22u
C0  a      b      0.134f
C1  vdd    z      0.053f
C2  vss    a      0.054f
C3  vdd    b      0.023f
C4  z      b      0.118f
C5  vss    vdd    0.004f
C6  vdd    w1     0.005f
C7  vss    z      0.160f
C8  vdd    a      0.018f
C9  vss    b      0.018f
C10 z      a      0.042f
C11 w1     b      0.007f
C14 z      vss    0.013f
C15 a      vss    0.021f
C16 b      vss    0.018f
.ends
