magic
tech scmos
timestamp 1179386605
<< checkpaint >>
rect -22 -22 134 94
<< ab >>
rect 0 0 112 72
<< pwell >>
rect -4 -4 116 32
<< nwell >>
rect -4 32 116 76
<< polysilicon >>
rect 10 58 12 63
rect 20 58 22 63
rect 30 58 32 63
rect 40 58 42 63
rect 50 58 52 63
rect 60 58 62 63
rect 70 58 72 63
rect 80 58 82 63
rect 90 58 92 63
rect 10 35 12 38
rect 20 35 22 38
rect 30 35 32 38
rect 10 34 32 35
rect 10 30 11 34
rect 15 30 18 34
rect 22 30 32 34
rect 10 29 32 30
rect 10 26 12 29
rect 20 26 22 29
rect 30 26 32 29
rect 40 35 42 38
rect 50 35 52 38
rect 60 35 62 38
rect 40 34 62 35
rect 40 30 42 34
rect 46 30 50 34
rect 54 30 62 34
rect 40 29 62 30
rect 40 26 42 29
rect 50 26 52 29
rect 60 26 62 29
rect 70 35 72 38
rect 80 35 82 38
rect 90 35 92 38
rect 70 34 103 35
rect 70 30 98 34
rect 102 30 103 34
rect 70 29 103 30
rect 70 26 72 29
rect 80 26 82 29
rect 90 26 92 29
rect 101 26 103 29
rect 90 11 92 16
rect 101 11 103 16
rect 10 2 12 6
rect 20 2 22 6
rect 30 2 32 6
rect 40 2 42 6
rect 50 2 52 6
rect 60 2 62 6
rect 70 2 72 6
rect 80 2 82 6
<< ndiffusion >>
rect 2 18 10 26
rect 2 14 3 18
rect 7 14 10 18
rect 2 11 10 14
rect 2 7 3 11
rect 7 7 10 11
rect 2 6 10 7
rect 12 25 20 26
rect 12 21 14 25
rect 18 21 20 25
rect 12 18 20 21
rect 12 14 14 18
rect 18 14 20 18
rect 12 6 20 14
rect 22 11 30 26
rect 22 7 24 11
rect 28 7 30 11
rect 22 6 30 7
rect 32 18 40 26
rect 32 14 34 18
rect 38 14 40 18
rect 32 6 40 14
rect 42 25 50 26
rect 42 21 44 25
rect 48 21 50 25
rect 42 6 50 21
rect 52 18 60 26
rect 52 14 54 18
rect 58 14 60 18
rect 52 6 60 14
rect 62 25 70 26
rect 62 21 64 25
rect 68 21 70 25
rect 62 18 70 21
rect 62 14 64 18
rect 68 14 70 18
rect 62 6 70 14
rect 72 25 80 26
rect 72 21 74 25
rect 78 21 80 25
rect 72 6 80 21
rect 82 21 90 26
rect 82 17 84 21
rect 88 17 90 21
rect 82 16 90 17
rect 92 25 101 26
rect 92 21 94 25
rect 98 21 101 25
rect 92 16 101 21
rect 103 22 108 26
rect 103 21 110 22
rect 103 17 105 21
rect 109 17 110 21
rect 103 16 110 17
rect 82 6 87 16
<< pdiffusion >>
rect 2 57 10 58
rect 2 53 3 57
rect 7 53 10 57
rect 2 50 10 53
rect 2 46 3 50
rect 7 46 10 50
rect 2 38 10 46
rect 12 50 20 58
rect 12 46 14 50
rect 18 46 20 50
rect 12 43 20 46
rect 12 39 14 43
rect 18 39 20 43
rect 12 38 20 39
rect 22 57 30 58
rect 22 53 24 57
rect 28 53 30 57
rect 22 50 30 53
rect 22 46 24 50
rect 28 46 30 50
rect 22 38 30 46
rect 32 50 40 58
rect 32 46 34 50
rect 38 46 40 50
rect 32 43 40 46
rect 32 39 34 43
rect 38 39 40 43
rect 32 38 40 39
rect 42 57 50 58
rect 42 53 44 57
rect 48 53 50 57
rect 42 50 50 53
rect 42 46 44 50
rect 48 46 50 50
rect 42 38 50 46
rect 52 50 60 58
rect 52 46 54 50
rect 58 46 60 50
rect 52 43 60 46
rect 52 39 54 43
rect 58 39 60 43
rect 52 38 60 39
rect 62 57 70 58
rect 62 53 64 57
rect 68 53 70 57
rect 62 50 70 53
rect 62 46 64 50
rect 68 46 70 50
rect 62 38 70 46
rect 72 50 80 58
rect 72 46 74 50
rect 78 46 80 50
rect 72 43 80 46
rect 72 39 74 43
rect 78 39 80 43
rect 72 38 80 39
rect 82 57 90 58
rect 82 53 84 57
rect 88 53 90 57
rect 82 50 90 53
rect 82 46 84 50
rect 88 46 90 50
rect 82 38 90 46
rect 92 51 97 58
rect 92 50 99 51
rect 92 46 94 50
rect 98 46 99 50
rect 92 43 99 46
rect 92 39 94 43
rect 98 39 99 43
rect 92 38 99 39
<< metal1 >>
rect -2 68 114 72
rect -2 64 104 68
rect 108 64 114 68
rect 2 57 8 64
rect 2 53 3 57
rect 7 53 8 57
rect 2 50 8 53
rect 23 57 29 64
rect 23 53 24 57
rect 28 53 29 57
rect 2 46 3 50
rect 7 46 8 50
rect 14 50 18 51
rect 23 50 29 53
rect 43 57 49 64
rect 43 53 44 57
rect 48 53 49 57
rect 23 46 24 50
rect 28 46 29 50
rect 34 50 38 51
rect 43 50 49 53
rect 63 57 69 64
rect 63 53 64 57
rect 68 53 69 57
rect 43 46 44 50
rect 48 46 49 50
rect 54 50 58 51
rect 63 50 69 53
rect 63 46 64 50
rect 68 46 69 50
rect 74 50 78 59
rect 83 57 89 64
rect 83 53 84 57
rect 88 53 89 57
rect 83 50 89 53
rect 83 46 84 50
rect 88 46 89 50
rect 94 50 98 51
rect 14 43 18 46
rect 2 34 6 43
rect 34 43 38 46
rect 18 39 34 42
rect 54 43 58 46
rect 38 39 54 42
rect 74 43 78 46
rect 94 43 98 46
rect 58 39 74 42
rect 90 42 94 43
rect 78 39 94 42
rect 14 38 98 39
rect 74 37 95 38
rect 2 30 11 34
rect 15 30 18 34
rect 22 30 23 34
rect 33 30 42 34
rect 46 30 50 34
rect 54 30 55 34
rect 2 21 6 30
rect 13 25 18 26
rect 13 21 14 25
rect 33 22 39 30
rect 74 25 78 37
rect 43 21 44 25
rect 48 21 64 25
rect 68 21 69 25
rect 13 18 18 21
rect 64 18 69 21
rect 91 25 95 37
rect 106 35 110 51
rect 98 34 110 35
rect 102 30 110 34
rect 98 29 110 30
rect 74 20 78 21
rect 84 21 88 22
rect 91 21 94 25
rect 98 21 99 25
rect 105 21 109 22
rect 2 14 3 18
rect 7 14 8 18
rect 13 14 14 18
rect 18 14 34 18
rect 38 14 54 18
rect 58 14 59 18
rect 68 17 69 18
rect 68 14 109 17
rect 2 11 8 14
rect 64 13 109 14
rect 2 8 3 11
rect -2 7 3 8
rect 7 8 8 11
rect 23 8 24 11
rect 7 7 24 8
rect 28 8 29 11
rect 28 7 96 8
rect -2 4 96 7
rect 100 4 104 8
rect 108 4 114 8
rect -2 0 114 4
<< ntransistor >>
rect 10 6 12 26
rect 20 6 22 26
rect 30 6 32 26
rect 40 6 42 26
rect 50 6 52 26
rect 60 6 62 26
rect 70 6 72 26
rect 80 6 82 26
rect 90 16 92 26
rect 101 16 103 26
<< ptransistor >>
rect 10 38 12 58
rect 20 38 22 58
rect 30 38 32 58
rect 40 38 42 58
rect 50 38 52 58
rect 60 38 62 58
rect 70 38 72 58
rect 80 38 82 58
rect 90 38 92 58
<< polycontact >>
rect 11 30 15 34
rect 18 30 22 34
rect 42 30 46 34
rect 50 30 54 34
rect 98 30 102 34
<< ndcontact >>
rect 3 14 7 18
rect 3 7 7 11
rect 14 21 18 25
rect 14 14 18 18
rect 24 7 28 11
rect 34 14 38 18
rect 44 21 48 25
rect 54 14 58 18
rect 64 21 68 25
rect 64 14 68 18
rect 74 21 78 25
rect 84 17 88 21
rect 94 21 98 25
rect 105 17 109 21
<< pdcontact >>
rect 3 53 7 57
rect 3 46 7 50
rect 14 46 18 50
rect 14 39 18 43
rect 24 53 28 57
rect 24 46 28 50
rect 34 46 38 50
rect 34 39 38 43
rect 44 53 48 57
rect 44 46 48 50
rect 54 46 58 50
rect 54 39 58 43
rect 64 53 68 57
rect 64 46 68 50
rect 74 46 78 50
rect 74 39 78 43
rect 84 53 88 57
rect 84 46 88 50
rect 94 46 98 50
rect 94 39 98 43
<< psubstratepcontact >>
rect 96 4 100 8
rect 104 4 108 8
<< nsubstratencontact >>
rect 104 64 108 68
<< psubstratepdiff >>
rect 95 8 109 9
rect 95 4 96 8
rect 100 4 104 8
rect 108 4 109 8
rect 95 3 109 4
<< nsubstratendiff >>
rect 103 68 109 69
rect 103 64 104 68
rect 108 64 109 68
rect 103 63 109 64
<< labels >>
rlabel metal1 15 20 15 20 6 n1
rlabel metal1 4 32 4 32 6 a
rlabel polycontact 12 32 12 32 6 a
rlabel metal1 36 28 36 28 6 b
rlabel polycontact 20 32 20 32 6 a
rlabel metal1 20 40 20 40 6 z
rlabel metal1 28 40 28 40 6 z
rlabel metal1 36 44 36 44 6 z
rlabel metal1 56 4 56 4 6 vss
rlabel ndcontact 36 16 36 16 6 n1
rlabel polycontact 52 32 52 32 6 b
rlabel polycontact 44 32 44 32 6 b
rlabel metal1 44 40 44 40 6 z
rlabel metal1 52 40 52 40 6 z
rlabel metal1 60 40 60 40 6 z
rlabel metal1 56 68 56 68 6 vdd
rlabel metal1 86 17 86 17 6 n2
rlabel metal1 66 19 66 19 6 n2
rlabel metal1 56 23 56 23 6 n2
rlabel metal1 68 40 68 40 6 z
rlabel pdcontact 76 40 76 40 6 z
rlabel metal1 84 40 84 40 6 z
rlabel metal1 107 17 107 17 6 n2
rlabel polycontact 100 32 100 32 6 c
rlabel metal1 92 40 92 40 6 z
rlabel metal1 108 40 108 40 6 c
<< end >>
