magic
tech scmos
timestamp 1185094650
<< checkpaint >>
rect -22 -22 92 122
<< ab >>
rect 0 0 70 100
<< pwell >>
rect -4 -4 74 48
<< nwell >>
rect -4 48 74 104
<< polysilicon >>
rect 11 93 13 98
rect 33 93 35 98
rect 45 93 47 98
rect 57 93 59 98
rect 11 52 13 55
rect 33 52 35 55
rect 45 52 47 55
rect 57 52 59 55
rect 11 51 22 52
rect 11 50 17 51
rect 15 47 17 50
rect 21 47 22 51
rect 15 46 22 47
rect 33 51 41 52
rect 33 47 36 51
rect 40 47 41 51
rect 33 46 41 47
rect 45 51 53 52
rect 45 47 48 51
rect 52 47 53 51
rect 45 46 53 47
rect 57 51 63 52
rect 57 47 58 51
rect 62 47 63 51
rect 57 46 63 47
rect 15 35 17 46
rect 33 35 35 46
rect 45 35 47 46
rect 57 40 59 46
rect 53 38 59 40
rect 53 35 55 38
rect 33 20 35 25
rect 15 11 17 16
rect 45 13 47 18
rect 53 13 55 18
<< ndiffusion >>
rect 7 34 15 35
rect 7 30 8 34
rect 12 30 15 34
rect 7 26 15 30
rect 7 22 8 26
rect 12 22 15 26
rect 7 21 15 22
rect 10 16 15 21
rect 17 32 33 35
rect 17 28 20 32
rect 24 28 33 32
rect 17 25 33 28
rect 35 34 45 35
rect 35 30 38 34
rect 42 30 45 34
rect 35 25 45 30
rect 17 22 31 25
rect 17 18 20 22
rect 24 18 31 22
rect 40 18 45 25
rect 47 18 53 35
rect 55 32 64 35
rect 55 28 58 32
rect 62 28 64 32
rect 55 23 64 28
rect 55 19 58 23
rect 62 19 64 23
rect 55 18 64 19
rect 17 16 31 18
<< pdiffusion >>
rect 6 73 11 93
rect 3 72 11 73
rect 3 68 4 72
rect 8 68 11 72
rect 3 62 11 68
rect 3 58 4 62
rect 8 58 11 62
rect 3 57 11 58
rect 6 55 11 57
rect 13 92 21 93
rect 13 88 16 92
rect 20 88 21 92
rect 13 82 21 88
rect 13 78 16 82
rect 20 78 21 82
rect 13 75 21 78
rect 13 55 19 75
rect 28 69 33 93
rect 25 68 33 69
rect 25 64 26 68
rect 30 64 33 68
rect 25 60 33 64
rect 25 56 26 60
rect 30 56 33 60
rect 25 55 33 56
rect 35 82 45 93
rect 35 78 38 82
rect 42 78 45 82
rect 35 55 45 78
rect 47 92 57 93
rect 47 88 50 92
rect 54 88 57 92
rect 47 55 57 88
rect 59 83 64 93
rect 59 82 67 83
rect 59 78 62 82
rect 66 78 67 82
rect 59 77 67 78
rect 59 55 64 77
<< metal1 >>
rect -2 92 72 100
rect -2 88 16 92
rect 20 88 50 92
rect 54 88 72 92
rect 16 82 20 88
rect 37 78 38 82
rect 42 78 62 82
rect 66 78 67 82
rect 16 77 20 78
rect 4 72 22 73
rect 8 68 22 72
rect 4 67 22 68
rect 26 68 30 69
rect 8 63 12 67
rect 4 62 12 63
rect 8 58 12 62
rect 4 57 12 58
rect 8 34 12 57
rect 26 60 30 64
rect 26 51 30 56
rect 38 68 53 73
rect 38 52 42 68
rect 58 63 62 73
rect 16 47 17 51
rect 21 47 30 51
rect 26 42 30 47
rect 36 51 42 52
rect 40 47 42 51
rect 36 46 42 47
rect 48 57 62 63
rect 48 51 52 57
rect 48 46 52 47
rect 57 51 63 52
rect 57 47 58 51
rect 62 47 63 51
rect 57 42 63 47
rect 26 38 42 42
rect 38 34 42 38
rect 8 26 12 30
rect 8 17 12 22
rect 20 32 24 33
rect 38 29 42 30
rect 47 38 63 42
rect 20 22 24 28
rect 47 18 53 38
rect 58 32 62 33
rect 58 23 62 28
rect 20 12 24 18
rect 58 12 62 19
rect -2 8 72 12
rect -2 4 8 8
rect 12 4 18 8
rect 22 4 72 8
rect -2 0 72 4
<< ntransistor >>
rect 15 16 17 35
rect 33 25 35 35
rect 45 18 47 35
rect 53 18 55 35
<< ptransistor >>
rect 11 55 13 93
rect 33 55 35 93
rect 45 55 47 93
rect 57 55 59 93
<< polycontact >>
rect 17 47 21 51
rect 36 47 40 51
rect 48 47 52 51
rect 58 47 62 51
<< ndcontact >>
rect 8 30 12 34
rect 8 22 12 26
rect 20 28 24 32
rect 38 30 42 34
rect 20 18 24 22
rect 58 28 62 32
rect 58 19 62 23
<< pdcontact >>
rect 4 68 8 72
rect 4 58 8 62
rect 16 88 20 92
rect 16 78 20 82
rect 26 64 30 68
rect 26 56 30 60
rect 38 78 42 82
rect 50 88 54 92
rect 62 78 66 82
<< psubstratepcontact >>
rect 8 4 12 8
rect 18 4 22 8
<< psubstratepdiff >>
rect 7 8 23 9
rect 7 4 8 8
rect 12 4 18 8
rect 22 4 23 8
rect 7 3 23 4
<< labels >>
rlabel polycontact 18 49 18 49 6 zn
rlabel metal1 10 45 10 45 6 z
rlabel metal1 20 70 20 70 6 z
rlabel metal1 35 6 35 6 6 vss
rlabel metal1 23 49 23 49 6 zn
rlabel metal1 28 53 28 53 6 zn
rlabel metal1 35 94 35 94 6 vdd
rlabel metal1 50 30 50 30 6 a1
rlabel metal1 40 35 40 35 6 zn
rlabel metal1 50 55 50 55 6 a2
rlabel metal1 40 60 40 60 6 b
rlabel metal1 50 70 50 70 6 b
rlabel metal1 60 45 60 45 6 a1
rlabel metal1 60 65 60 65 6 a2
rlabel metal1 52 80 52 80 6 n2
<< end >>
