.subckt rowend_x0 vdd vss
*   SPICE3 file   created from rowend_x0.ext -      technology: scmos
.ends
