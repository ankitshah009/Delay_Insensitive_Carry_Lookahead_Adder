magic
tech scmos
timestamp 1179386942
<< checkpaint >>
rect -22 -25 134 105
<< ab >>
rect 0 0 112 80
<< pwell >>
rect -4 -7 116 36
<< nwell >>
rect -4 36 116 87
<< polysilicon >>
rect 14 69 16 74
rect 21 69 23 74
rect 28 69 30 74
rect 35 69 37 74
rect 47 69 49 74
rect 54 69 56 74
rect 61 69 63 74
rect 68 69 70 74
rect 78 69 80 74
rect 85 69 87 74
rect 92 69 94 74
rect 99 69 101 74
rect 14 41 16 44
rect 9 40 16 41
rect 9 36 10 40
rect 14 36 16 40
rect 9 35 16 36
rect 10 22 12 35
rect 21 31 23 44
rect 17 30 23 31
rect 17 26 18 30
rect 22 26 23 30
rect 17 25 23 26
rect 28 31 30 44
rect 35 39 37 44
rect 47 39 49 42
rect 35 38 49 39
rect 35 37 39 38
rect 38 34 39 37
rect 43 37 49 38
rect 43 34 44 37
rect 38 33 44 34
rect 28 30 34 31
rect 28 26 29 30
rect 33 26 34 30
rect 28 25 34 26
rect 20 22 22 25
rect 32 22 34 25
rect 42 22 44 33
rect 54 31 56 42
rect 61 33 63 42
rect 68 39 70 42
rect 78 39 80 42
rect 68 38 81 39
rect 68 37 76 38
rect 75 34 76 37
rect 80 34 81 38
rect 75 33 81 34
rect 61 32 71 33
rect 61 31 66 32
rect 48 30 56 31
rect 48 26 49 30
rect 53 26 56 30
rect 65 28 66 31
rect 70 29 71 32
rect 85 29 87 42
rect 70 28 87 29
rect 65 27 87 28
rect 48 25 56 26
rect 54 23 56 25
rect 92 23 94 42
rect 10 6 12 11
rect 20 6 22 11
rect 54 21 94 23
rect 99 23 101 42
rect 99 22 105 23
rect 99 18 100 22
rect 104 18 105 22
rect 99 17 105 18
rect 32 6 34 11
rect 42 6 44 11
<< ndiffusion >>
rect 2 12 10 22
rect 2 8 3 12
rect 7 11 10 12
rect 12 21 20 22
rect 12 17 14 21
rect 18 17 20 21
rect 12 11 20 17
rect 22 12 32 22
rect 22 11 25 12
rect 7 8 8 11
rect 2 7 8 8
rect 24 8 25 11
rect 29 11 32 12
rect 34 21 42 22
rect 34 17 36 21
rect 40 17 42 21
rect 34 11 42 17
rect 44 12 52 22
rect 44 11 47 12
rect 29 8 30 11
rect 24 7 30 8
rect 46 8 47 11
rect 51 8 52 12
rect 46 7 52 8
<< pdiffusion >>
rect 39 72 45 73
rect 39 69 40 72
rect 9 63 14 69
rect 7 62 14 63
rect 7 58 8 62
rect 12 58 14 62
rect 7 57 14 58
rect 9 44 14 57
rect 16 44 21 69
rect 23 44 28 69
rect 30 44 35 69
rect 37 68 40 69
rect 44 69 45 72
rect 44 68 47 69
rect 37 44 47 68
rect 39 42 47 44
rect 49 42 54 69
rect 56 42 61 69
rect 63 42 68 69
rect 70 62 78 69
rect 70 58 72 62
rect 76 58 78 62
rect 70 42 78 58
rect 80 42 85 69
rect 87 42 92 69
rect 94 42 99 69
rect 101 68 108 69
rect 101 64 103 68
rect 107 64 108 68
rect 101 61 108 64
rect 101 57 103 61
rect 107 57 108 61
rect 101 42 108 57
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect -2 72 114 78
rect -2 68 40 72
rect 44 68 114 72
rect 102 64 103 68
rect 107 64 108 68
rect 2 58 8 62
rect 12 58 72 62
rect 76 58 79 62
rect 102 61 108 64
rect 2 23 6 58
rect 102 57 103 61
rect 107 57 108 61
rect 10 50 80 54
rect 10 40 14 50
rect 10 33 14 36
rect 18 42 70 46
rect 18 30 22 42
rect 38 34 39 38
rect 43 34 62 38
rect 28 26 29 30
rect 33 26 49 30
rect 53 26 54 30
rect 18 25 22 26
rect 2 17 14 23
rect 33 21 41 22
rect 18 17 36 21
rect 40 17 41 21
rect 50 17 54 26
rect 58 22 62 34
rect 66 32 70 42
rect 74 38 80 50
rect 74 34 76 38
rect 74 33 80 34
rect 66 27 70 28
rect 58 18 100 22
rect 104 18 105 22
rect -2 8 3 12
rect 7 8 25 12
rect 29 8 47 12
rect 51 8 114 12
rect -2 2 114 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
<< ntransistor >>
rect 10 11 12 22
rect 20 11 22 22
rect 32 11 34 22
rect 42 11 44 22
<< ptransistor >>
rect 14 44 16 69
rect 21 44 23 69
rect 28 44 30 69
rect 35 44 37 69
rect 47 42 49 69
rect 54 42 56 69
rect 61 42 63 69
rect 68 42 70 69
rect 78 42 80 69
rect 85 42 87 69
rect 92 42 94 69
rect 99 42 101 69
<< polycontact >>
rect 10 36 14 40
rect 18 26 22 30
rect 39 34 43 38
rect 29 26 33 30
rect 76 34 80 38
rect 49 26 53 30
rect 66 28 70 32
rect 100 18 104 22
<< ndcontact >>
rect 3 8 7 12
rect 14 17 18 21
rect 25 8 29 12
rect 36 17 40 21
rect 47 8 51 12
<< pdcontact >>
rect 8 58 12 62
rect 40 68 44 72
rect 72 58 76 62
rect 103 64 107 68
rect 103 57 107 61
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
rect 90 -2 94 2
rect 98 -2 102 2
rect 106 -2 110 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
rect 90 78 94 82
rect 98 78 102 82
rect 106 78 110 82
<< psubstratepdiff >>
rect 0 2 112 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 112 2
rect 0 -3 112 -2
<< nsubstratendiff >>
rect 0 82 112 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 112 82
rect 0 77 112 78
<< labels >>
rlabel metal1 12 20 12 20 6 z
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 40 12 40 6 d
rlabel metal1 12 60 12 60 6 z
rlabel metal1 36 20 36 20 6 z
rlabel metal1 36 28 36 28 6 b
rlabel metal1 20 32 20 32 6 c
rlabel metal1 28 44 28 44 6 c
rlabel metal1 36 44 36 44 6 c
rlabel metal1 28 52 28 52 6 d
rlabel metal1 36 52 36 52 6 d
rlabel metal1 20 52 20 52 6 d
rlabel metal1 20 60 20 60 6 z
rlabel metal1 28 60 28 60 6 z
rlabel metal1 36 60 36 60 6 z
rlabel metal1 56 6 56 6 6 vss
rlabel metal1 44 28 44 28 6 b
rlabel metal1 52 20 52 20 6 b
rlabel metal1 60 28 60 28 6 a
rlabel metal1 44 36 44 36 6 a
rlabel metal1 44 44 44 44 6 c
rlabel metal1 52 36 52 36 6 a
rlabel metal1 52 44 52 44 6 c
rlabel metal1 60 44 60 44 6 c
rlabel metal1 52 52 52 52 6 d
rlabel metal1 60 52 60 52 6 d
rlabel metal1 44 52 44 52 6 d
rlabel metal1 44 60 44 60 6 z
rlabel metal1 52 60 52 60 6 z
rlabel metal1 60 60 60 60 6 z
rlabel metal1 56 74 56 74 6 vdd
rlabel metal1 68 20 68 20 6 a
rlabel metal1 76 20 76 20 6 a
rlabel metal1 84 20 84 20 6 a
rlabel metal1 68 36 68 36 6 c
rlabel metal1 76 44 76 44 6 d
rlabel metal1 68 52 68 52 6 d
rlabel metal1 68 60 68 60 6 z
rlabel metal1 76 60 76 60 6 z
rlabel metal1 92 20 92 20 6 a
rlabel metal1 100 20 100 20 6 a
<< end >>
