magic
tech scmos
timestamp 1179385929
<< checkpaint >>
rect -22 -22 94 94
<< ab >>
rect 0 0 72 72
<< pwell >>
rect -4 -4 76 32
<< nwell >>
rect -4 32 76 76
<< polysilicon >>
rect 9 66 11 70
rect 19 66 21 70
rect 29 66 31 70
rect 39 66 41 70
rect 49 66 51 70
rect 59 57 61 61
rect 9 35 11 38
rect 19 35 21 38
rect 29 35 31 38
rect 39 35 41 38
rect 9 34 41 35
rect 9 33 36 34
rect 22 26 24 33
rect 32 30 36 33
rect 40 30 41 34
rect 32 29 41 30
rect 49 35 51 38
rect 59 35 61 38
rect 49 34 61 35
rect 49 30 50 34
rect 54 33 61 34
rect 54 30 55 33
rect 49 29 55 30
rect 32 26 34 29
rect 22 2 24 6
rect 32 2 34 6
<< ndiffusion >>
rect 14 19 22 26
rect 14 15 16 19
rect 20 15 22 19
rect 14 11 22 15
rect 14 7 16 11
rect 20 7 22 11
rect 14 6 22 7
rect 24 25 32 26
rect 24 21 26 25
rect 30 21 32 25
rect 24 18 32 21
rect 24 14 26 18
rect 30 14 32 18
rect 24 6 32 14
rect 34 19 42 26
rect 34 15 36 19
rect 40 15 42 19
rect 34 11 42 15
rect 34 7 36 11
rect 40 7 42 11
rect 34 6 42 7
<< pdiffusion >>
rect 2 65 9 66
rect 2 61 3 65
rect 7 61 9 65
rect 2 58 9 61
rect 2 54 3 58
rect 7 54 9 58
rect 2 51 9 54
rect 2 47 3 51
rect 7 47 9 51
rect 2 38 9 47
rect 11 50 19 66
rect 11 46 13 50
rect 17 46 19 50
rect 11 43 19 46
rect 11 39 13 43
rect 17 39 19 43
rect 11 38 19 39
rect 21 65 29 66
rect 21 61 23 65
rect 27 61 29 65
rect 21 57 29 61
rect 21 53 23 57
rect 27 53 29 57
rect 21 38 29 53
rect 31 50 39 66
rect 31 46 33 50
rect 37 46 39 50
rect 31 43 39 46
rect 31 39 33 43
rect 37 39 39 43
rect 31 38 39 39
rect 41 65 49 66
rect 41 61 43 65
rect 47 61 49 65
rect 41 57 49 61
rect 41 53 43 57
rect 47 53 49 57
rect 41 38 49 53
rect 51 57 56 66
rect 51 50 59 57
rect 51 46 53 50
rect 57 46 59 50
rect 51 43 59 46
rect 51 39 53 43
rect 57 39 59 43
rect 51 38 59 39
rect 61 56 68 57
rect 61 52 63 56
rect 67 52 68 56
rect 61 49 68 52
rect 61 45 63 49
rect 67 45 68 49
rect 61 38 68 45
<< metal1 >>
rect -2 68 74 72
rect -2 65 62 68
rect -2 64 3 65
rect 7 64 23 65
rect 3 58 7 61
rect 3 51 7 54
rect 27 64 43 65
rect 23 57 27 61
rect 23 52 27 53
rect 47 64 62 65
rect 66 64 74 68
rect 43 57 47 61
rect 43 52 47 53
rect 62 56 68 64
rect 62 52 63 56
rect 67 52 68 56
rect 3 46 7 47
rect 13 50 17 51
rect 13 43 17 46
rect 9 39 13 42
rect 33 50 38 51
rect 37 46 38 50
rect 33 43 38 46
rect 17 39 33 42
rect 37 42 38 43
rect 53 50 57 51
rect 62 49 68 52
rect 62 46 63 49
rect 53 43 57 46
rect 67 46 68 49
rect 37 39 53 42
rect 57 39 63 42
rect 9 38 63 39
rect 26 25 30 38
rect 35 30 36 34
rect 40 30 50 34
rect 54 30 55 34
rect 49 22 55 30
rect 16 19 20 20
rect 16 11 20 15
rect 26 18 30 21
rect 26 13 30 14
rect 36 19 40 20
rect -2 4 4 8
rect 8 7 16 8
rect 36 11 40 15
rect 20 7 36 8
rect 40 7 63 8
rect 8 4 63 7
rect 67 4 74 8
rect -2 0 74 4
<< ntransistor >>
rect 22 6 24 26
rect 32 6 34 26
<< ptransistor >>
rect 9 38 11 66
rect 19 38 21 66
rect 29 38 31 66
rect 39 38 41 66
rect 49 38 51 66
rect 59 38 61 57
<< polycontact >>
rect 36 30 40 34
rect 50 30 54 34
<< ndcontact >>
rect 16 15 20 19
rect 16 7 20 11
rect 26 21 30 25
rect 26 14 30 18
rect 36 15 40 19
rect 36 7 40 11
<< pdcontact >>
rect 3 61 7 65
rect 3 54 7 58
rect 3 47 7 51
rect 13 46 17 50
rect 13 39 17 43
rect 23 61 27 65
rect 23 53 27 57
rect 33 46 37 50
rect 33 39 37 43
rect 43 61 47 65
rect 43 53 47 57
rect 53 46 57 50
rect 53 39 57 43
rect 63 52 67 56
rect 63 45 67 49
<< psubstratepcontact >>
rect 4 4 8 8
rect 63 4 67 8
<< nsubstratencontact >>
rect 62 64 66 68
<< psubstratepdiff >>
rect 3 8 9 24
rect 3 4 4 8
rect 8 4 9 8
rect 62 8 68 24
rect 3 3 9 4
rect 62 4 63 8
rect 67 4 68 8
rect 62 3 68 4
<< nsubstratendiff >>
rect 61 68 67 69
rect 61 64 62 68
rect 66 64 67 68
rect 61 63 67 64
<< labels >>
rlabel metal1 12 40 12 40 6 z
rlabel metal1 28 32 28 32 6 z
rlabel metal1 20 40 20 40 6 z
rlabel metal1 36 4 36 4 6 vss
rlabel metal1 44 32 44 32 6 a
rlabel metal1 52 28 52 28 6 a
rlabel metal1 44 40 44 40 6 z
rlabel metal1 52 40 52 40 6 z
rlabel metal1 36 44 36 44 6 z
rlabel metal1 36 68 36 68 6 vdd
rlabel metal1 60 40 60 40 6 z
<< end >>
