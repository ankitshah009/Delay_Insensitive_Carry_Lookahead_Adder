magic
tech scmos
timestamp 1179387182
<< checkpaint >>
rect -22 -25 86 105
<< ab >>
rect 0 0 64 80
<< pwell >>
rect -4 -7 68 36
<< nwell >>
rect -4 36 68 87
<< polysilicon >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 36 70 38 74
rect 46 60 48 65
rect 53 60 55 65
rect 9 39 11 42
rect 19 39 21 42
rect 9 38 21 39
rect 9 34 16 38
rect 20 34 21 38
rect 9 33 21 34
rect 9 30 11 33
rect 19 30 21 33
rect 29 35 31 44
rect 36 41 38 44
rect 46 41 48 44
rect 36 39 48 41
rect 53 41 55 44
rect 53 40 62 41
rect 53 39 57 40
rect 41 38 48 39
rect 29 34 37 35
rect 29 32 32 34
rect 31 30 32 32
rect 36 30 37 34
rect 31 29 37 30
rect 41 34 42 38
rect 46 34 48 38
rect 56 36 57 39
rect 61 36 62 40
rect 56 35 62 36
rect 41 33 48 34
rect 31 26 33 29
rect 41 26 43 33
rect 9 11 11 16
rect 19 11 21 16
rect 31 9 33 14
rect 41 9 43 14
<< ndiffusion >>
rect 2 21 9 30
rect 2 17 3 21
rect 7 17 9 21
rect 2 16 9 17
rect 11 29 19 30
rect 11 25 13 29
rect 17 25 19 29
rect 11 22 19 25
rect 11 18 13 22
rect 17 18 19 22
rect 11 16 19 18
rect 21 26 28 30
rect 21 16 31 26
rect 23 14 31 16
rect 33 22 41 26
rect 33 18 35 22
rect 39 18 41 22
rect 33 14 41 18
rect 43 19 51 26
rect 43 15 45 19
rect 49 15 51 19
rect 43 14 51 15
rect 23 12 29 14
rect 23 8 24 12
rect 28 8 29 12
rect 23 7 29 8
<< pdiffusion >>
rect 2 69 9 70
rect 2 65 3 69
rect 7 65 9 69
rect 2 62 9 65
rect 2 58 3 62
rect 7 58 9 62
rect 2 42 9 58
rect 11 55 19 70
rect 11 51 13 55
rect 17 51 19 55
rect 11 47 19 51
rect 11 43 13 47
rect 17 43 19 47
rect 11 42 19 43
rect 21 69 29 70
rect 21 65 23 69
rect 27 65 29 69
rect 21 62 29 65
rect 21 58 23 62
rect 27 58 29 62
rect 21 44 29 58
rect 31 44 36 70
rect 38 60 43 70
rect 38 54 46 60
rect 38 50 40 54
rect 44 50 46 54
rect 38 44 46 50
rect 48 44 53 60
rect 55 59 62 60
rect 55 55 57 59
rect 61 55 62 59
rect 55 44 62 55
rect 21 42 27 44
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect -2 69 66 78
rect -2 68 3 69
rect 2 65 3 68
rect 7 68 23 69
rect 7 65 8 68
rect 2 62 8 65
rect 2 58 3 62
rect 7 58 8 62
rect 22 65 23 68
rect 27 68 66 69
rect 27 65 28 68
rect 22 62 28 65
rect 22 58 23 62
rect 27 58 28 62
rect 57 59 61 68
rect 13 55 17 56
rect 57 54 61 55
rect 13 47 17 51
rect 2 43 13 47
rect 2 42 17 43
rect 23 50 40 54
rect 44 50 45 54
rect 2 30 6 42
rect 23 38 27 50
rect 58 46 62 47
rect 15 34 16 38
rect 20 34 27 38
rect 2 29 17 30
rect 2 25 13 29
rect 13 22 17 25
rect 2 17 3 21
rect 7 17 8 21
rect 23 22 27 34
rect 32 42 62 46
rect 32 34 36 42
rect 57 40 62 42
rect 32 29 36 30
rect 41 34 42 38
rect 46 34 47 38
rect 41 31 47 34
rect 61 36 62 40
rect 57 33 62 36
rect 41 25 54 31
rect 23 18 35 22
rect 39 18 40 22
rect 45 19 49 20
rect 13 17 17 18
rect 2 12 8 17
rect 45 12 49 15
rect -2 8 24 12
rect 28 8 66 12
rect -2 2 66 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
<< ntransistor >>
rect 9 16 11 30
rect 19 16 21 30
rect 31 14 33 26
rect 41 14 43 26
<< ptransistor >>
rect 9 42 11 70
rect 19 42 21 70
rect 29 44 31 70
rect 36 44 38 70
rect 46 44 48 60
rect 53 44 55 60
<< polycontact >>
rect 16 34 20 38
rect 32 30 36 34
rect 42 34 46 38
rect 57 36 61 40
<< ndcontact >>
rect 3 17 7 21
rect 13 25 17 29
rect 13 18 17 22
rect 35 18 39 22
rect 45 15 49 19
rect 24 8 28 12
<< pdcontact >>
rect 3 65 7 69
rect 3 58 7 62
rect 13 51 17 55
rect 13 43 17 47
rect 23 65 27 69
rect 23 58 27 62
rect 40 50 44 54
rect 57 55 61 59
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
<< psubstratepdiff >>
rect 0 2 64 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 64 2
rect 0 -3 64 -2
<< nsubstratendiff >>
rect 0 82 64 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 64 82
rect 0 77 64 78
<< labels >>
rlabel polysilicon 15 36 15 36 6 zn
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 28 12 28 6 z
rlabel metal1 12 44 12 44 6 z
rlabel metal1 32 6 32 6 6 vss
rlabel metal1 21 36 21 36 6 zn
rlabel metal1 36 44 36 44 6 a
rlabel metal1 32 74 32 74 6 vdd
rlabel metal1 31 20 31 20 6 zn
rlabel metal1 44 32 44 32 6 b
rlabel metal1 44 44 44 44 6 a
rlabel metal1 34 52 34 52 6 zn
rlabel metal1 52 28 52 28 6 b
rlabel metal1 52 44 52 44 6 a
rlabel metal1 60 40 60 40 6 a
<< end >>
