.subckt nr2av0x1 a b vdd vss z
*   SPICE3 file   created from nr2av0x1.ext -      technology: scmos
m00 vdd    vdd    w1     vdd p w=26u  l=2.3636u ad=147.333p pd=46u      as=182p     ps=66u
m01 w2     a      vdd    vdd p w=26u  l=2.3636u ad=182p     pd=66u      as=147.333p ps=46u
m02 w3     w2     vdd    vdd p w=26u  l=2.3636u ad=130p     pd=36u      as=147.333p ps=46u
m03 z      b      w3     vdd p w=26u  l=2.3636u ad=182p     pd=66u      as=130p     ps=36u
m04 vss    vss    w4     vss n w=18u  l=2.3636u ad=108p     pd=39u      as=126p     ps=50u
m05 w2     a      vss    vss n w=18u  l=2.3636u ad=126p     pd=50u      as=108p     ps=39u
m06 z      w2     vss    vss n w=18u  l=2.3636u ad=90p      pd=28u      as=108p     ps=39u
m07 vss    b      z      vss n w=18u  l=2.3636u ad=108p     pd=39u      as=90p      ps=28u
C0  w2     vdd    0.123f
C1  z      w3     0.022f
C2  z      b      0.249f
C3  vss    w2     0.191f
C4  z      a      0.033f
C5  vss    vdd    0.047f
C6  b      w2     0.181f
C7  b      vdd    0.014f
C8  w2     a      0.178f
C9  a      vdd    0.092f
C10 vss    b      0.045f
C11 z      w2     0.193f
C12 vss    a      0.102f
C13 z      vdd    0.011f
C14 b      a      0.046f
C15 vss    z      0.055f
C17 z      vss    0.006f
C18 b      vss    0.061f
C19 w2     vss    0.067f
C20 a      vss    0.062f
.ends
