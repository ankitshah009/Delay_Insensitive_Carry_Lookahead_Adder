magic
tech scmos
timestamp 1179385854
<< checkpaint >>
rect -22 -22 78 94
<< ab >>
rect 0 0 56 72
<< pwell >>
rect -4 -4 60 32
<< nwell >>
rect -4 32 60 76
<< polysilicon >>
rect 9 66 11 70
rect 19 66 21 70
rect 29 66 31 70
rect 39 58 41 63
rect 9 35 11 38
rect 19 35 21 38
rect 29 35 31 38
rect 39 35 41 38
rect 9 34 41 35
rect 9 33 27 34
rect 9 26 11 33
rect 19 26 21 33
rect 26 30 27 33
rect 31 30 36 34
rect 40 30 41 34
rect 26 29 41 30
rect 29 26 31 29
rect 39 26 41 29
rect 9 11 11 16
rect 19 7 21 12
rect 29 7 31 12
rect 39 7 41 12
<< ndiffusion >>
rect 2 21 9 26
rect 2 17 3 21
rect 7 17 9 21
rect 2 16 9 17
rect 11 25 19 26
rect 11 21 13 25
rect 17 21 19 25
rect 11 16 19 21
rect 14 12 19 16
rect 21 17 29 26
rect 21 13 23 17
rect 27 13 29 17
rect 21 12 29 13
rect 31 25 39 26
rect 31 21 33 25
rect 37 21 39 25
rect 31 18 39 21
rect 31 14 33 18
rect 37 14 39 18
rect 31 12 39 14
rect 41 25 48 26
rect 41 21 43 25
rect 47 21 48 25
rect 41 17 48 21
rect 41 13 43 17
rect 47 13 48 17
rect 41 12 48 13
<< pdiffusion >>
rect 2 65 9 66
rect 2 61 3 65
rect 7 61 9 65
rect 2 58 9 61
rect 2 54 3 58
rect 7 54 9 58
rect 2 38 9 54
rect 11 50 19 66
rect 11 46 13 50
rect 17 46 19 50
rect 11 43 19 46
rect 11 39 13 43
rect 17 39 19 43
rect 11 38 19 39
rect 21 65 29 66
rect 21 61 23 65
rect 27 61 29 65
rect 21 57 29 61
rect 21 53 23 57
rect 27 53 29 57
rect 21 38 29 53
rect 31 58 36 66
rect 31 50 39 58
rect 31 46 33 50
rect 37 46 39 50
rect 31 43 39 46
rect 31 39 33 43
rect 37 39 39 43
rect 31 38 39 39
rect 41 57 48 58
rect 41 53 43 57
rect 47 53 48 57
rect 41 50 48 53
rect 41 46 43 50
rect 47 46 48 50
rect 41 38 48 46
<< metal1 >>
rect -2 68 58 72
rect -2 65 48 68
rect -2 64 3 65
rect 2 61 3 64
rect 7 64 23 65
rect 7 61 8 64
rect 2 58 8 61
rect 2 54 3 58
rect 7 54 8 58
rect 27 64 48 65
rect 52 64 58 68
rect 23 57 27 61
rect 23 52 27 53
rect 42 57 48 64
rect 42 53 43 57
rect 47 53 48 57
rect 13 50 17 51
rect 13 43 17 46
rect 10 39 13 43
rect 33 50 38 51
rect 37 46 38 50
rect 42 50 48 53
rect 42 46 43 50
rect 47 46 48 50
rect 33 43 38 46
rect 17 39 33 42
rect 37 39 38 43
rect 10 38 38 39
rect 10 26 14 38
rect 42 34 47 43
rect 25 30 27 34
rect 31 30 36 34
rect 40 30 47 34
rect 10 25 38 26
rect 3 21 7 22
rect 10 21 13 25
rect 17 22 33 25
rect 17 21 18 22
rect 37 21 38 25
rect 33 18 38 21
rect 3 8 7 17
rect 23 17 27 18
rect 37 14 38 18
rect 33 13 38 14
rect 43 25 47 26
rect 43 17 47 21
rect 23 8 27 13
rect 43 8 47 13
rect -2 4 4 8
rect 8 4 58 8
rect -2 0 58 4
<< ntransistor >>
rect 9 16 11 26
rect 19 12 21 26
rect 29 12 31 26
rect 39 12 41 26
<< ptransistor >>
rect 9 38 11 66
rect 19 38 21 66
rect 29 38 31 66
rect 39 38 41 58
<< polycontact >>
rect 27 30 31 34
rect 36 30 40 34
<< ndcontact >>
rect 3 17 7 21
rect 13 21 17 25
rect 23 13 27 17
rect 33 21 37 25
rect 33 14 37 18
rect 43 21 47 25
rect 43 13 47 17
<< pdcontact >>
rect 3 61 7 65
rect 3 54 7 58
rect 13 46 17 50
rect 13 39 17 43
rect 23 61 27 65
rect 23 53 27 57
rect 33 46 37 50
rect 33 39 37 43
rect 43 53 47 57
rect 43 46 47 50
<< psubstratepcontact >>
rect 4 4 8 8
<< nsubstratencontact >>
rect 48 64 52 68
<< psubstratepdiff >>
rect 3 8 9 9
rect 3 4 4 8
rect 8 4 9 8
rect 3 3 9 4
<< nsubstratendiff >>
rect 47 68 53 69
rect 47 64 48 68
rect 52 64 53 68
rect 47 63 53 64
<< labels >>
rlabel metal1 12 32 12 32 6 z
rlabel metal1 20 24 20 24 6 z
rlabel metal1 20 40 20 40 6 z
rlabel metal1 28 4 28 4 6 vss
rlabel ndcontact 36 16 36 16 6 z
rlabel metal1 28 24 28 24 6 z
rlabel polycontact 28 32 28 32 6 a
rlabel metal1 36 32 36 32 6 a
rlabel metal1 28 40 28 40 6 z
rlabel pdcontact 36 48 36 48 6 z
rlabel metal1 28 68 28 68 6 vdd
rlabel metal1 44 36 44 36 6 a
<< end >>
