magic
tech scmos
timestamp 1179387181
<< checkpaint >>
rect -22 -22 86 94
<< ab >>
rect 0 0 64 72
<< pwell >>
rect -4 -4 68 32
<< nwell >>
rect -4 32 68 76
<< polysilicon >>
rect 9 66 11 70
rect 19 66 21 70
rect 29 66 31 70
rect 36 66 38 70
rect 46 56 48 61
rect 53 56 55 61
rect 9 35 11 38
rect 19 35 21 38
rect 9 34 21 35
rect 9 30 16 34
rect 20 30 21 34
rect 9 29 21 30
rect 9 26 11 29
rect 19 26 21 29
rect 29 31 31 40
rect 36 37 38 40
rect 46 37 48 40
rect 36 35 48 37
rect 53 37 55 40
rect 53 36 62 37
rect 53 35 57 36
rect 41 34 48 35
rect 29 30 37 31
rect 29 28 32 30
rect 31 26 32 28
rect 36 26 37 30
rect 31 25 37 26
rect 41 30 42 34
rect 46 30 48 34
rect 56 32 57 35
rect 61 32 62 36
rect 56 31 62 32
rect 41 29 48 30
rect 31 22 33 25
rect 41 22 43 29
rect 9 7 11 12
rect 19 7 21 12
rect 31 5 33 10
rect 41 5 43 10
<< ndiffusion >>
rect 2 17 9 26
rect 2 13 3 17
rect 7 13 9 17
rect 2 12 9 13
rect 11 25 19 26
rect 11 21 13 25
rect 17 21 19 25
rect 11 18 19 21
rect 11 14 13 18
rect 17 14 19 18
rect 11 12 19 14
rect 21 22 28 26
rect 21 12 31 22
rect 23 10 31 12
rect 33 18 41 22
rect 33 14 35 18
rect 39 14 41 18
rect 33 10 41 14
rect 43 15 51 22
rect 43 11 45 15
rect 49 11 51 15
rect 43 10 51 11
rect 23 8 29 10
rect 23 4 24 8
rect 28 4 29 8
rect 23 3 29 4
<< pdiffusion >>
rect 2 65 9 66
rect 2 61 3 65
rect 7 61 9 65
rect 2 58 9 61
rect 2 54 3 58
rect 7 54 9 58
rect 2 38 9 54
rect 11 51 19 66
rect 11 47 13 51
rect 17 47 19 51
rect 11 43 19 47
rect 11 39 13 43
rect 17 39 19 43
rect 11 38 19 39
rect 21 65 29 66
rect 21 61 23 65
rect 27 61 29 65
rect 21 58 29 61
rect 21 54 23 58
rect 27 54 29 58
rect 21 40 29 54
rect 31 40 36 66
rect 38 56 43 66
rect 38 50 46 56
rect 38 46 40 50
rect 44 46 46 50
rect 38 40 46 46
rect 48 40 53 56
rect 55 55 62 56
rect 55 51 57 55
rect 61 51 62 55
rect 55 40 62 51
rect 21 38 27 40
<< metal1 >>
rect -2 68 66 72
rect -2 65 48 68
rect -2 64 3 65
rect 2 61 3 64
rect 7 64 23 65
rect 7 61 8 64
rect 2 58 8 61
rect 2 54 3 58
rect 7 54 8 58
rect 22 61 23 64
rect 27 64 48 65
rect 52 64 56 68
rect 60 64 66 68
rect 27 61 28 64
rect 22 58 28 61
rect 22 54 23 58
rect 27 54 28 58
rect 57 55 61 64
rect 13 51 17 52
rect 57 50 61 51
rect 13 43 17 47
rect 2 39 13 43
rect 2 38 17 39
rect 23 46 40 50
rect 44 46 45 50
rect 2 26 6 38
rect 23 34 27 46
rect 58 42 62 43
rect 15 30 16 34
rect 20 30 27 34
rect 2 25 17 26
rect 2 21 13 25
rect 13 18 17 21
rect 2 13 3 17
rect 7 13 8 17
rect 23 18 27 30
rect 32 38 62 42
rect 32 30 36 38
rect 57 36 62 38
rect 32 25 36 26
rect 41 30 42 34
rect 46 30 47 34
rect 41 27 47 30
rect 61 32 62 36
rect 57 29 62 32
rect 41 21 54 27
rect 23 14 35 18
rect 39 14 40 18
rect 45 15 49 16
rect 13 13 17 14
rect 2 8 8 13
rect 45 8 49 11
rect -2 4 24 8
rect 28 4 56 8
rect 60 4 66 8
rect -2 0 66 4
<< ntransistor >>
rect 9 12 11 26
rect 19 12 21 26
rect 31 10 33 22
rect 41 10 43 22
<< ptransistor >>
rect 9 38 11 66
rect 19 38 21 66
rect 29 40 31 66
rect 36 40 38 66
rect 46 40 48 56
rect 53 40 55 56
<< polycontact >>
rect 16 30 20 34
rect 32 26 36 30
rect 42 30 46 34
rect 57 32 61 36
<< ndcontact >>
rect 3 13 7 17
rect 13 21 17 25
rect 13 14 17 18
rect 35 14 39 18
rect 45 11 49 15
rect 24 4 28 8
<< pdcontact >>
rect 3 61 7 65
rect 3 54 7 58
rect 13 47 17 51
rect 13 39 17 43
rect 23 61 27 65
rect 23 54 27 58
rect 40 46 44 50
rect 57 51 61 55
<< psubstratepcontact >>
rect 56 4 60 8
<< nsubstratencontact >>
rect 48 64 52 68
rect 56 64 60 68
<< psubstratepdiff >>
rect 55 8 61 24
rect 55 4 56 8
rect 60 4 61 8
rect 55 3 61 4
<< nsubstratendiff >>
rect 47 68 61 69
rect 47 64 48 68
rect 52 64 56 68
rect 60 64 61 68
rect 47 63 61 64
<< labels >>
rlabel polysilicon 15 32 15 32 6 zn
rlabel metal1 4 32 4 32 6 z
rlabel metal1 12 24 12 24 6 z
rlabel metal1 12 40 12 40 6 z
rlabel metal1 21 32 21 32 6 zn
rlabel metal1 32 4 32 4 6 vss
rlabel metal1 31 16 31 16 6 zn
rlabel metal1 44 28 44 28 6 b
rlabel metal1 44 40 44 40 6 a
rlabel metal1 36 40 36 40 6 a
rlabel metal1 34 48 34 48 6 zn
rlabel metal1 32 68 32 68 6 vdd
rlabel metal1 52 24 52 24 6 b
rlabel metal1 60 36 60 36 6 a
rlabel metal1 52 40 52 40 6 a
<< end >>
