magic
tech scmos
timestamp 1179385656
<< checkpaint >>
rect -22 -25 94 105
<< ab >>
rect 0 0 72 80
<< pwell >>
rect -4 -7 76 36
<< nwell >>
rect -4 36 76 87
<< polysilicon >>
rect 26 67 48 69
rect 9 58 11 63
rect 19 58 21 63
rect 26 58 28 67
rect 36 58 38 63
rect 46 58 48 67
rect 58 62 60 67
rect 9 37 11 42
rect 19 37 21 42
rect 9 35 21 37
rect 9 32 11 35
rect 5 31 11 32
rect 5 27 6 31
rect 10 27 11 31
rect 19 30 21 35
rect 26 30 28 42
rect 36 39 38 42
rect 32 38 38 39
rect 32 34 33 38
rect 37 34 38 38
rect 32 33 38 34
rect 36 30 38 33
rect 46 39 48 42
rect 58 39 60 42
rect 46 38 53 39
rect 46 34 48 38
rect 52 34 53 38
rect 46 33 53 34
rect 57 38 63 39
rect 57 34 58 38
rect 62 34 63 38
rect 57 33 63 34
rect 46 30 48 33
rect 58 30 60 33
rect 5 26 11 27
rect 9 23 11 26
rect 19 18 21 23
rect 26 18 28 23
rect 36 18 38 23
rect 46 18 48 23
rect 9 11 11 16
rect 58 15 60 20
<< ndiffusion >>
rect 13 23 19 30
rect 21 23 26 30
rect 28 29 36 30
rect 28 25 30 29
rect 34 25 36 29
rect 28 23 36 25
rect 38 28 46 30
rect 38 24 40 28
rect 44 24 46 28
rect 38 23 46 24
rect 48 23 58 30
rect 2 21 9 23
rect 2 17 3 21
rect 7 17 9 21
rect 2 16 9 17
rect 11 16 17 23
rect 50 20 58 23
rect 60 29 67 30
rect 60 25 62 29
rect 66 25 67 29
rect 60 24 67 25
rect 60 20 65 24
rect 50 16 51 20
rect 55 16 56 20
rect 13 12 19 16
rect 50 15 56 16
rect 13 8 14 12
rect 18 8 19 12
rect 13 7 19 8
<< pdiffusion >>
rect 13 72 19 73
rect 13 68 14 72
rect 18 68 19 72
rect 13 65 19 68
rect 13 58 17 65
rect 50 61 58 62
rect 50 58 51 61
rect 2 57 9 58
rect 2 53 3 57
rect 7 53 9 57
rect 2 50 9 53
rect 2 46 3 50
rect 7 46 9 50
rect 2 45 9 46
rect 4 42 9 45
rect 11 42 19 58
rect 21 42 26 58
rect 28 55 36 58
rect 28 51 30 55
rect 34 51 36 55
rect 28 42 36 51
rect 38 57 46 58
rect 38 53 40 57
rect 44 53 46 57
rect 38 50 46 53
rect 38 46 40 50
rect 44 46 46 50
rect 38 42 46 46
rect 48 57 51 58
rect 55 57 58 61
rect 48 42 58 57
rect 60 61 67 62
rect 60 57 62 61
rect 66 57 67 61
rect 60 54 67 57
rect 60 50 62 54
rect 66 50 67 54
rect 60 49 67 50
rect 60 42 65 49
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect -2 72 74 78
rect -2 68 14 72
rect 18 68 74 72
rect 3 59 44 63
rect 3 57 7 59
rect 40 57 44 59
rect 50 61 56 68
rect 50 57 51 61
rect 55 57 56 61
rect 62 61 66 62
rect 3 50 7 53
rect 10 51 30 55
rect 34 51 35 55
rect 62 54 66 57
rect 10 49 22 51
rect 3 45 7 46
rect 2 27 6 39
rect 10 27 14 31
rect 2 25 14 27
rect 18 30 22 49
rect 40 50 44 53
rect 26 38 30 47
rect 40 45 44 46
rect 49 46 55 54
rect 66 50 70 53
rect 62 49 70 50
rect 49 42 63 46
rect 48 38 52 39
rect 26 34 33 38
rect 37 34 39 38
rect 57 38 63 42
rect 57 34 58 38
rect 62 34 63 38
rect 18 29 35 30
rect 48 29 52 34
rect 18 25 30 29
rect 34 25 35 29
rect 40 28 44 29
rect 48 25 62 29
rect 66 25 70 49
rect 40 21 44 24
rect 2 17 3 21
rect 7 17 44 21
rect 51 20 55 21
rect 51 12 55 16
rect -2 8 14 12
rect 18 8 74 12
rect -2 2 74 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
<< ntransistor >>
rect 19 23 21 30
rect 26 23 28 30
rect 36 23 38 30
rect 46 23 48 30
rect 9 16 11 23
rect 58 20 60 30
<< ptransistor >>
rect 9 42 11 58
rect 19 42 21 58
rect 26 42 28 58
rect 36 42 38 58
rect 46 42 48 58
rect 58 42 60 62
<< polycontact >>
rect 6 27 10 31
rect 33 34 37 38
rect 48 34 52 38
rect 58 34 62 38
<< ndcontact >>
rect 30 25 34 29
rect 40 24 44 28
rect 3 17 7 21
rect 62 25 66 29
rect 51 16 55 20
rect 14 8 18 12
<< pdcontact >>
rect 14 68 18 72
rect 3 53 7 57
rect 3 46 7 50
rect 30 51 34 55
rect 40 53 44 57
rect 40 46 44 50
rect 51 57 55 61
rect 62 57 66 61
rect 62 50 66 54
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
<< psubstratepdiff >>
rect 0 2 72 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 72 2
rect 0 -3 72 -2
<< nsubstratendiff >>
rect 0 82 72 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 72 82
rect 0 77 72 78
<< labels >>
rlabel polycontact 49 36 49 36 6 bn
rlabel metal1 4 32 4 32 6 a
rlabel pdcontact 5 54 5 54 6 n1
rlabel metal1 12 28 12 28 6 a
rlabel metal1 20 40 20 40 6 z
rlabel metal1 12 52 12 52 6 z
rlabel metal1 36 6 36 6 6 vss
rlabel metal1 28 28 28 28 6 z
rlabel metal1 28 44 28 44 6 c
rlabel polycontact 36 36 36 36 6 c
rlabel metal1 36 74 36 74 6 vdd
rlabel metal1 42 23 42 23 6 n3
rlabel metal1 23 19 23 19 6 n3
rlabel metal1 50 32 50 32 6 bn
rlabel metal1 52 48 52 48 6 b
rlabel pdcontact 42 54 42 54 6 n1
rlabel metal1 59 27 59 27 6 bn
rlabel metal1 60 40 60 40 6 b
rlabel metal1 64 55 64 55 6 bn
<< end >>
