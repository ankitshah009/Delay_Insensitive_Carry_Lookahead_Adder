magic
tech scmos
timestamp 1179387350
<< checkpaint >>
rect -22 -25 38 105
<< ab >>
rect 0 0 16 80
<< pwell >>
rect -4 -7 20 36
<< nwell >>
rect -4 36 20 87
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect -2 68 18 78
rect -2 2 18 12
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
<< psubstratepdiff >>
rect 0 2 16 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 16 2
rect 0 -3 16 -2
<< nsubstratendiff >>
rect 0 82 16 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 16 82
rect 0 77 16 78
<< labels >>
rlabel metal1 8 6 8 6 6 vss
rlabel metal1 8 74 8 74 6 vdd
<< end >>
