magic
tech scmos
timestamp 1179387410
<< checkpaint >>
rect -22 -22 102 94
<< ab >>
rect 0 0 80 72
<< pwell >>
rect -4 -4 84 32
<< nwell >>
rect -4 32 84 76
<< polysilicon >>
rect 9 66 11 70
rect 27 66 29 70
rect 37 66 39 70
rect 44 66 46 70
rect 57 66 59 70
rect 67 66 69 70
rect 9 35 11 38
rect 27 35 29 38
rect 9 34 29 35
rect 9 30 10 34
rect 14 33 29 34
rect 14 30 15 33
rect 37 31 39 38
rect 44 35 46 38
rect 57 35 59 38
rect 9 29 15 30
rect 33 30 39 31
rect 11 22 13 29
rect 33 27 34 30
rect 21 26 34 27
rect 38 26 39 30
rect 43 34 49 35
rect 43 30 44 34
rect 48 31 49 34
rect 57 34 63 35
rect 48 30 52 31
rect 43 29 52 30
rect 57 30 58 34
rect 62 30 63 34
rect 57 29 63 30
rect 67 32 69 38
rect 67 31 73 32
rect 21 25 39 26
rect 21 22 23 25
rect 50 23 52 29
rect 60 23 62 29
rect 67 27 68 31
rect 72 27 73 31
rect 67 26 73 27
rect 67 23 69 26
rect 11 4 13 9
rect 21 4 23 9
rect 50 2 52 6
rect 60 2 62 6
rect 67 2 69 6
<< ndiffusion >>
rect 4 14 11 22
rect 4 10 5 14
rect 9 10 11 14
rect 4 9 11 10
rect 13 21 21 22
rect 13 17 15 21
rect 19 17 21 21
rect 13 9 21 17
rect 23 21 31 22
rect 23 17 26 21
rect 30 17 31 21
rect 45 19 50 23
rect 23 16 31 17
rect 42 18 50 19
rect 23 9 28 16
rect 42 14 43 18
rect 47 14 50 18
rect 42 13 50 14
rect 45 6 50 13
rect 52 22 60 23
rect 52 18 54 22
rect 58 18 60 22
rect 52 6 60 18
rect 62 6 67 23
rect 69 11 76 23
rect 69 7 71 11
rect 75 7 76 11
rect 69 6 76 7
<< pdiffusion >>
rect 2 65 9 66
rect 2 61 3 65
rect 7 61 9 65
rect 2 58 9 61
rect 2 54 3 58
rect 7 54 9 58
rect 2 38 9 54
rect 11 44 16 66
rect 22 59 27 66
rect 20 58 27 59
rect 20 54 21 58
rect 25 54 27 58
rect 20 53 27 54
rect 11 43 18 44
rect 11 39 13 43
rect 17 39 18 43
rect 11 38 18 39
rect 22 38 27 53
rect 29 43 37 66
rect 29 39 31 43
rect 35 39 37 43
rect 29 38 37 39
rect 39 38 44 66
rect 46 65 57 66
rect 46 61 49 65
rect 53 61 57 65
rect 46 38 57 61
rect 59 58 67 66
rect 59 54 61 58
rect 65 54 67 58
rect 59 51 67 54
rect 59 47 61 51
rect 65 47 67 51
rect 59 38 67 47
rect 69 65 77 66
rect 69 61 71 65
rect 75 61 77 65
rect 69 58 77 61
rect 69 54 71 58
rect 75 54 77 58
rect 69 38 77 54
<< metal1 >>
rect -2 65 82 72
rect -2 64 3 65
rect 2 61 3 64
rect 7 64 49 65
rect 7 61 8 64
rect 48 61 49 64
rect 53 64 71 65
rect 53 61 54 64
rect 70 61 71 64
rect 75 64 82 65
rect 75 61 76 64
rect 2 58 8 61
rect 61 58 66 59
rect 2 54 3 58
rect 7 54 8 58
rect 20 54 21 58
rect 25 54 55 58
rect 51 51 55 54
rect 65 54 66 58
rect 70 58 76 61
rect 70 54 71 58
rect 75 54 76 58
rect 61 51 66 54
rect 18 46 46 50
rect 18 43 22 46
rect 2 35 6 43
rect 12 39 13 43
rect 17 39 22 43
rect 2 34 14 35
rect 2 30 10 34
rect 2 29 14 30
rect 2 21 6 29
rect 18 21 22 39
rect 14 17 15 21
rect 19 17 22 21
rect 26 39 31 43
rect 35 39 36 43
rect 26 21 30 39
rect 42 35 46 46
rect 51 47 61 51
rect 65 47 66 51
rect 42 34 48 35
rect 34 30 38 31
rect 42 30 44 34
rect 42 29 48 30
rect 51 26 55 47
rect 58 37 78 43
rect 58 34 62 37
rect 58 29 62 30
rect 68 31 72 32
rect 34 22 55 26
rect 66 25 78 27
rect 51 18 54 22
rect 58 18 59 22
rect 65 21 78 25
rect 30 17 43 18
rect 5 14 9 15
rect 26 14 43 17
rect 47 14 48 18
rect 65 14 71 21
rect 5 8 9 10
rect 70 8 71 11
rect -2 4 33 8
rect 37 7 71 8
rect 75 8 76 11
rect 75 7 82 8
rect 37 4 82 7
rect -2 0 82 4
<< ntransistor >>
rect 11 9 13 22
rect 21 9 23 22
rect 50 6 52 23
rect 60 6 62 23
rect 67 6 69 23
<< ptransistor >>
rect 9 38 11 66
rect 27 38 29 66
rect 37 38 39 66
rect 44 38 46 66
rect 57 38 59 66
rect 67 38 69 66
<< polycontact >>
rect 10 30 14 34
rect 34 26 38 30
rect 44 30 48 34
rect 58 30 62 34
rect 68 27 72 31
<< ndcontact >>
rect 5 10 9 14
rect 15 17 19 21
rect 26 17 30 21
rect 43 14 47 18
rect 54 18 58 22
rect 71 7 75 11
<< pdcontact >>
rect 3 61 7 65
rect 3 54 7 58
rect 21 54 25 58
rect 13 39 17 43
rect 31 39 35 43
rect 49 61 53 65
rect 61 54 65 58
rect 61 47 65 51
rect 71 61 75 65
rect 71 54 75 58
<< psubstratepcontact >>
rect 33 4 37 8
<< psubstratepdiff >>
rect 32 8 38 9
rect 32 4 33 8
rect 37 4 38 8
rect 32 3 38 4
<< labels >>
rlabel polycontact 36 28 36 28 6 an
rlabel ptransistor 45 49 45 49 6 bn
rlabel metal1 4 32 4 32 6 b
rlabel polycontact 12 32 12 32 6 b
rlabel metal1 36 16 36 16 6 z
rlabel metal1 36 26 36 26 6 an
rlabel metal1 28 32 28 32 6 z
rlabel metal1 20 33 20 33 6 bn
rlabel metal1 17 41 17 41 6 bn
rlabel metal1 40 4 40 4 6 vss
rlabel ndcontact 44 16 44 16 6 z
rlabel metal1 44 39 44 39 6 bn
rlabel metal1 37 56 37 56 6 an
rlabel metal1 53 38 53 38 6 an
rlabel metal1 40 68 40 68 6 vdd
rlabel metal1 68 20 68 20 6 a1
rlabel metal1 76 24 76 24 6 a1
rlabel metal1 68 40 68 40 6 a2
rlabel metal1 76 40 76 40 6 a2
rlabel metal1 60 36 60 36 6 a2
rlabel metal1 63 53 63 53 6 an
<< end >>
