.subckt nd2v3x4 a b vdd vss z
*   SPICE3 file   created from nd2v3x4.ext -      technology: scmos
m00 z      a      vdd    vdd p w=24u  l=2.3636u ad=96p      pd=32u      as=138p     ps=47.5u
m01 vdd    b      z      vdd p w=24u  l=2.3636u ad=138p     pd=47.5u    as=96p      ps=32u
m02 z      b      vdd    vdd p w=24u  l=2.3636u ad=96p      pd=32u      as=138p     ps=47.5u
m03 vdd    a      z      vdd p w=24u  l=2.3636u ad=138p     pd=47.5u    as=96p      ps=32u
m04 w1     a      vss    vss n w=20u  l=2.3636u ad=50p      pd=25u      as=135p     ps=43.5u
m05 z      b      w1     vss n w=20u  l=2.3636u ad=80p      pd=28u      as=50p      ps=25u
m06 w2     b      z      vss n w=20u  l=2.3636u ad=50p      pd=25u      as=80p      ps=28u
m07 vss    a      w2     vss n w=20u  l=2.3636u ad=135p     pd=43.5u    as=50p      ps=25u
m08 w3     a      vss    vss n w=20u  l=2.3636u ad=50p      pd=25u      as=135p     ps=43.5u
m09 z      b      w3     vss n w=20u  l=2.3636u ad=80p      pd=28u      as=50p      ps=25u
m10 w4     b      z      vss n w=20u  l=2.3636u ad=50p      pd=25u      as=80p      ps=28u
m11 vss    a      w4     vss n w=20u  l=2.3636u ad=135p     pd=43.5u    as=50p      ps=25u
C0  vss    z      0.472f
C1  w2     a      0.007f
C2  vss    a      0.218f
C3  z      b      0.225f
C4  z      vdd    0.294f
C5  b      a      0.542f
C6  w4     vss    0.005f
C7  a      vdd    0.070f
C8  w2     vss    0.005f
C9  w3     z      0.010f
C10 w1     z      0.010f
C11 w3     a      0.007f
C12 w1     a      0.007f
C13 vss    b      0.058f
C14 vss    vdd    0.003f
C15 z      a      0.606f
C16 b      vdd    0.094f
C17 w3     vss    0.005f
C18 w2     z      0.010f
C19 w1     vss    0.005f
C20 w4     a      0.007f
C22 z      vss    0.007f
C23 b      vss    0.054f
C24 a      vss    0.052f
.ends
