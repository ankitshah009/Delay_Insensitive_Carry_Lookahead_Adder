magic
tech scmos
timestamp 1182409234
<< checkpaint >>
rect -22 -22 222 94
<< ab >>
rect 0 0 200 72
<< pwell >>
rect -4 -4 204 32
<< nwell >>
rect -4 32 204 76
<< polysilicon >>
rect 9 66 11 70
rect 19 66 21 70
rect 29 66 31 70
rect 39 66 41 70
rect 49 66 51 70
rect 59 66 61 70
rect 69 66 71 70
rect 79 66 81 70
rect 89 66 91 70
rect 99 66 101 70
rect 109 66 111 70
rect 119 66 121 70
rect 126 66 128 70
rect 136 66 138 70
rect 143 66 145 70
rect 153 66 155 70
rect 160 66 162 70
rect 170 66 172 70
rect 177 66 179 70
rect 79 43 81 46
rect 89 43 91 46
rect 99 43 101 46
rect 79 42 101 43
rect 79 38 80 42
rect 84 41 101 42
rect 84 38 85 41
rect 9 35 11 38
rect 19 35 21 38
rect 29 35 31 38
rect 9 34 31 35
rect 9 33 20 34
rect 9 26 11 33
rect 19 30 20 33
rect 24 33 31 34
rect 39 35 41 38
rect 49 35 51 38
rect 59 35 61 38
rect 69 35 71 38
rect 79 37 85 38
rect 99 39 101 41
rect 109 39 111 42
rect 99 37 111 39
rect 79 35 81 37
rect 39 34 64 35
rect 39 33 59 34
rect 24 30 25 33
rect 19 29 25 30
rect 58 30 59 33
rect 63 30 64 34
rect 58 29 64 30
rect 19 26 21 29
rect 42 25 44 29
rect 52 25 54 29
rect 62 25 64 29
rect 69 33 81 35
rect 69 25 71 33
rect 79 25 81 33
rect 89 35 95 36
rect 89 32 90 35
rect 86 31 90 32
rect 94 31 95 35
rect 119 33 121 38
rect 126 35 128 38
rect 136 35 138 38
rect 126 34 138 35
rect 126 33 130 34
rect 86 30 95 31
rect 114 32 121 33
rect 86 25 88 30
rect 114 28 115 32
rect 119 28 121 32
rect 129 30 130 33
rect 134 33 138 34
rect 143 35 145 38
rect 153 35 155 38
rect 143 34 155 35
rect 134 30 135 33
rect 129 29 135 30
rect 114 27 121 28
rect 9 6 11 9
rect 19 6 21 9
rect 42 6 44 9
rect 52 6 54 9
rect 9 4 54 6
rect 62 4 64 9
rect 69 4 71 9
rect 79 4 81 9
rect 86 4 88 9
rect 133 23 135 29
rect 143 30 146 34
rect 150 30 155 34
rect 143 29 155 30
rect 160 35 162 38
rect 170 35 172 38
rect 160 34 172 35
rect 160 30 162 34
rect 166 33 172 34
rect 166 30 167 33
rect 160 29 167 30
rect 143 23 145 29
rect 153 23 155 29
rect 163 23 165 29
rect 177 27 179 38
rect 177 26 183 27
rect 177 22 178 26
rect 182 22 183 26
rect 177 21 183 22
rect 133 2 135 6
rect 143 2 145 6
rect 153 2 155 6
rect 163 2 165 6
<< ndiffusion >>
rect 2 22 9 26
rect 2 18 3 22
rect 7 18 9 22
rect 2 14 9 18
rect 2 10 3 14
rect 7 10 9 14
rect 2 9 9 10
rect 11 25 19 26
rect 11 21 13 25
rect 17 21 19 25
rect 11 18 19 21
rect 11 14 13 18
rect 17 14 19 18
rect 11 9 19 14
rect 21 14 29 26
rect 21 10 23 14
rect 27 10 29 14
rect 35 24 42 25
rect 35 20 36 24
rect 40 20 42 24
rect 35 17 42 20
rect 35 13 36 17
rect 40 13 42 17
rect 35 12 42 13
rect 21 9 29 10
rect 37 9 42 12
rect 44 24 52 25
rect 44 20 46 24
rect 50 20 52 24
rect 44 9 52 20
rect 54 24 62 25
rect 54 20 56 24
rect 60 20 62 24
rect 54 17 62 20
rect 54 13 56 17
rect 60 13 62 17
rect 54 9 62 13
rect 64 9 69 25
rect 71 14 79 25
rect 71 10 73 14
rect 77 10 79 14
rect 71 9 79 10
rect 81 9 86 25
rect 88 24 95 25
rect 88 20 90 24
rect 94 20 95 24
rect 88 17 95 20
rect 88 13 90 17
rect 94 13 95 17
rect 88 12 95 13
rect 88 9 93 12
rect 124 18 133 23
rect 124 14 126 18
rect 130 14 133 18
rect 124 11 133 14
rect 124 7 126 11
rect 130 7 133 11
rect 124 6 133 7
rect 135 18 143 23
rect 135 14 137 18
rect 141 14 143 18
rect 135 6 143 14
rect 145 11 153 23
rect 145 7 147 11
rect 151 7 153 11
rect 145 6 153 7
rect 155 18 163 23
rect 155 14 157 18
rect 161 14 163 18
rect 155 6 163 14
rect 165 11 173 23
rect 165 7 167 11
rect 171 7 173 11
rect 165 6 173 7
<< pdiffusion >>
rect 2 65 9 66
rect 2 61 3 65
rect 7 61 9 65
rect 2 58 9 61
rect 2 54 3 58
rect 7 54 9 58
rect 2 38 9 54
rect 11 51 19 66
rect 11 47 13 51
rect 17 47 19 51
rect 11 44 19 47
rect 11 40 13 44
rect 17 40 19 44
rect 11 38 19 40
rect 21 65 29 66
rect 21 61 23 65
rect 27 61 29 65
rect 21 58 29 61
rect 21 54 23 58
rect 27 54 29 58
rect 21 38 29 54
rect 31 58 39 66
rect 31 54 33 58
rect 37 54 39 58
rect 31 51 39 54
rect 31 47 33 51
rect 37 47 39 51
rect 31 38 39 47
rect 41 59 49 66
rect 41 55 43 59
rect 47 55 49 59
rect 41 43 49 55
rect 41 39 43 43
rect 47 39 49 43
rect 41 38 49 39
rect 51 50 59 66
rect 51 46 53 50
rect 57 46 59 50
rect 51 43 59 46
rect 51 39 53 43
rect 57 39 59 43
rect 51 38 59 39
rect 61 59 69 66
rect 61 55 63 59
rect 67 55 69 59
rect 61 52 69 55
rect 61 48 63 52
rect 67 48 69 52
rect 61 38 69 48
rect 71 51 79 66
rect 71 47 73 51
rect 77 47 79 51
rect 71 46 79 47
rect 81 59 89 66
rect 81 55 83 59
rect 87 55 89 59
rect 81 46 89 55
rect 91 51 99 66
rect 91 47 93 51
rect 97 47 99 51
rect 91 46 99 47
rect 101 59 109 66
rect 101 55 103 59
rect 107 55 109 59
rect 101 46 109 55
rect 71 38 76 46
rect 104 42 109 46
rect 111 58 119 66
rect 111 54 113 58
rect 117 54 119 58
rect 111 51 119 54
rect 111 47 113 51
rect 117 47 119 51
rect 111 42 119 47
rect 114 38 119 42
rect 121 38 126 66
rect 128 65 136 66
rect 128 61 130 65
rect 134 61 136 65
rect 128 58 136 61
rect 128 54 130 58
rect 134 54 136 58
rect 128 38 136 54
rect 138 38 143 66
rect 145 58 153 66
rect 145 54 147 58
rect 151 54 153 58
rect 145 51 153 54
rect 145 47 147 51
rect 151 47 153 51
rect 145 38 153 47
rect 155 38 160 66
rect 162 65 170 66
rect 162 61 164 65
rect 168 61 170 65
rect 162 58 170 61
rect 162 54 164 58
rect 168 54 170 58
rect 162 38 170 54
rect 172 38 177 66
rect 179 51 184 66
rect 179 50 186 51
rect 179 46 181 50
rect 185 46 186 50
rect 179 43 186 46
rect 179 39 181 43
rect 185 39 186 43
rect 179 38 186 39
<< metal1 >>
rect -2 68 202 72
rect -2 65 189 68
rect -2 64 3 65
rect 2 61 3 64
rect 7 64 23 65
rect 7 61 8 64
rect 2 58 8 61
rect 2 54 3 58
rect 7 54 8 58
rect 22 61 23 64
rect 27 64 130 65
rect 27 61 28 64
rect 22 58 28 61
rect 129 61 130 64
rect 134 64 164 65
rect 134 61 135 64
rect 22 54 23 58
rect 27 54 28 58
rect 33 58 37 59
rect 42 55 43 59
rect 47 55 63 59
rect 67 55 83 59
rect 87 55 103 59
rect 107 55 108 59
rect 113 58 117 59
rect 33 51 37 54
rect 63 52 67 55
rect 12 47 13 51
rect 17 47 33 51
rect 37 50 57 51
rect 37 47 53 50
rect 12 44 17 47
rect 12 43 13 44
rect 10 40 13 43
rect 129 58 135 61
rect 163 61 164 64
rect 168 64 189 65
rect 193 64 202 68
rect 168 61 169 64
rect 129 54 130 58
rect 134 54 135 58
rect 147 58 151 59
rect 163 58 169 61
rect 163 54 164 58
rect 168 54 169 58
rect 189 60 193 64
rect 189 55 193 56
rect 113 51 117 54
rect 147 51 151 54
rect 63 47 67 48
rect 72 47 73 51
rect 77 47 93 51
rect 97 47 113 51
rect 117 47 147 51
rect 151 50 185 51
rect 151 47 181 50
rect 53 43 57 46
rect 10 39 17 40
rect 10 25 14 39
rect 26 35 30 43
rect 18 34 30 35
rect 18 30 20 34
rect 24 30 30 34
rect 18 29 30 30
rect 3 22 7 23
rect 10 21 13 25
rect 17 21 18 25
rect 26 21 30 29
rect 34 39 43 43
rect 47 39 48 43
rect 34 38 48 39
rect 57 39 80 42
rect 53 38 80 39
rect 84 38 85 42
rect 34 25 38 38
rect 90 35 94 47
rect 181 43 185 46
rect 45 30 59 34
rect 63 31 90 34
rect 129 38 167 42
rect 185 39 190 42
rect 181 38 190 39
rect 129 34 135 38
rect 161 34 167 38
rect 63 30 94 31
rect 113 32 119 34
rect 34 24 40 25
rect 3 14 7 18
rect 12 18 18 21
rect 12 14 13 18
rect 17 14 18 18
rect 34 20 36 24
rect 45 24 51 30
rect 113 28 115 32
rect 129 30 130 34
rect 134 30 135 34
rect 145 30 146 34
rect 150 30 151 34
rect 161 30 162 34
rect 166 30 167 34
rect 113 26 119 28
rect 145 26 151 30
rect 45 20 46 24
rect 50 20 51 24
rect 56 24 95 26
rect 60 22 90 24
rect 60 20 61 22
rect 34 17 40 20
rect 56 17 61 20
rect 23 14 27 15
rect 3 8 7 10
rect 34 13 36 17
rect 40 13 56 17
rect 60 13 61 17
rect 89 20 90 22
rect 94 20 95 24
rect 89 17 95 20
rect 73 14 77 15
rect 23 8 27 10
rect 89 13 90 17
rect 94 13 95 17
rect 113 22 178 26
rect 182 22 183 26
rect 113 14 119 22
rect 126 18 130 19
rect 186 18 190 38
rect 136 14 137 18
rect 141 14 157 18
rect 161 14 190 18
rect 73 8 77 10
rect 126 11 130 14
rect -2 4 102 8
rect 106 7 126 8
rect 146 8 147 11
rect 130 7 147 8
rect 151 8 152 11
rect 166 8 167 11
rect 151 7 167 8
rect 171 8 172 11
rect 171 7 188 8
rect 106 4 188 7
rect 192 4 202 8
rect -2 0 202 4
<< ntransistor >>
rect 9 9 11 26
rect 19 9 21 26
rect 42 9 44 25
rect 52 9 54 25
rect 62 9 64 25
rect 69 9 71 25
rect 79 9 81 25
rect 86 9 88 25
rect 133 6 135 23
rect 143 6 145 23
rect 153 6 155 23
rect 163 6 165 23
<< ptransistor >>
rect 9 38 11 66
rect 19 38 21 66
rect 29 38 31 66
rect 39 38 41 66
rect 49 38 51 66
rect 59 38 61 66
rect 69 38 71 66
rect 79 46 81 66
rect 89 46 91 66
rect 99 46 101 66
rect 109 42 111 66
rect 119 38 121 66
rect 126 38 128 66
rect 136 38 138 66
rect 143 38 145 66
rect 153 38 155 66
rect 160 38 162 66
rect 170 38 172 66
rect 177 38 179 66
<< polycontact >>
rect 80 38 84 42
rect 20 30 24 34
rect 59 30 63 34
rect 90 31 94 35
rect 115 28 119 32
rect 130 30 134 34
rect 146 30 150 34
rect 162 30 166 34
rect 178 22 182 26
<< ndcontact >>
rect 3 18 7 22
rect 3 10 7 14
rect 13 21 17 25
rect 13 14 17 18
rect 23 10 27 14
rect 36 20 40 24
rect 36 13 40 17
rect 46 20 50 24
rect 56 20 60 24
rect 56 13 60 17
rect 73 10 77 14
rect 90 20 94 24
rect 90 13 94 17
rect 126 14 130 18
rect 126 7 130 11
rect 137 14 141 18
rect 147 7 151 11
rect 157 14 161 18
rect 167 7 171 11
<< pdcontact >>
rect 3 61 7 65
rect 3 54 7 58
rect 13 47 17 51
rect 13 40 17 44
rect 23 61 27 65
rect 23 54 27 58
rect 33 54 37 58
rect 33 47 37 51
rect 43 55 47 59
rect 43 39 47 43
rect 53 46 57 50
rect 53 39 57 43
rect 63 55 67 59
rect 63 48 67 52
rect 73 47 77 51
rect 83 55 87 59
rect 93 47 97 51
rect 103 55 107 59
rect 113 54 117 58
rect 113 47 117 51
rect 130 61 134 65
rect 130 54 134 58
rect 147 54 151 58
rect 147 47 151 51
rect 164 61 168 65
rect 164 54 168 58
rect 181 46 185 50
rect 181 39 185 43
<< psubstratepcontact >>
rect 102 4 106 8
rect 188 4 192 8
<< nsubstratencontact >>
rect 189 64 193 68
rect 189 56 193 60
<< psubstratepdiff >>
rect 101 8 107 24
rect 101 4 102 8
rect 106 4 107 8
rect 187 8 193 24
rect 101 3 107 4
rect 187 4 188 8
rect 192 4 193 8
rect 187 3 193 4
<< nsubstratendiff >>
rect 188 68 194 69
rect 188 64 189 68
rect 193 64 194 68
rect 188 60 194 64
rect 188 56 189 60
rect 193 56 194 60
rect 188 55 194 56
<< labels >>
rlabel polycontact 82 40 82 40 6 bn
rlabel metal1 15 19 15 19 6 bn
rlabel metal1 20 32 20 32 6 b
rlabel metal1 28 32 28 32 6 b
rlabel metal1 14 45 14 45 6 bn
rlabel metal1 35 53 35 53 6 bn
rlabel metal1 60 24 60 24 6 z
rlabel metal1 68 24 68 24 6 z
rlabel metal1 76 24 76 24 6 z
rlabel metal1 48 27 48 27 6 an
rlabel metal1 36 28 36 28 6 z
rlabel pdcontact 44 40 44 40 6 z
rlabel metal1 55 44 55 44 6 bn
rlabel pdcontact 34 49 34 49 6 bn
rlabel metal1 100 4 100 4 6 vss
rlabel metal1 116 24 116 24 6 a2
rlabel metal1 84 24 84 24 6 z
rlabel metal1 92 20 92 20 6 z
rlabel metal1 69 40 69 40 6 bn
rlabel metal1 115 53 115 53 6 an
rlabel metal1 100 68 100 68 6 vdd
rlabel metal1 124 24 124 24 6 a2
rlabel metal1 132 24 132 24 6 a2
rlabel metal1 140 24 140 24 6 a2
rlabel metal1 156 24 156 24 6 a2
rlabel metal1 148 28 148 28 6 a2
rlabel metal1 140 40 140 40 6 a1
rlabel metal1 148 40 148 40 6 a1
rlabel metal1 156 40 156 40 6 a1
rlabel metal1 132 36 132 36 6 a1
rlabel metal1 149 53 149 53 6 an
rlabel metal1 163 16 163 16 6 an
rlabel metal1 164 24 164 24 6 a2
rlabel metal1 172 24 172 24 6 a2
rlabel polycontact 180 24 180 24 6 a2
rlabel metal1 164 36 164 36 6 a1
rlabel metal1 164 40 164 40 6 a1
rlabel metal1 183 44 183 44 6 an
rlabel metal1 128 49 128 49 6 an
<< end >>
