.subckt noa2a22_x4 i0 i1 i2 i3 nq vdd vss
*   SPICE3 file   created from noa2a22_x4.ext -      technology: scmos
m00 w1     i0     w2     vdd p w=20u  l=2.3636u ad=100p     pd=30u      as=130p     ps=43u
m01 w2     i1     w1     vdd p w=20u  l=2.3636u ad=130p     pd=43u      as=100p     ps=30u
m02 vdd    i3     w2     vdd p w=20u  l=2.3636u ad=131.739p pd=38.8406u as=130p     ps=43u
m03 w2     i2     vdd    vdd p w=20u  l=2.3636u ad=130p     pd=43u      as=131.739p ps=38.8406u
m04 vdd    w1     w3     vdd p w=20u  l=2.3636u ad=131.739p pd=38.8406u as=160p     ps=56u
m05 nq     w3     vdd    vdd p w=39u  l=2.3636u ad=195p     pd=49u      as=256.891p ps=75.7391u
m06 vdd    w3     nq     vdd p w=39u  l=2.3636u ad=256.891p pd=75.7391u as=195p     ps=49u
m07 w4     i0     vss    vss n w=10u  l=2.3636u ad=50p      pd=20u      as=85.2941p ps=31.7647u
m08 w1     i1     w4     vss n w=10u  l=2.3636u ad=50p      pd=20u      as=50p      ps=20u
m09 w5     i3     w1     vss n w=10u  l=2.3636u ad=50p      pd=20u      as=50p      ps=20u
m10 vss    i2     w5     vss n w=10u  l=2.3636u ad=85.2941p pd=31.7647u as=50p      ps=20u
m11 vss    w1     w3     vss n w=10u  l=2.3636u ad=85.2941p pd=31.7647u as=80p      ps=36u
m12 nq     w3     vss    vss n w=19u  l=2.3636u ad=95p      pd=29u      as=162.059p ps=60.3529u
m13 vss    w3     nq     vss n w=19u  l=2.3636u ad=162.059p pd=60.3529u as=95p      ps=29u
C0  vss    nq     0.089f
C1  w2     vdd    0.319f
C2  i2     i0     0.062f
C3  w3     i1     0.033f
C4  nq     w1     0.076f
C5  w3     vdd    0.025f
C6  i3     i0     0.090f
C7  nq     i2     0.039f
C8  vss    w3     0.083f
C9  w1     w2     0.271f
C10 i1     vdd    0.008f
C11 vss    i1     0.029f
C12 w2     i2     0.013f
C13 w1     w3     0.309f
C14 w2     i3     0.013f
C15 i2     w3     0.132f
C16 w1     i1     0.262f
C17 vss    vdd    0.004f
C18 w3     i3     0.066f
C19 w2     i0     0.013f
C20 w1     vdd    0.212f
C21 i2     i1     0.090f
C22 vss    w1     0.036f
C23 i2     vdd    0.007f
C24 i3     i1     0.167f
C25 vss    i2     0.046f
C26 nq     w2     0.004f
C27 i3     vdd    0.007f
C28 i1     i0     0.327f
C29 w1     i2     0.166f
C30 w4     i1     0.018f
C31 nq     w3     0.105f
C32 vss    i3     0.034f
C33 w5     i3     0.018f
C34 i0     vdd    0.007f
C35 vss    i0     0.038f
C36 w1     i3     0.295f
C37 i2     i3     0.327f
C38 w2     i1     0.013f
C39 w1     i0     0.087f
C40 nq     vdd    0.165f
C42 nq     vss    0.012f
C43 w1     vss    0.048f
C44 i2     vss    0.037f
C45 w3     vss    0.071f
C46 i3     vss    0.043f
C47 i1     vss    0.043f
C48 i0     vss    0.037f
.ends
