.subckt nr4_x05 a b c d vdd vss z
*   SPICE3 file   created from nr4_x05.ext -      technology: scmos
m00 w1     d      z      vdd p w=39u  l=2.3636u ad=117p     pd=45u      as=243p     ps=94u
m01 w2     c      w1     vdd p w=39u  l=2.3636u ad=117p     pd=45u      as=117p     ps=45u
m02 w3     b      w2     vdd p w=39u  l=2.3636u ad=117p     pd=45u      as=117p     ps=45u
m03 vdd    a      w3     vdd p w=39u  l=2.3636u ad=312p     pd=94u      as=117p     ps=45u
m04 z      d      vss    vss n w=6u   l=2.3636u ad=30p      pd=16u      as=69p      ps=32u
m05 vss    c      z      vss n w=6u   l=2.3636u ad=69p      pd=32u      as=30p      ps=16u
m06 z      b      vss    vss n w=6u   l=2.3636u ad=30p      pd=16u      as=69p      ps=32u
m07 vss    a      z      vss n w=6u   l=2.3636u ad=69p      pd=32u      as=30p      ps=16u
C0  z      b      0.070f
C1  w3     vdd    0.011f
C2  w1     vdd    0.011f
C3  a      c      0.087f
C4  z      d      0.206f
C5  b      d      0.042f
C6  a      vdd    0.066f
C7  vss    a      0.009f
C8  c      vdd    0.008f
C9  vss    c      0.023f
C10 w2     a      0.006f
C11 z      a      0.030f
C12 w2     vdd    0.011f
C13 a      b      0.177f
C14 z      c      0.092f
C15 w1     d      0.011f
C16 a      d      0.056f
C17 b      c      0.208f
C18 z      vdd    0.031f
C19 vss    z      0.279f
C20 c      d      0.204f
C21 b      vdd    0.005f
C22 vss    b      0.037f
C23 w3     a      0.018f
C24 d      vdd    0.018f
C25 vss    d      0.016f
C27 z      vss    0.019f
C28 a      vss    0.024f
C29 b      vss    0.033f
C30 c      vss    0.036f
C31 d      vss    0.036f
.ends
