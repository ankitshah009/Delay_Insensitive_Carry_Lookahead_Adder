.subckt ts_x8 cmd i q vdd vss
*   SPICE3 file   created from ts_x8.ext -      technology: scmos
m00 q      w1     vdd    vdd p w=39u  l=2.3636u ad=195p     pd=49u      as=235.27p  ps=66.3907u
m01 vdd    w1     q      vdd p w=39u  l=2.3636u ad=235.27p  pd=66.3907u as=195p     ps=49u
m02 q      w1     vdd    vdd p w=39u  l=2.3636u ad=195p     pd=49u      as=235.27p  ps=66.3907u
m03 vdd    w1     q      vdd p w=39u  l=2.3636u ad=235.27p  pd=66.3907u as=195p     ps=49u
m04 w2     cmd    vdd    vdd p w=19u  l=2.3636u ad=152p     pd=54u      as=114.619p ps=32.3442u
m05 w1     w2     w3     vdd p w=19u  l=2.3636u ad=114.322p pd=37.3559u as=152p     ps=54u
m06 vdd    cmd    w1     vdd p w=20u  l=2.3636u ad=120.651p pd=34.0465u as=120.339p ps=39.322u
m07 w1     i      vdd    vdd p w=20u  l=2.3636u ad=120.339p pd=39.322u  as=120.651p ps=34.0465u
m08 q      w3     vss    vss n w=19u  l=2.3636u ad=95p      pd=29u      as=119.35p  ps=41.3204u
m09 vss    w3     q      vss n w=19u  l=2.3636u ad=119.35p  pd=41.3204u as=95p      ps=29u
m10 q      w3     vss    vss n w=19u  l=2.3636u ad=95p      pd=29u      as=119.35p  ps=41.3204u
m11 vss    w3     q      vss n w=19u  l=2.3636u ad=119.35p  pd=41.3204u as=95p      ps=29u
m12 w2     cmd    vss    vss n w=9u   l=2.3636u ad=72p      pd=34u      as=56.534p  ps=19.5728u
m13 vss    w2     w3     vss n w=9u   l=2.3636u ad=56.534p  pd=19.5728u as=53.6786p ps=23.7857u
m14 w3     i      vss    vss n w=9u   l=2.3636u ad=53.6786p pd=23.7857u as=56.534p  ps=19.5728u
m15 w1     cmd    w3     vss n w=10u  l=2.3636u ad=80p      pd=36u      as=59.6429p ps=26.4286u
C0  w3     q      0.070f
C1  i      w2     0.075f
C2  vss    vdd    0.007f
C3  w2     q      0.091f
C4  w3     cmd    0.364f
C5  vss    w1     0.029f
C6  i      vdd    0.034f
C7  w2     cmd    0.387f
C8  i      w1     0.253f
C9  q      vdd    0.436f
C10 q      w1     0.011f
C11 vdd    cmd    0.143f
C12 vss    i      0.012f
C13 cmd    w1     0.262f
C14 w3     w2     0.424f
C15 vss    q      0.203f
C16 w3     vdd    0.024f
C17 vss    cmd    0.067f
C18 w3     w1     0.346f
C19 i      cmd    0.224f
C20 w2     vdd    0.094f
C21 q      cmd    0.393f
C22 w2     w1     0.123f
C23 vss    w3     0.198f
C24 vdd    w1     0.193f
C25 w3     i      0.110f
C26 vss    w2     0.067f
C28 w3     vss    0.077f
C29 i      vss    0.039f
C30 w2     vss    0.056f
C31 q      vss    0.036f
C33 cmd    vss    0.094f
C34 w1     vss    0.089f
.ends
