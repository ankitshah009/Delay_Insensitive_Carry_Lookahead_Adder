magic
tech scmos
timestamp 1179385553
<< checkpaint >>
rect -22 -22 94 94
<< ab >>
rect 0 0 72 72
<< pwell >>
rect -4 -4 76 32
<< nwell >>
rect -4 32 76 76
<< polysilicon >>
rect 9 64 11 69
rect 19 64 21 69
rect 29 64 31 69
rect 39 64 41 69
rect 49 64 51 69
rect 59 56 61 61
rect 9 35 11 38
rect 19 35 21 38
rect 29 35 31 38
rect 39 35 41 38
rect 9 34 41 35
rect 9 33 29 34
rect 9 26 11 33
rect 19 30 29 33
rect 33 30 36 34
rect 40 30 41 34
rect 19 29 41 30
rect 19 26 21 29
rect 29 26 31 29
rect 39 26 41 29
rect 49 35 51 38
rect 59 35 61 38
rect 49 34 70 35
rect 49 33 65 34
rect 49 26 51 33
rect 59 30 65 33
rect 69 30 70 34
rect 59 29 70 30
rect 59 26 61 29
rect 9 8 11 13
rect 19 8 21 13
rect 29 8 31 13
rect 39 8 41 13
rect 49 10 51 15
rect 59 11 61 15
<< ndiffusion >>
rect 2 25 9 26
rect 2 21 3 25
rect 7 21 9 25
rect 2 18 9 21
rect 2 14 3 18
rect 7 14 9 18
rect 2 13 9 14
rect 11 25 19 26
rect 11 21 13 25
rect 17 21 19 25
rect 11 18 19 21
rect 11 14 13 18
rect 17 14 19 18
rect 11 13 19 14
rect 21 18 29 26
rect 21 14 23 18
rect 27 14 29 18
rect 21 13 29 14
rect 31 25 39 26
rect 31 21 33 25
rect 37 21 39 25
rect 31 18 39 21
rect 31 14 33 18
rect 37 14 39 18
rect 31 13 39 14
rect 41 20 49 26
rect 41 16 43 20
rect 47 16 49 20
rect 41 15 49 16
rect 51 25 59 26
rect 51 21 53 25
rect 57 21 59 25
rect 51 15 59 21
rect 61 20 69 26
rect 61 16 63 20
rect 67 16 69 20
rect 61 15 69 16
rect 41 13 47 15
<< pdiffusion >>
rect 2 63 9 64
rect 2 59 3 63
rect 7 59 9 63
rect 2 55 9 59
rect 2 51 3 55
rect 7 51 9 55
rect 2 38 9 51
rect 11 50 19 64
rect 11 46 13 50
rect 17 46 19 50
rect 11 43 19 46
rect 11 39 13 43
rect 17 39 19 43
rect 11 38 19 39
rect 21 63 29 64
rect 21 59 23 63
rect 27 59 29 63
rect 21 55 29 59
rect 21 51 23 55
rect 27 51 29 55
rect 21 38 29 51
rect 31 50 39 64
rect 31 46 33 50
rect 37 46 39 50
rect 31 43 39 46
rect 31 39 33 43
rect 37 39 39 43
rect 31 38 39 39
rect 41 63 49 64
rect 41 59 43 63
rect 47 59 49 63
rect 41 55 49 59
rect 41 51 43 55
rect 47 51 49 55
rect 41 38 49 51
rect 51 56 56 64
rect 51 51 59 56
rect 51 47 53 51
rect 57 47 59 51
rect 51 38 59 47
rect 61 55 69 56
rect 61 51 63 55
rect 67 51 69 55
rect 61 38 69 51
<< metal1 >>
rect -2 68 74 72
rect -2 64 62 68
rect 66 64 74 68
rect 3 63 7 64
rect 3 55 7 59
rect 23 63 27 64
rect 23 55 27 59
rect 43 63 47 64
rect 43 55 47 59
rect 63 55 67 64
rect 3 50 7 51
rect 13 50 17 51
rect 23 50 27 51
rect 33 50 39 51
rect 43 50 47 51
rect 13 43 17 46
rect 9 39 13 42
rect 37 46 39 50
rect 33 43 39 46
rect 17 39 33 42
rect 37 39 39 43
rect 9 38 39 39
rect 50 47 53 51
rect 57 47 58 51
rect 63 50 67 51
rect 18 26 22 38
rect 50 34 54 47
rect 58 37 70 43
rect 65 34 70 37
rect 28 30 29 34
rect 33 30 36 34
rect 40 30 57 34
rect 3 25 7 26
rect 3 18 7 21
rect 3 8 7 14
rect 13 25 39 26
rect 17 22 33 25
rect 13 18 17 21
rect 37 21 39 25
rect 53 25 57 30
rect 69 30 70 34
rect 65 29 70 30
rect 33 18 39 21
rect 13 13 17 14
rect 22 14 23 18
rect 27 14 28 18
rect 22 8 28 14
rect 37 14 39 18
rect 33 13 39 14
rect 43 20 47 21
rect 53 20 57 21
rect 63 20 67 21
rect 43 8 47 16
rect 63 8 67 16
rect -2 4 54 8
rect 58 4 62 8
rect 66 4 74 8
rect -2 0 74 4
<< ntransistor >>
rect 9 13 11 26
rect 19 13 21 26
rect 29 13 31 26
rect 39 13 41 26
rect 49 15 51 26
rect 59 15 61 26
<< ptransistor >>
rect 9 38 11 64
rect 19 38 21 64
rect 29 38 31 64
rect 39 38 41 64
rect 49 38 51 64
rect 59 38 61 56
<< polycontact >>
rect 29 30 33 34
rect 36 30 40 34
rect 65 30 69 34
<< ndcontact >>
rect 3 21 7 25
rect 3 14 7 18
rect 13 21 17 25
rect 13 14 17 18
rect 23 14 27 18
rect 33 21 37 25
rect 33 14 37 18
rect 43 16 47 20
rect 53 21 57 25
rect 63 16 67 20
<< pdcontact >>
rect 3 59 7 63
rect 3 51 7 55
rect 13 46 17 50
rect 13 39 17 43
rect 23 59 27 63
rect 23 51 27 55
rect 33 46 37 50
rect 33 39 37 43
rect 43 59 47 63
rect 43 51 47 55
rect 53 47 57 51
rect 63 51 67 55
<< psubstratepcontact >>
rect 54 4 58 8
rect 62 4 66 8
<< nsubstratencontact >>
rect 62 64 66 68
<< psubstratepdiff >>
rect 53 8 67 9
rect 53 4 54 8
rect 58 4 62 8
rect 66 4 67 8
rect 53 3 67 4
<< nsubstratendiff >>
rect 61 68 67 69
rect 61 64 62 68
rect 66 64 67 68
rect 61 63 67 64
<< labels >>
rlabel polycontact 30 32 30 32 6 an
rlabel metal1 12 40 12 40 6 z
rlabel metal1 20 32 20 32 6 z
rlabel metal1 28 24 28 24 6 z
rlabel metal1 28 40 28 40 6 z
rlabel metal1 36 4 36 4 6 vss
rlabel metal1 36 20 36 20 6 z
rlabel metal1 36 44 36 44 6 z
rlabel metal1 36 68 36 68 6 vdd
rlabel metal1 55 27 55 27 6 an
rlabel metal1 42 32 42 32 6 an
rlabel metal1 60 40 60 40 6 a
rlabel metal1 68 36 68 36 6 a
rlabel pdcontact 54 49 54 49 6 an
<< end >>
