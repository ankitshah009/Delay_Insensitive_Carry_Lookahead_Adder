magic
tech scmos
timestamp 1179386184
<< checkpaint >>
rect -22 -22 78 94
<< ab >>
rect 0 0 56 72
<< pwell >>
rect -4 -4 60 32
<< nwell >>
rect -4 32 60 76
<< polysilicon >>
rect 22 64 24 69
rect 32 64 34 69
rect 45 66 47 70
rect 9 57 11 61
rect 45 45 47 48
rect 41 44 47 45
rect 41 40 42 44
rect 46 40 47 44
rect 9 27 11 39
rect 22 37 24 40
rect 16 36 24 37
rect 16 32 17 36
rect 21 32 24 36
rect 32 37 34 40
rect 41 39 47 40
rect 32 35 37 37
rect 16 31 24 32
rect 35 34 41 35
rect 22 29 30 31
rect 9 26 16 27
rect 28 26 30 29
rect 35 30 36 34
rect 40 30 41 34
rect 35 29 41 30
rect 35 26 37 29
rect 45 26 47 39
rect 9 22 11 26
rect 15 22 16 26
rect 9 21 16 22
rect 9 18 11 21
rect 9 4 11 9
rect 45 12 47 17
rect 28 2 30 6
rect 35 2 37 6
<< ndiffusion >>
rect 21 25 28 26
rect 21 21 22 25
rect 26 21 28 25
rect 21 20 28 21
rect 2 17 9 18
rect 2 13 3 17
rect 7 13 9 17
rect 2 12 9 13
rect 4 9 9 12
rect 11 16 17 18
rect 11 9 19 16
rect 13 8 19 9
rect 13 4 14 8
rect 18 4 19 8
rect 23 6 28 20
rect 30 6 35 26
rect 37 22 45 26
rect 37 18 39 22
rect 43 18 45 22
rect 37 17 45 18
rect 47 25 54 26
rect 47 21 49 25
rect 53 21 54 25
rect 47 20 54 21
rect 47 17 52 20
rect 37 6 43 17
rect 13 3 19 4
<< pdiffusion >>
rect 36 65 45 66
rect 36 64 37 65
rect 14 58 22 64
rect 14 57 15 58
rect 4 52 9 57
rect 2 51 9 52
rect 2 47 3 51
rect 7 47 9 51
rect 2 44 9 47
rect 2 40 3 44
rect 7 40 9 44
rect 2 39 9 40
rect 11 54 15 57
rect 19 54 22 58
rect 11 40 22 54
rect 24 53 32 64
rect 24 49 26 53
rect 30 49 32 53
rect 24 45 32 49
rect 24 41 26 45
rect 30 41 32 45
rect 24 40 32 41
rect 34 61 37 64
rect 41 61 45 65
rect 34 58 45 61
rect 34 54 37 58
rect 41 54 45 58
rect 34 48 45 54
rect 47 54 52 66
rect 47 53 54 54
rect 47 49 49 53
rect 53 49 54 53
rect 47 48 54 49
rect 34 40 39 48
rect 11 39 16 40
<< metal1 >>
rect -2 68 58 72
rect -2 64 4 68
rect 8 65 58 68
rect 8 64 37 65
rect 14 58 20 64
rect 14 54 15 58
rect 19 54 20 58
rect 36 61 37 64
rect 41 64 58 65
rect 41 61 42 64
rect 36 58 42 61
rect 36 54 37 58
rect 41 54 42 58
rect 26 53 30 54
rect 3 51 7 52
rect 3 44 7 47
rect 17 49 26 50
rect 49 53 53 54
rect 17 46 30 49
rect 3 36 7 40
rect 26 45 30 46
rect 34 45 46 51
rect 2 32 17 36
rect 21 32 22 36
rect 2 17 6 32
rect 26 26 30 41
rect 42 44 46 45
rect 42 37 46 40
rect 49 34 53 49
rect 35 30 36 34
rect 40 30 53 34
rect 9 22 11 26
rect 15 22 18 26
rect 14 18 18 22
rect 21 25 30 26
rect 21 21 22 25
rect 26 22 30 25
rect 49 25 53 30
rect 39 22 43 23
rect 26 21 27 22
rect 49 20 53 21
rect 2 13 3 17
rect 7 13 8 17
rect 14 14 31 18
rect 39 8 43 18
rect -2 4 14 8
rect 18 4 48 8
rect 52 4 58 8
rect -2 0 58 4
<< ntransistor >>
rect 9 9 11 18
rect 28 6 30 26
rect 35 6 37 26
rect 45 17 47 26
<< ptransistor >>
rect 9 39 11 57
rect 22 40 24 64
rect 32 40 34 64
rect 45 48 47 66
<< polycontact >>
rect 42 40 46 44
rect 17 32 21 36
rect 36 30 40 34
rect 11 22 15 26
<< ndcontact >>
rect 22 21 26 25
rect 3 13 7 17
rect 14 4 18 8
rect 39 18 43 22
rect 49 21 53 25
<< pdcontact >>
rect 3 47 7 51
rect 3 40 7 44
rect 15 54 19 58
rect 26 49 30 53
rect 26 41 30 45
rect 37 61 41 65
rect 37 54 41 58
rect 49 49 53 53
<< psubstratepcontact >>
rect 48 4 52 8
<< nsubstratencontact >>
rect 4 64 8 68
<< psubstratepdiff >>
rect 47 8 53 9
rect 47 4 48 8
rect 52 4 53 8
rect 47 3 53 4
<< nsubstratendiff >>
rect 3 68 9 69
rect 3 64 4 68
rect 8 64 9 68
rect 3 63 9 64
<< labels >>
rlabel polycontact 20 34 20 34 6 bn
rlabel polycontact 38 32 38 32 6 an
rlabel pdcontact 5 42 5 42 6 bn
rlabel metal1 4 24 4 24 6 bn
rlabel metal1 20 16 20 16 6 b
rlabel polycontact 12 24 12 24 6 b
rlabel metal1 12 34 12 34 6 bn
rlabel metal1 20 48 20 48 6 z
rlabel metal1 28 4 28 4 6 vss
rlabel metal1 28 16 28 16 6 b
rlabel metal1 28 40 28 40 6 z
rlabel metal1 36 48 36 48 6 a
rlabel metal1 28 68 28 68 6 vdd
rlabel metal1 44 32 44 32 6 an
rlabel metal1 51 37 51 37 6 an
rlabel metal1 44 44 44 44 6 a
<< end >>
