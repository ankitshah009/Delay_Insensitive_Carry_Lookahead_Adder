magic
tech scmos
timestamp 1179386530
<< checkpaint >>
rect -22 -25 62 105
<< ab >>
rect 0 0 40 80
<< pwell >>
rect -4 -7 44 36
<< nwell >>
rect -4 36 44 87
<< polysilicon >>
rect 9 63 11 68
rect 19 63 21 68
rect 29 63 31 68
rect 9 36 11 53
rect 19 47 21 53
rect 19 46 25 47
rect 19 42 20 46
rect 24 42 25 46
rect 19 41 25 42
rect 9 35 17 36
rect 9 31 10 35
rect 14 31 17 35
rect 9 30 17 31
rect 15 27 17 30
rect 22 27 24 41
rect 29 39 31 53
rect 29 38 35 39
rect 29 34 30 38
rect 34 34 35 38
rect 29 33 35 34
rect 29 27 31 33
rect 15 12 17 17
rect 22 12 24 17
rect 29 12 31 17
<< ndiffusion >>
rect 10 23 15 27
rect 8 22 15 23
rect 8 18 9 22
rect 13 18 15 22
rect 8 17 15 18
rect 17 17 22 27
rect 24 17 29 27
rect 31 22 38 27
rect 31 18 33 22
rect 37 18 38 22
rect 31 17 38 18
<< pdiffusion >>
rect 4 59 9 63
rect 2 58 9 59
rect 2 54 3 58
rect 7 54 9 58
rect 2 53 9 54
rect 11 62 19 63
rect 11 58 13 62
rect 17 58 19 62
rect 11 53 19 58
rect 21 58 29 63
rect 21 54 23 58
rect 27 54 29 58
rect 21 53 29 54
rect 31 62 38 63
rect 31 58 33 62
rect 37 58 38 62
rect 31 53 38 58
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect -2 68 42 78
rect 2 58 7 63
rect 12 62 18 68
rect 12 58 13 62
rect 17 58 18 62
rect 32 62 38 68
rect 23 58 27 59
rect 32 58 33 62
rect 37 58 38 62
rect 2 54 3 58
rect 2 50 27 54
rect 2 22 6 50
rect 34 46 38 55
rect 17 42 20 46
rect 24 42 38 46
rect 10 35 14 36
rect 25 34 30 38
rect 10 30 14 31
rect 10 25 23 30
rect 34 25 38 38
rect 2 18 9 22
rect 13 18 14 22
rect 2 17 6 18
rect 18 17 23 25
rect 32 18 33 22
rect 37 18 38 22
rect 32 12 38 18
rect -2 2 42 12
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
<< ntransistor >>
rect 15 17 17 27
rect 22 17 24 27
rect 29 17 31 27
<< ptransistor >>
rect 9 53 11 63
rect 19 53 21 63
rect 29 53 31 63
<< polycontact >>
rect 20 42 24 46
rect 10 31 14 35
rect 30 34 34 38
<< ndcontact >>
rect 9 18 13 22
rect 33 18 37 22
<< pdcontact >>
rect 3 54 7 58
rect 13 58 17 62
rect 23 54 27 58
rect 33 58 37 62
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
<< psubstratepdiff >>
rect 0 2 40 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 40 2
rect 0 -3 40 -2
<< nsubstratendiff >>
rect 0 82 40 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 40 82
rect 0 77 40 78
<< labels >>
rlabel metal1 4 40 4 40 6 z
rlabel metal1 12 28 12 28 6 c
rlabel metal1 12 52 12 52 6 z
rlabel metal1 20 6 20 6 6 vss
rlabel metal1 20 24 20 24 6 c
rlabel metal1 28 36 28 36 6 a
rlabel metal1 28 44 28 44 6 b
rlabel metal1 20 44 20 44 6 b
rlabel metal1 20 52 20 52 6 z
rlabel metal1 20 74 20 74 6 vdd
rlabel metal1 36 28 36 28 6 a
rlabel metal1 36 52 36 52 6 b
<< end >>
