magic
tech scmos
timestamp 1182409238
<< checkpaint >>
rect -22 -25 222 105
<< ab >>
rect 0 0 200 80
<< pwell >>
rect -4 -7 204 36
<< nwell >>
rect -4 36 204 87
<< polysilicon >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 39 70 41 74
rect 49 70 51 74
rect 59 70 61 74
rect 69 70 71 74
rect 79 70 81 74
rect 89 70 91 74
rect 99 70 101 74
rect 109 70 111 74
rect 119 70 121 74
rect 126 70 128 74
rect 136 70 138 74
rect 143 70 145 74
rect 153 70 155 74
rect 160 70 162 74
rect 170 70 172 74
rect 177 70 179 74
rect 79 47 81 50
rect 89 47 91 50
rect 99 47 101 50
rect 79 46 101 47
rect 79 42 80 46
rect 84 45 101 46
rect 84 42 85 45
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 9 38 31 39
rect 9 37 20 38
rect 9 30 11 37
rect 19 34 20 37
rect 24 37 31 38
rect 39 39 41 42
rect 49 39 51 42
rect 59 39 61 42
rect 69 39 71 42
rect 79 41 85 42
rect 99 43 101 45
rect 109 43 111 46
rect 99 41 111 43
rect 79 39 81 41
rect 39 38 64 39
rect 39 37 59 38
rect 24 34 25 37
rect 19 33 25 34
rect 58 34 59 37
rect 63 34 64 38
rect 58 33 64 34
rect 19 30 21 33
rect 42 29 44 33
rect 52 29 54 33
rect 62 29 64 33
rect 69 37 81 39
rect 69 29 71 37
rect 79 29 81 37
rect 89 39 95 40
rect 89 36 90 39
rect 86 35 90 36
rect 94 35 95 39
rect 119 37 121 42
rect 126 39 128 42
rect 136 39 138 42
rect 126 38 138 39
rect 126 37 130 38
rect 86 34 95 35
rect 114 36 121 37
rect 86 29 88 34
rect 114 32 115 36
rect 119 32 121 36
rect 129 34 130 37
rect 134 37 138 38
rect 143 39 145 42
rect 153 39 155 42
rect 143 38 155 39
rect 134 34 135 37
rect 129 33 135 34
rect 114 31 121 32
rect 133 27 135 33
rect 143 34 146 38
rect 150 34 155 38
rect 143 33 155 34
rect 160 39 162 42
rect 170 39 172 42
rect 160 38 172 39
rect 160 34 162 38
rect 166 37 172 38
rect 166 34 167 37
rect 160 33 167 34
rect 143 27 145 33
rect 153 27 155 33
rect 163 27 165 33
rect 177 31 179 42
rect 177 30 183 31
rect 9 10 11 13
rect 19 10 21 13
rect 42 10 44 13
rect 52 10 54 13
rect 9 8 54 10
rect 62 8 64 13
rect 69 8 71 13
rect 79 8 81 13
rect 86 8 88 13
rect 177 26 178 30
rect 182 26 183 30
rect 177 25 183 26
rect 133 6 135 10
rect 143 6 145 10
rect 153 6 155 10
rect 163 6 165 10
<< ndiffusion >>
rect 2 26 9 30
rect 2 22 3 26
rect 7 22 9 26
rect 2 18 9 22
rect 2 14 3 18
rect 7 14 9 18
rect 2 13 9 14
rect 11 29 19 30
rect 11 25 13 29
rect 17 25 19 29
rect 11 22 19 25
rect 11 18 13 22
rect 17 18 19 22
rect 11 13 19 18
rect 21 18 29 30
rect 21 14 23 18
rect 27 14 29 18
rect 35 28 42 29
rect 35 24 36 28
rect 40 24 42 28
rect 35 21 42 24
rect 35 17 36 21
rect 40 17 42 21
rect 35 16 42 17
rect 21 13 29 14
rect 37 13 42 16
rect 44 28 52 29
rect 44 24 46 28
rect 50 24 52 28
rect 44 13 52 24
rect 54 28 62 29
rect 54 24 56 28
rect 60 24 62 28
rect 54 21 62 24
rect 54 17 56 21
rect 60 17 62 21
rect 54 13 62 17
rect 64 13 69 29
rect 71 18 79 29
rect 71 14 73 18
rect 77 14 79 18
rect 71 13 79 14
rect 81 13 86 29
rect 88 28 95 29
rect 88 24 90 28
rect 94 24 95 28
rect 88 21 95 24
rect 88 17 90 21
rect 94 17 95 21
rect 88 16 95 17
rect 124 22 133 27
rect 124 18 126 22
rect 130 18 133 22
rect 88 13 93 16
rect 124 15 133 18
rect 124 11 126 15
rect 130 11 133 15
rect 124 10 133 11
rect 135 22 143 27
rect 135 18 137 22
rect 141 18 143 22
rect 135 10 143 18
rect 145 15 153 27
rect 145 11 147 15
rect 151 11 153 15
rect 145 10 153 11
rect 155 22 163 27
rect 155 18 157 22
rect 161 18 163 22
rect 155 10 163 18
rect 165 15 173 27
rect 165 11 167 15
rect 171 11 173 15
rect 165 10 173 11
<< pdiffusion >>
rect 2 69 9 70
rect 2 65 3 69
rect 7 65 9 69
rect 2 62 9 65
rect 2 58 3 62
rect 7 58 9 62
rect 2 42 9 58
rect 11 55 19 70
rect 11 51 13 55
rect 17 51 19 55
rect 11 48 19 51
rect 11 44 13 48
rect 17 44 19 48
rect 11 42 19 44
rect 21 69 29 70
rect 21 65 23 69
rect 27 65 29 69
rect 21 62 29 65
rect 21 58 23 62
rect 27 58 29 62
rect 21 42 29 58
rect 31 62 39 70
rect 31 58 33 62
rect 37 58 39 62
rect 31 55 39 58
rect 31 51 33 55
rect 37 51 39 55
rect 31 42 39 51
rect 41 63 49 70
rect 41 59 43 63
rect 47 59 49 63
rect 41 47 49 59
rect 41 43 43 47
rect 47 43 49 47
rect 41 42 49 43
rect 51 54 59 70
rect 51 50 53 54
rect 57 50 59 54
rect 51 47 59 50
rect 51 43 53 47
rect 57 43 59 47
rect 51 42 59 43
rect 61 63 69 70
rect 61 59 63 63
rect 67 59 69 63
rect 61 56 69 59
rect 61 52 63 56
rect 67 52 69 56
rect 61 42 69 52
rect 71 55 79 70
rect 71 51 73 55
rect 77 51 79 55
rect 71 50 79 51
rect 81 63 89 70
rect 81 59 83 63
rect 87 59 89 63
rect 81 50 89 59
rect 91 55 99 70
rect 91 51 93 55
rect 97 51 99 55
rect 91 50 99 51
rect 101 63 109 70
rect 101 59 103 63
rect 107 59 109 63
rect 101 50 109 59
rect 71 42 76 50
rect 104 46 109 50
rect 111 62 119 70
rect 111 58 113 62
rect 117 58 119 62
rect 111 55 119 58
rect 111 51 113 55
rect 117 51 119 55
rect 111 46 119 51
rect 114 42 119 46
rect 121 42 126 70
rect 128 69 136 70
rect 128 65 130 69
rect 134 65 136 69
rect 128 62 136 65
rect 128 58 130 62
rect 134 58 136 62
rect 128 42 136 58
rect 138 42 143 70
rect 145 62 153 70
rect 145 58 147 62
rect 151 58 153 62
rect 145 55 153 58
rect 145 51 147 55
rect 151 51 153 55
rect 145 42 153 51
rect 155 42 160 70
rect 162 69 170 70
rect 162 65 164 69
rect 168 65 170 69
rect 162 62 170 65
rect 162 58 164 62
rect 168 58 170 62
rect 162 42 170 58
rect 172 42 177 70
rect 179 55 184 70
rect 179 54 186 55
rect 179 50 181 54
rect 185 50 186 54
rect 179 47 186 50
rect 179 43 181 47
rect 185 43 186 47
rect 179 42 186 43
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect 118 78 122 82
rect 126 78 130 82
rect 134 78 138 82
rect 142 78 146 82
rect 150 78 154 82
rect 158 78 162 82
rect 166 78 170 82
rect 174 78 178 82
rect 182 78 186 82
rect 190 78 194 82
rect 198 78 202 82
rect -2 69 202 78
rect -2 68 3 69
rect 2 65 3 68
rect 7 68 23 69
rect 7 65 8 68
rect 2 62 8 65
rect 2 58 3 62
rect 7 58 8 62
rect 22 65 23 68
rect 27 68 130 69
rect 27 65 28 68
rect 22 62 28 65
rect 129 65 130 68
rect 134 68 164 69
rect 134 65 135 68
rect 22 58 23 62
rect 27 58 28 62
rect 33 62 37 63
rect 42 59 43 63
rect 47 59 63 63
rect 67 59 83 63
rect 87 59 103 63
rect 107 59 108 63
rect 113 62 117 63
rect 33 55 37 58
rect 63 56 67 59
rect 12 51 13 55
rect 17 51 33 55
rect 37 54 57 55
rect 37 51 53 54
rect 12 48 17 51
rect 12 47 13 48
rect 10 44 13 47
rect 129 62 135 65
rect 163 65 164 68
rect 168 68 202 69
rect 168 65 169 68
rect 129 58 130 62
rect 134 58 135 62
rect 147 62 151 63
rect 163 62 169 65
rect 163 58 164 62
rect 168 58 169 62
rect 189 59 193 68
rect 113 55 117 58
rect 147 55 151 58
rect 63 51 67 52
rect 72 51 73 55
rect 77 51 93 55
rect 97 51 113 55
rect 117 51 147 55
rect 151 54 185 55
rect 151 51 181 54
rect 53 47 57 50
rect 10 43 17 44
rect 10 29 14 43
rect 26 39 30 47
rect 18 38 30 39
rect 18 34 20 38
rect 24 34 30 38
rect 18 33 30 34
rect 3 26 7 27
rect 10 25 13 29
rect 17 25 18 29
rect 26 25 30 33
rect 34 43 43 47
rect 47 43 48 47
rect 34 42 48 43
rect 57 43 80 46
rect 53 42 80 43
rect 84 42 85 46
rect 34 29 38 42
rect 90 39 94 51
rect 181 47 185 50
rect 45 34 59 38
rect 63 35 90 38
rect 129 42 167 46
rect 185 43 190 46
rect 181 42 190 43
rect 129 38 135 42
rect 161 38 167 42
rect 63 34 94 35
rect 113 36 119 38
rect 34 28 40 29
rect 3 18 7 22
rect 12 22 18 25
rect 12 18 13 22
rect 17 18 18 22
rect 34 24 36 28
rect 45 28 51 34
rect 113 32 115 36
rect 129 34 130 38
rect 134 34 135 38
rect 145 34 146 38
rect 150 34 151 38
rect 161 34 162 38
rect 166 34 167 38
rect 113 30 119 32
rect 145 30 151 34
rect 45 24 46 28
rect 50 24 51 28
rect 56 28 95 30
rect 60 26 90 28
rect 60 24 61 26
rect 34 21 40 24
rect 56 21 61 24
rect 23 18 27 19
rect 3 12 7 14
rect 34 17 36 21
rect 40 17 56 21
rect 60 17 61 21
rect 89 24 90 26
rect 94 24 95 28
rect 89 21 95 24
rect 73 18 77 19
rect 23 12 27 14
rect 89 17 90 21
rect 94 17 95 21
rect 113 26 178 30
rect 182 26 183 30
rect 113 18 119 26
rect 126 22 130 23
rect 186 22 190 42
rect 136 18 137 22
rect 141 18 157 22
rect 161 18 190 22
rect 73 12 77 14
rect 126 15 130 18
rect -2 11 126 12
rect 146 12 147 15
rect 130 11 147 12
rect 151 12 152 15
rect 166 12 167 15
rect 151 11 167 12
rect 171 12 172 15
rect 171 11 202 12
rect -2 2 202 11
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 122 2
rect 126 -2 130 2
rect 134 -2 138 2
rect 142 -2 146 2
rect 150 -2 154 2
rect 158 -2 162 2
rect 166 -2 170 2
rect 174 -2 178 2
rect 182 -2 186 2
rect 190 -2 194 2
rect 198 -2 202 2
<< ntransistor >>
rect 9 13 11 30
rect 19 13 21 30
rect 42 13 44 29
rect 52 13 54 29
rect 62 13 64 29
rect 69 13 71 29
rect 79 13 81 29
rect 86 13 88 29
rect 133 10 135 27
rect 143 10 145 27
rect 153 10 155 27
rect 163 10 165 27
<< ptransistor >>
rect 9 42 11 70
rect 19 42 21 70
rect 29 42 31 70
rect 39 42 41 70
rect 49 42 51 70
rect 59 42 61 70
rect 69 42 71 70
rect 79 50 81 70
rect 89 50 91 70
rect 99 50 101 70
rect 109 46 111 70
rect 119 42 121 70
rect 126 42 128 70
rect 136 42 138 70
rect 143 42 145 70
rect 153 42 155 70
rect 160 42 162 70
rect 170 42 172 70
rect 177 42 179 70
<< polycontact >>
rect 80 42 84 46
rect 20 34 24 38
rect 59 34 63 38
rect 90 35 94 39
rect 115 32 119 36
rect 130 34 134 38
rect 146 34 150 38
rect 162 34 166 38
rect 178 26 182 30
<< ndcontact >>
rect 3 22 7 26
rect 3 14 7 18
rect 13 25 17 29
rect 13 18 17 22
rect 23 14 27 18
rect 36 24 40 28
rect 36 17 40 21
rect 46 24 50 28
rect 56 24 60 28
rect 56 17 60 21
rect 73 14 77 18
rect 90 24 94 28
rect 90 17 94 21
rect 126 18 130 22
rect 126 11 130 15
rect 137 18 141 22
rect 147 11 151 15
rect 157 18 161 22
rect 167 11 171 15
<< pdcontact >>
rect 3 65 7 69
rect 3 58 7 62
rect 13 51 17 55
rect 13 44 17 48
rect 23 65 27 69
rect 23 58 27 62
rect 33 58 37 62
rect 33 51 37 55
rect 43 59 47 63
rect 43 43 47 47
rect 53 50 57 54
rect 53 43 57 47
rect 63 59 67 63
rect 63 52 67 56
rect 73 51 77 55
rect 83 59 87 63
rect 93 51 97 55
rect 103 59 107 63
rect 113 58 117 62
rect 113 51 117 55
rect 130 65 134 69
rect 130 58 134 62
rect 147 58 151 62
rect 147 51 151 55
rect 164 65 168 69
rect 164 58 168 62
rect 181 50 185 54
rect 181 43 185 47
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
rect 90 -2 94 2
rect 98 -2 102 2
rect 106 -2 110 2
rect 114 -2 118 2
rect 122 -2 126 2
rect 130 -2 134 2
rect 138 -2 142 2
rect 146 -2 150 2
rect 154 -2 158 2
rect 162 -2 166 2
rect 170 -2 174 2
rect 178 -2 182 2
rect 186 -2 190 2
rect 194 -2 198 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
rect 90 78 94 82
rect 98 78 102 82
rect 106 78 110 82
rect 114 78 118 82
rect 122 78 126 82
rect 130 78 134 82
rect 138 78 142 82
rect 146 78 150 82
rect 154 78 158 82
rect 162 78 166 82
rect 170 78 174 82
rect 178 78 182 82
rect 186 78 190 82
rect 194 78 198 82
<< psubstratepdiff >>
rect 0 2 200 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 122 2
rect 126 -2 130 2
rect 134 -2 138 2
rect 142 -2 146 2
rect 150 -2 154 2
rect 158 -2 162 2
rect 166 -2 170 2
rect 174 -2 178 2
rect 182 -2 186 2
rect 190 -2 194 2
rect 198 -2 200 2
rect 0 -3 200 -2
<< nsubstratendiff >>
rect 0 82 200 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect 118 78 122 82
rect 126 78 130 82
rect 134 78 138 82
rect 142 78 146 82
rect 150 78 154 82
rect 158 78 162 82
rect 166 78 170 82
rect 174 78 178 82
rect 182 78 186 82
rect 190 78 194 82
rect 198 78 200 82
rect 0 77 200 78
<< labels >>
rlabel polycontact 82 44 82 44 6 bn
rlabel metal1 15 23 15 23 6 bn
rlabel metal1 20 36 20 36 6 b
rlabel metal1 28 36 28 36 6 b
rlabel metal1 14 49 14 49 6 bn
rlabel metal1 60 28 60 28 6 z
rlabel metal1 48 31 48 31 6 an
rlabel metal1 36 32 36 32 6 z
rlabel pdcontact 44 44 44 44 6 z
rlabel pdcontact 34 53 34 53 6 bn
rlabel metal1 35 57 35 57 6 bn
rlabel metal1 55 48 55 48 6 bn
rlabel metal1 76 28 76 28 6 z
rlabel metal1 92 24 92 24 6 z
rlabel metal1 84 28 84 28 6 z
rlabel metal1 68 28 68 28 6 z
rlabel metal1 69 44 69 44 6 bn
rlabel metal1 100 6 100 6 6 vss
rlabel metal1 116 28 116 28 6 a2
rlabel metal1 124 28 124 28 6 a2
rlabel metal1 132 28 132 28 6 a2
rlabel metal1 132 40 132 40 6 a1
rlabel metal1 115 57 115 57 6 an
rlabel metal1 100 74 100 74 6 vdd
rlabel metal1 156 28 156 28 6 a2
rlabel metal1 140 28 140 28 6 a2
rlabel metal1 164 28 164 28 6 a2
rlabel metal1 148 32 148 32 6 a2
rlabel metal1 156 44 156 44 6 a1
rlabel metal1 148 44 148 44 6 a1
rlabel metal1 140 44 140 44 6 a1
rlabel metal1 164 40 164 40 6 a1
rlabel metal1 164 44 164 44 6 a1
rlabel metal1 149 57 149 57 6 an
rlabel metal1 163 20 163 20 6 an
rlabel polycontact 180 28 180 28 6 a2
rlabel metal1 172 28 172 28 6 a2
rlabel metal1 128 53 128 53 6 an
rlabel metal1 183 48 183 48 6 an
<< end >>
