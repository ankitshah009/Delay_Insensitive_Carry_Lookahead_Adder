magic
tech scmos
timestamp 1179386133
<< checkpaint >>
rect -22 -25 246 105
<< ab >>
rect 0 0 224 80
<< pwell >>
rect -4 -7 228 36
<< nwell >>
rect -4 36 228 87
<< polysilicon >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 39 70 41 74
rect 59 71 81 73
rect 59 65 61 71
rect 69 68 71 71
rect 79 68 81 71
rect 139 72 205 74
rect 139 69 141 72
rect 49 63 61 65
rect 49 60 51 63
rect 59 60 61 63
rect 89 64 91 69
rect 99 67 141 69
rect 99 64 101 67
rect 109 64 111 67
rect 119 64 121 67
rect 129 64 131 67
rect 139 64 141 67
rect 149 64 151 68
rect 163 64 165 68
rect 173 64 175 68
rect 183 64 185 68
rect 193 64 195 68
rect 203 64 205 72
rect 213 58 215 63
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 39 39 41 42
rect 9 38 41 39
rect 49 38 51 42
rect 59 38 61 42
rect 69 38 71 42
rect 79 39 81 42
rect 89 39 91 42
rect 79 38 91 39
rect 99 38 101 42
rect 109 38 111 42
rect 119 39 121 42
rect 119 38 125 39
rect 9 34 10 38
rect 14 34 18 38
rect 22 34 41 38
rect 79 34 84 38
rect 88 34 91 38
rect 119 34 120 38
rect 124 34 125 38
rect 129 37 131 42
rect 139 37 141 42
rect 149 39 151 42
rect 163 39 165 42
rect 173 39 175 42
rect 183 39 185 42
rect 193 39 195 42
rect 149 38 195 39
rect 9 33 41 34
rect 19 30 21 33
rect 29 30 31 33
rect 39 30 41 33
rect 49 30 51 34
rect 59 30 61 34
rect 69 30 71 34
rect 79 33 91 34
rect 79 30 81 33
rect 89 30 91 33
rect 99 30 101 34
rect 109 30 111 34
rect 119 33 125 34
rect 149 34 150 38
rect 154 34 158 38
rect 162 37 195 38
rect 203 39 205 42
rect 213 39 215 42
rect 162 34 181 37
rect 149 33 181 34
rect 79 13 81 17
rect 89 14 91 17
rect 99 14 101 17
rect 109 14 111 17
rect 89 12 111 14
rect 19 7 21 12
rect 29 7 31 12
rect 39 7 41 12
rect 49 8 51 12
rect 59 8 61 12
rect 69 8 71 12
rect 120 8 122 33
rect 149 30 151 33
rect 159 30 161 33
rect 169 30 171 33
rect 179 30 181 33
rect 203 33 215 39
rect 203 30 205 33
rect 213 30 215 33
rect 49 6 122 8
rect 149 11 151 16
rect 159 11 161 16
rect 169 11 171 16
rect 179 11 181 16
rect 203 14 205 19
rect 213 15 215 19
<< ndiffusion >>
rect 11 25 19 30
rect 11 21 13 25
rect 17 21 19 25
rect 11 17 19 21
rect 11 13 13 17
rect 17 13 19 17
rect 11 12 19 13
rect 21 29 29 30
rect 21 25 23 29
rect 27 25 29 29
rect 21 22 29 25
rect 21 18 23 22
rect 27 18 29 22
rect 21 12 29 18
rect 31 17 39 30
rect 31 13 33 17
rect 37 13 39 17
rect 31 12 39 13
rect 41 29 49 30
rect 41 25 43 29
rect 47 25 49 29
rect 41 22 49 25
rect 41 18 43 22
rect 47 18 49 22
rect 41 12 49 18
rect 51 29 59 30
rect 51 25 53 29
rect 57 25 59 29
rect 51 12 59 25
rect 61 21 69 30
rect 61 17 63 21
rect 67 17 69 21
rect 61 12 69 17
rect 71 29 79 30
rect 71 25 73 29
rect 77 25 79 29
rect 71 22 79 25
rect 71 18 73 22
rect 77 18 79 22
rect 71 17 79 18
rect 81 22 89 30
rect 81 18 83 22
rect 87 18 89 22
rect 81 17 89 18
rect 91 29 99 30
rect 91 25 93 29
rect 97 25 99 29
rect 91 17 99 25
rect 101 22 109 30
rect 101 18 103 22
rect 107 18 109 22
rect 101 17 109 18
rect 111 29 118 30
rect 111 25 113 29
rect 117 25 118 29
rect 111 24 118 25
rect 111 17 116 24
rect 71 12 76 17
rect 141 16 149 30
rect 151 29 159 30
rect 151 25 153 29
rect 157 25 159 29
rect 151 22 159 25
rect 151 18 153 22
rect 157 18 159 22
rect 151 16 159 18
rect 161 21 169 30
rect 161 17 163 21
rect 167 17 169 21
rect 161 16 169 17
rect 171 29 179 30
rect 171 25 173 29
rect 177 25 179 29
rect 171 22 179 25
rect 171 18 173 22
rect 177 18 179 22
rect 171 16 179 18
rect 181 29 189 30
rect 181 25 183 29
rect 187 25 189 29
rect 181 21 189 25
rect 181 17 183 21
rect 187 17 189 21
rect 195 24 203 30
rect 195 20 197 24
rect 201 20 203 24
rect 195 19 203 20
rect 205 29 213 30
rect 205 25 207 29
rect 211 25 213 29
rect 205 19 213 25
rect 215 24 222 30
rect 215 20 217 24
rect 221 20 222 24
rect 215 19 222 20
rect 181 16 189 17
rect 141 12 147 16
rect 141 8 142 12
rect 146 8 147 12
rect 141 7 147 8
<< pdiffusion >>
rect 4 55 9 70
rect 2 54 9 55
rect 2 50 3 54
rect 7 50 9 54
rect 2 47 9 50
rect 2 43 3 47
rect 7 43 9 47
rect 2 42 9 43
rect 11 69 19 70
rect 11 65 13 69
rect 17 65 19 69
rect 11 62 19 65
rect 11 58 13 62
rect 17 58 19 62
rect 11 42 19 58
rect 21 54 29 70
rect 21 50 23 54
rect 27 50 29 54
rect 21 47 29 50
rect 21 43 23 47
rect 27 43 29 47
rect 21 42 29 43
rect 31 69 39 70
rect 31 65 33 69
rect 37 65 39 69
rect 31 62 39 65
rect 31 58 33 62
rect 37 58 39 62
rect 31 42 39 58
rect 41 60 46 70
rect 64 60 69 68
rect 41 54 49 60
rect 41 50 43 54
rect 47 50 49 54
rect 41 47 49 50
rect 41 43 43 47
rect 47 43 49 47
rect 41 42 49 43
rect 51 54 59 60
rect 51 50 53 54
rect 57 50 59 54
rect 51 47 59 50
rect 51 43 53 47
rect 57 43 59 47
rect 51 42 59 43
rect 61 59 69 60
rect 61 55 63 59
rect 67 55 69 59
rect 61 52 69 55
rect 61 48 63 52
rect 67 48 69 52
rect 61 42 69 48
rect 71 54 79 68
rect 71 50 73 54
rect 77 50 79 54
rect 71 47 79 50
rect 71 43 73 47
rect 77 43 79 47
rect 71 42 79 43
rect 81 64 86 68
rect 81 63 89 64
rect 81 59 83 63
rect 87 59 89 63
rect 81 42 89 59
rect 91 47 99 64
rect 91 43 93 47
rect 97 43 99 47
rect 91 42 99 43
rect 101 55 109 64
rect 101 51 103 55
rect 107 51 109 55
rect 101 42 109 51
rect 111 47 119 64
rect 111 43 113 47
rect 117 43 119 47
rect 111 42 119 43
rect 121 55 129 64
rect 121 51 123 55
rect 127 51 129 55
rect 121 42 129 51
rect 131 47 139 64
rect 131 43 133 47
rect 137 43 139 47
rect 131 42 139 43
rect 141 54 149 64
rect 141 50 143 54
rect 147 50 149 54
rect 141 47 149 50
rect 141 43 143 47
rect 147 43 149 47
rect 141 42 149 43
rect 151 63 163 64
rect 151 59 157 63
rect 161 59 163 63
rect 151 42 163 59
rect 165 47 173 64
rect 165 43 167 47
rect 171 43 173 47
rect 165 42 173 43
rect 175 63 183 64
rect 175 59 177 63
rect 181 59 183 63
rect 175 42 183 59
rect 185 47 193 64
rect 185 43 187 47
rect 191 43 193 47
rect 185 42 193 43
rect 195 63 203 64
rect 195 59 197 63
rect 201 59 203 63
rect 195 42 203 59
rect 205 58 210 64
rect 205 54 213 58
rect 205 50 207 54
rect 211 50 213 54
rect 205 47 213 50
rect 205 43 207 47
rect 211 43 213 47
rect 205 42 213 43
rect 215 57 222 58
rect 215 53 217 57
rect 221 53 222 57
rect 215 49 222 53
rect 215 45 217 49
rect 221 45 222 49
rect 215 42 222 45
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect 118 78 122 82
rect 126 78 130 82
rect 134 78 138 82
rect 142 78 146 82
rect 150 78 154 82
rect 158 78 162 82
rect 166 78 170 82
rect 174 78 178 82
rect 182 78 186 82
rect 190 78 194 82
rect 198 78 202 82
rect 206 78 210 82
rect 214 78 218 82
rect 222 78 226 82
rect -2 69 226 78
rect -2 68 13 69
rect 17 68 33 69
rect 13 62 17 65
rect 13 57 17 58
rect 37 68 226 69
rect 33 62 37 65
rect 157 63 161 68
rect 33 57 37 58
rect 43 59 83 63
rect 87 59 88 63
rect 93 59 154 63
rect 3 54 7 55
rect 3 47 7 50
rect 23 54 27 55
rect 23 47 27 50
rect 7 43 23 46
rect 43 54 47 59
rect 43 47 47 50
rect 27 43 43 46
rect 3 42 47 43
rect 2 38 22 39
rect 2 34 10 38
rect 14 34 18 38
rect 2 33 22 34
rect 2 17 6 33
rect 43 30 47 42
rect 23 29 47 30
rect 13 25 17 26
rect 13 17 17 21
rect 27 26 43 29
rect 23 22 27 25
rect 43 22 47 25
rect 53 54 57 55
rect 53 47 57 50
rect 63 52 67 55
rect 63 47 67 48
rect 73 54 78 56
rect 93 55 97 59
rect 150 55 154 59
rect 157 58 161 59
rect 177 63 181 68
rect 196 63 202 68
rect 196 59 197 63
rect 201 59 202 63
rect 177 58 181 59
rect 217 57 221 68
rect 77 50 78 54
rect 73 47 78 50
rect 53 30 57 43
rect 77 43 78 47
rect 73 30 78 43
rect 84 51 97 55
rect 102 51 103 55
rect 107 51 123 55
rect 127 54 147 55
rect 127 51 143 54
rect 84 38 88 51
rect 142 50 143 51
rect 150 54 211 55
rect 150 51 207 54
rect 142 47 147 50
rect 207 47 211 50
rect 92 43 93 47
rect 97 46 98 47
rect 112 46 113 47
rect 97 43 113 46
rect 117 46 118 47
rect 132 46 133 47
rect 117 43 133 46
rect 137 43 138 47
rect 142 43 143 47
rect 147 43 167 47
rect 171 43 187 47
rect 191 43 192 47
rect 217 49 221 53
rect 217 44 221 45
rect 92 42 138 43
rect 84 33 88 34
rect 98 30 102 42
rect 146 38 166 39
rect 119 34 120 38
rect 124 34 135 38
rect 53 29 119 30
rect 57 26 73 29
rect 53 24 57 25
rect 77 26 93 29
rect 77 25 78 26
rect 92 25 93 26
rect 97 26 113 29
rect 97 25 98 26
rect 112 25 113 26
rect 117 25 119 29
rect 129 26 135 34
rect 146 34 150 38
rect 154 34 158 38
rect 162 34 166 38
rect 146 33 166 34
rect 146 25 150 33
rect 173 30 177 43
rect 153 29 177 30
rect 157 26 173 29
rect 157 25 158 26
rect 73 22 78 25
rect 153 22 158 25
rect 173 22 177 25
rect 47 18 63 21
rect 23 17 27 18
rect 33 17 37 18
rect 43 17 63 18
rect 67 17 68 21
rect 77 18 78 22
rect 82 18 83 22
rect 87 18 103 22
rect 107 18 153 22
rect 157 18 158 22
rect 163 21 167 22
rect 73 17 78 18
rect 173 17 177 18
rect 183 29 187 30
rect 207 29 211 43
rect 183 21 187 25
rect 13 12 17 13
rect 33 12 37 13
rect 163 12 167 17
rect 183 12 187 17
rect 197 24 201 25
rect 207 24 211 25
rect 217 24 221 25
rect 197 12 201 20
rect 217 12 221 20
rect -2 8 142 12
rect 146 8 226 12
rect -2 2 226 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 122 2
rect 126 -2 130 2
rect 134 -2 138 2
rect 142 -2 146 2
rect 150 -2 154 2
rect 158 -2 162 2
rect 166 -2 170 2
rect 174 -2 178 2
rect 182 -2 186 2
rect 190 -2 194 2
rect 198 -2 202 2
rect 206 -2 210 2
rect 214 -2 218 2
rect 222 -2 226 2
<< ntransistor >>
rect 19 12 21 30
rect 29 12 31 30
rect 39 12 41 30
rect 49 12 51 30
rect 59 12 61 30
rect 69 12 71 30
rect 79 17 81 30
rect 89 17 91 30
rect 99 17 101 30
rect 109 17 111 30
rect 149 16 151 30
rect 159 16 161 30
rect 169 16 171 30
rect 179 16 181 30
rect 203 19 205 30
rect 213 19 215 30
<< ptransistor >>
rect 9 42 11 70
rect 19 42 21 70
rect 29 42 31 70
rect 39 42 41 70
rect 49 42 51 60
rect 59 42 61 60
rect 69 42 71 68
rect 79 42 81 68
rect 89 42 91 64
rect 99 42 101 64
rect 109 42 111 64
rect 119 42 121 64
rect 129 42 131 64
rect 139 42 141 64
rect 149 42 151 64
rect 163 42 165 64
rect 173 42 175 64
rect 183 42 185 64
rect 193 42 195 64
rect 203 42 205 64
rect 213 42 215 58
<< polycontact >>
rect 10 34 14 38
rect 18 34 22 38
rect 84 34 88 38
rect 120 34 124 38
rect 150 34 154 38
rect 158 34 162 38
<< ndcontact >>
rect 13 21 17 25
rect 13 13 17 17
rect 23 25 27 29
rect 23 18 27 22
rect 33 13 37 17
rect 43 25 47 29
rect 43 18 47 22
rect 53 25 57 29
rect 63 17 67 21
rect 73 25 77 29
rect 73 18 77 22
rect 83 18 87 22
rect 93 25 97 29
rect 103 18 107 22
rect 113 25 117 29
rect 153 25 157 29
rect 153 18 157 22
rect 163 17 167 21
rect 173 25 177 29
rect 173 18 177 22
rect 183 25 187 29
rect 183 17 187 21
rect 197 20 201 24
rect 207 25 211 29
rect 217 20 221 24
rect 142 8 146 12
<< pdcontact >>
rect 3 50 7 54
rect 3 43 7 47
rect 13 65 17 69
rect 13 58 17 62
rect 23 50 27 54
rect 23 43 27 47
rect 33 65 37 69
rect 33 58 37 62
rect 43 50 47 54
rect 43 43 47 47
rect 53 50 57 54
rect 53 43 57 47
rect 63 55 67 59
rect 63 48 67 52
rect 73 50 77 54
rect 73 43 77 47
rect 83 59 87 63
rect 93 43 97 47
rect 103 51 107 55
rect 113 43 117 47
rect 123 51 127 55
rect 133 43 137 47
rect 143 50 147 54
rect 143 43 147 47
rect 157 59 161 63
rect 167 43 171 47
rect 177 59 181 63
rect 187 43 191 47
rect 197 59 201 63
rect 207 50 211 54
rect 207 43 211 47
rect 217 53 221 57
rect 217 45 221 49
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
rect 90 -2 94 2
rect 98 -2 102 2
rect 106 -2 110 2
rect 114 -2 118 2
rect 122 -2 126 2
rect 130 -2 134 2
rect 138 -2 142 2
rect 146 -2 150 2
rect 154 -2 158 2
rect 162 -2 166 2
rect 170 -2 174 2
rect 178 -2 182 2
rect 186 -2 190 2
rect 194 -2 198 2
rect 202 -2 206 2
rect 210 -2 214 2
rect 218 -2 222 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
rect 90 78 94 82
rect 98 78 102 82
rect 106 78 110 82
rect 114 78 118 82
rect 122 78 126 82
rect 130 78 134 82
rect 138 78 142 82
rect 146 78 150 82
rect 154 78 158 82
rect 162 78 166 82
rect 170 78 174 82
rect 178 78 182 82
rect 186 78 190 82
rect 194 78 198 82
rect 202 78 206 82
rect 210 78 214 82
rect 218 78 222 82
<< psubstratepdiff >>
rect 0 2 224 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 122 2
rect 126 -2 130 2
rect 134 -2 138 2
rect 142 -2 146 2
rect 150 -2 154 2
rect 158 -2 162 2
rect 166 -2 170 2
rect 174 -2 178 2
rect 182 -2 186 2
rect 190 -2 194 2
rect 198 -2 202 2
rect 206 -2 210 2
rect 214 -2 218 2
rect 222 -2 224 2
rect 0 -3 224 -2
<< nsubstratendiff >>
rect 0 82 224 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect 118 78 122 82
rect 126 78 130 82
rect 134 78 138 82
rect 142 78 146 82
rect 150 78 154 82
rect 158 78 162 82
rect 166 78 170 82
rect 174 78 178 82
rect 182 78 186 82
rect 190 78 194 82
rect 198 78 202 82
rect 206 78 210 82
rect 214 78 218 82
rect 222 78 224 82
rect 0 77 224 78
<< labels >>
rlabel metal1 4 28 4 28 6 a1
rlabel metal1 25 23 25 23 6 a1n
rlabel polycontact 12 36 12 36 6 a1
rlabel polycontact 20 36 20 36 6 a1
rlabel metal1 5 48 5 48 6 a1n
rlabel metal1 25 48 25 48 6 a1n
rlabel metal1 55 19 55 19 6 a1n
rlabel metal1 68 28 68 28 6 z
rlabel metal1 60 28 60 28 6 z
rlabel metal1 65 55 65 55 6 a1n
rlabel metal1 45 40 45 40 6 a1n
rlabel metal1 84 28 84 28 6 z
rlabel metal1 92 28 92 28 6 z
rlabel metal1 108 28 108 28 6 z
rlabel metal1 76 36 76 36 6 z
rlabel metal1 100 36 100 36 6 z
rlabel metal1 108 44 108 44 6 z
rlabel metal1 86 44 86 44 6 sn
rlabel metal1 65 61 65 61 6 a1n
rlabel metal1 112 6 112 6 6 vss
rlabel ndcontact 116 28 116 28 6 z
rlabel metal1 148 32 148 32 6 a0
rlabel metal1 124 36 124 36 6 s
rlabel metal1 132 32 132 32 6 s
rlabel metal1 132 44 132 44 6 z
rlabel metal1 124 44 124 44 6 z
rlabel pdcontact 116 44 116 44 6 z
rlabel metal1 144 49 144 49 6 a0n
rlabel pdcontact 124 53 124 53 6 a0n
rlabel metal1 112 74 112 74 6 vdd
rlabel metal1 120 20 120 20 6 a0n
rlabel metal1 155 24 155 24 6 a0n
rlabel metal1 164 36 164 36 6 a0
rlabel metal1 156 36 156 36 6 a0
rlabel metal1 175 32 175 32 6 a0n
rlabel metal1 167 45 167 45 6 a0n
rlabel metal1 209 39 209 39 6 sn
<< end >>
