.subckt xor2_x05 a b vdd vss z
*   SPICE3 file   created from xor2_x05.ext -      technology: scmos
m00 z      an     bn     vdd p w=20u  l=2.3636u ad=100p     pd=30u      as=118p     ps=56u
m01 an     bn     z      vdd p w=20u  l=2.3636u ad=100p     pd=30u      as=100p     ps=30u
m02 vdd    a      an     vdd p w=20u  l=2.3636u ad=300p     pd=58u      as=100p     ps=30u
m03 bn     b      vdd    vdd p w=20u  l=2.3636u ad=118p     pd=56u      as=300p     ps=58u
m04 w1     an     vss    vss n w=9u   l=2.3636u ad=27p      pd=15u      as=77p      ps=31.3333u
m05 z      bn     w1     vss n w=9u   l=2.3636u ad=45p      pd=19u      as=27p      ps=15u
m06 an     b      z      vss n w=9u   l=2.3636u ad=45p      pd=19u      as=45p      ps=19u
m07 vss    a      an     vss n w=9u   l=2.3636u ad=77p      pd=31.3333u as=45p      ps=19u
m08 bn     b      vss    vss n w=9u   l=2.3636u ad=63p      pd=34u      as=77p      ps=31.3333u
C0  vss    b      0.015f
C1  w1     z      0.011f
C2  vss    a      0.063f
C3  b      z      0.021f
C4  z      a      0.033f
C5  b      bn     0.207f
C6  vss    an     0.066f
C7  z      an     0.306f
C8  a      bn     0.304f
C9  b      vdd    0.162f
C10 bn     an     0.427f
C11 a      vdd    0.004f
C12 an     vdd    0.019f
C13 vss    z      0.152f
C14 b      a      0.097f
C15 vss    bn     0.048f
C16 z      bn     0.195f
C17 b      an     0.053f
C18 a      an     0.171f
C19 z      vdd    0.036f
C20 bn     vdd    0.262f
C22 b      vss    0.049f
C23 z      vss    0.021f
C24 a      vss    0.040f
C25 bn     vss    0.060f
C26 an     vss    0.053f
.ends
