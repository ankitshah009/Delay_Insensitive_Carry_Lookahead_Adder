.subckt oa22_x2 i0 i1 i2 q vdd vss
*   SPICE3 file   created from oa22_x2.ext -      technology: scmos
m00 w1     i0     w2     vdd p w=20u  l=2.3636u ad=100p     pd=30.7692u as=120.339p ps=39.322u
m01 w2     i1     w1     vdd p w=19u  l=2.3636u ad=114.322p pd=37.3559u as=95p      ps=29.2308u
m02 vdd    i2     w2     vdd p w=20u  l=2.3636u ad=119.322p pd=33.2203u as=120.339p ps=39.322u
m03 q      w1     vdd    vdd p w=39u  l=2.3636u ad=312p     pd=94u      as=232.678p ps=64.7797u
m04 w3     i0     vss    vss n w=10u  l=2.3636u ad=50p      pd=21.0526u as=77.6316p ps=28.9474u
m05 w1     i1     w3     vss n w=9u   l=2.3636u ad=45p      pd=19u      as=45p      ps=18.9474u
m06 vss    i2     w1     vss n w=9u   l=2.3636u ad=69.8684p pd=26.0526u as=45p      ps=19u
m07 q      w1     vss    vss n w=19u  l=2.3636u ad=152p     pd=54u      as=147.5p   ps=55u
C0  w2     i1     0.013f
C1  q      i0     0.039f
C2  vss    w1     0.034f
C3  q      vdd    0.080f
C4  i2     i0     0.079f
C5  w2     w1     0.143f
C6  i1     w1     0.268f
C7  i2     vdd    0.076f
C8  vss    q      0.065f
C9  i0     vdd    0.007f
C10 q      w2     0.017f
C11 w3     i1     0.016f
C12 vss    i2     0.043f
C13 q      i1     0.054f
C14 vss    i0     0.038f
C15 w2     i2     0.036f
C16 i2     i1     0.129f
C17 w2     i0     0.013f
C18 q      w1     0.186f
C19 i2     w1     0.385f
C20 i1     i0     0.302f
C21 w2     vdd    0.164f
C22 i0     w1     0.108f
C23 i1     vdd    0.008f
C24 w1     vdd    0.042f
C25 vss    i1     0.029f
C26 q      i2     0.334f
C28 q      vss    0.011f
C29 i2     vss    0.039f
C30 i1     vss    0.039f
C31 i0     vss    0.037f
C32 w1     vss    0.047f
.ends
