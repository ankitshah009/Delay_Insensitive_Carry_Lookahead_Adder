magic
tech scmos
timestamp 1179385433
<< checkpaint >>
rect -22 -25 118 105
<< ab >>
rect 0 0 96 80
<< pwell >>
rect -4 -7 100 36
<< nwell >>
rect -4 36 100 87
<< polysilicon >>
rect 9 69 11 74
rect 19 69 21 74
rect 29 69 31 74
rect 39 69 41 74
rect 50 69 52 74
rect 60 69 62 74
rect 71 61 73 66
rect 81 61 83 65
rect 50 47 52 52
rect 9 39 11 43
rect 19 39 21 43
rect 29 39 31 47
rect 39 39 41 47
rect 50 46 56 47
rect 50 42 51 46
rect 55 42 56 46
rect 50 41 56 42
rect 60 43 62 52
rect 71 43 73 46
rect 60 41 73 43
rect 81 43 83 46
rect 81 42 87 43
rect 9 38 15 39
rect 9 34 10 38
rect 14 34 15 38
rect 9 33 15 34
rect 19 38 31 39
rect 19 34 26 38
rect 30 34 31 38
rect 19 33 31 34
rect 12 30 14 33
rect 19 30 21 33
rect 29 30 31 33
rect 36 38 46 39
rect 36 34 41 38
rect 45 34 46 38
rect 36 33 46 34
rect 36 30 38 33
rect 51 29 53 41
rect 64 37 70 41
rect 64 34 65 37
rect 58 33 65 34
rect 69 33 70 37
rect 81 38 82 42
rect 86 38 87 42
rect 81 37 87 38
rect 81 34 83 37
rect 58 32 70 33
rect 58 29 60 32
rect 68 29 70 32
rect 75 32 83 34
rect 75 29 77 32
rect 12 6 14 10
rect 19 6 21 10
rect 29 6 31 10
rect 36 6 38 10
rect 51 9 53 14
rect 58 9 60 14
rect 68 13 70 18
rect 75 13 77 18
<< ndiffusion >>
rect 3 12 12 30
rect 3 8 5 12
rect 9 10 12 12
rect 14 10 19 30
rect 21 22 29 30
rect 21 18 23 22
rect 27 18 29 22
rect 21 10 29 18
rect 31 10 36 30
rect 38 29 49 30
rect 38 22 51 29
rect 38 18 43 22
rect 47 18 51 22
rect 38 15 51 18
rect 38 11 43 15
rect 47 14 51 15
rect 53 14 58 29
rect 60 23 68 29
rect 60 19 62 23
rect 66 19 68 23
rect 60 18 68 19
rect 70 18 75 29
rect 77 23 88 29
rect 77 19 82 23
rect 86 19 88 23
rect 77 18 88 19
rect 60 14 65 18
rect 47 11 49 14
rect 38 10 49 11
rect 9 8 10 10
rect 3 7 10 8
<< pdiffusion >>
rect 2 68 9 69
rect 2 64 3 68
rect 7 64 9 68
rect 2 61 9 64
rect 2 57 3 61
rect 7 57 9 61
rect 2 43 9 57
rect 11 62 19 69
rect 11 58 13 62
rect 17 58 19 62
rect 11 55 19 58
rect 11 51 13 55
rect 17 51 19 55
rect 11 43 19 51
rect 21 68 29 69
rect 21 64 23 68
rect 27 64 29 68
rect 21 61 29 64
rect 21 57 23 61
rect 27 57 29 61
rect 21 47 29 57
rect 31 62 39 69
rect 31 58 33 62
rect 37 58 39 62
rect 31 55 39 58
rect 31 51 33 55
rect 37 51 39 55
rect 31 47 39 51
rect 41 68 50 69
rect 41 64 43 68
rect 47 64 50 68
rect 41 61 50 64
rect 41 57 43 61
rect 47 57 50 61
rect 41 52 50 57
rect 52 57 60 69
rect 52 53 54 57
rect 58 53 60 57
rect 52 52 60 53
rect 62 68 69 69
rect 62 64 64 68
rect 68 64 69 68
rect 62 61 69 64
rect 62 57 64 61
rect 68 57 71 61
rect 62 52 71 57
rect 41 47 48 52
rect 21 43 27 47
rect 64 46 71 52
rect 73 60 81 61
rect 73 56 75 60
rect 79 56 81 60
rect 73 53 81 56
rect 73 49 75 53
rect 79 49 81 53
rect 73 46 81 49
rect 83 60 90 61
rect 83 56 85 60
rect 89 56 90 60
rect 83 53 90 56
rect 83 49 85 53
rect 89 49 90 53
rect 83 46 90 49
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect -2 68 98 78
rect 2 64 3 68
rect 7 64 8 68
rect 2 61 8 64
rect 22 64 23 68
rect 27 64 28 68
rect 2 57 3 61
rect 7 57 8 61
rect 13 62 17 63
rect 13 55 17 58
rect 22 61 28 64
rect 42 64 43 68
rect 47 64 48 68
rect 22 57 23 61
rect 27 57 28 61
rect 33 62 39 63
rect 37 58 39 62
rect 2 51 13 54
rect 33 55 39 58
rect 42 61 48 64
rect 42 57 43 61
rect 47 57 48 61
rect 63 64 64 68
rect 68 64 69 68
rect 63 61 69 64
rect 54 57 58 58
rect 63 57 64 61
rect 68 57 69 61
rect 75 60 80 61
rect 17 51 33 54
rect 37 51 39 55
rect 79 56 80 60
rect 75 53 80 56
rect 2 50 39 51
rect 2 22 6 50
rect 42 49 75 53
rect 79 49 80 53
rect 84 60 90 68
rect 84 56 85 60
rect 89 56 90 60
rect 84 53 90 56
rect 84 49 85 53
rect 89 49 90 53
rect 17 42 31 46
rect 10 38 14 39
rect 25 38 31 42
rect 42 39 46 49
rect 49 42 51 46
rect 55 42 87 46
rect 25 34 26 38
rect 30 34 31 38
rect 41 38 46 39
rect 81 38 82 42
rect 86 38 87 42
rect 45 34 46 38
rect 10 30 14 34
rect 41 30 46 34
rect 65 37 71 38
rect 69 33 71 37
rect 81 34 87 38
rect 65 30 71 33
rect 10 26 58 30
rect 65 26 87 30
rect 54 23 58 26
rect 2 18 23 22
rect 27 18 28 22
rect 42 18 43 22
rect 47 18 48 22
rect 54 19 62 23
rect 66 19 67 23
rect 42 15 48 18
rect 74 17 78 26
rect 81 19 82 23
rect 86 19 87 23
rect 42 12 43 15
rect -2 8 5 12
rect 9 11 43 12
rect 47 12 48 15
rect 81 12 87 19
rect 47 11 98 12
rect 9 8 98 11
rect -2 2 98 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
<< ntransistor >>
rect 12 10 14 30
rect 19 10 21 30
rect 29 10 31 30
rect 36 10 38 30
rect 51 14 53 29
rect 58 14 60 29
rect 68 18 70 29
rect 75 18 77 29
<< ptransistor >>
rect 9 43 11 69
rect 19 43 21 69
rect 29 47 31 69
rect 39 47 41 69
rect 50 52 52 69
rect 60 52 62 69
rect 71 46 73 61
rect 81 46 83 61
<< polycontact >>
rect 51 42 55 46
rect 10 34 14 38
rect 26 34 30 38
rect 41 34 45 38
rect 65 33 69 37
rect 82 38 86 42
<< ndcontact >>
rect 5 8 9 12
rect 23 18 27 22
rect 43 18 47 22
rect 43 11 47 15
rect 62 19 66 23
rect 82 19 86 23
<< pdcontact >>
rect 3 64 7 68
rect 3 57 7 61
rect 13 58 17 62
rect 13 51 17 55
rect 23 64 27 68
rect 23 57 27 61
rect 33 58 37 62
rect 33 51 37 55
rect 43 64 47 68
rect 43 57 47 61
rect 54 53 58 57
rect 64 64 68 68
rect 64 57 68 61
rect 75 56 79 60
rect 75 49 79 53
rect 85 56 89 60
rect 85 49 89 53
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
rect 90 -2 94 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
rect 90 78 94 82
<< psubstratepdiff >>
rect 0 2 96 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 96 2
rect 0 -3 96 -2
<< nsubstratendiff >>
rect 0 82 96 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 96 82
rect 0 77 96 78
<< labels >>
rlabel ntransistor 13 22 13 22 6 an
rlabel ptransistor 40 53 40 53 6 an
rlabel metal1 12 20 12 20 6 z
rlabel metal1 12 32 12 32 6 an
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 52 12 52 6 z
rlabel metal1 20 20 20 20 6 z
rlabel metal1 20 44 20 44 6 b
rlabel metal1 28 40 28 40 6 b
rlabel metal1 28 52 28 52 6 z
rlabel metal1 20 52 20 52 6 z
rlabel metal1 48 6 48 6 6 vss
rlabel polycontact 52 44 52 44 6 a1
rlabel metal1 56 53 56 53 6 an
rlabel metal1 44 39 44 39 6 an
rlabel metal1 36 56 36 56 6 z
rlabel metal1 48 74 48 74 6 vdd
rlabel metal1 60 21 60 21 6 an
rlabel metal1 76 24 76 24 6 a2
rlabel metal1 68 32 68 32 6 a2
rlabel metal1 60 44 60 44 6 a1
rlabel metal1 68 44 68 44 6 a1
rlabel metal1 76 44 76 44 6 a1
rlabel metal1 84 28 84 28 6 a2
rlabel polycontact 84 40 84 40 6 a1
rlabel metal1 77 55 77 55 6 an
rlabel metal1 61 51 61 51 6 an
<< end >>
