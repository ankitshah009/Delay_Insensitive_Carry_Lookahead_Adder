.subckt iv1v0x6 a vdd vss z
*   SPICE3 file   created from iv1v0x6.ext -      technology: scmos
m00 z      a      vdd    vdd p w=26u  l=2.3636u ad=130p     pd=36u      as=182p     ps=66u
m01 vdd    a      z      vdd p w=26u  l=2.3636u ad=182p     pd=66u      as=130p     ps=36u
m02 z      a      vdd    vdd p w=26u  l=2.3636u ad=130p     pd=36u      as=182p     ps=66u
m03 w1     vdd    z      vdd p w=26u  l=2.3636u ad=182p     pd=66u      as=130p     ps=36u
m04 z      a      vss    vss n w=18u  l=2.3636u ad=90p      pd=28u      as=126p     ps=50u
m05 vss    a      z      vss n w=18u  l=2.3636u ad=126p     pd=50u      as=90p      ps=28u
m06 z      a      vss    vss n w=18u  l=2.3636u ad=90p      pd=28u      as=126p     ps=50u
m07 w2     vss    z      vss n w=18u  l=2.3636u ad=126p     pd=50u      as=90p      ps=28u
C0  vss    z      0.222f
C1  vss    vdd    0.047f
C2  z      vdd    0.179f
C3  vss    a      0.145f
C4  z      a      0.392f
C5  a      vdd    0.141f
C7  z      vss    0.010f
C8  a      vss    0.194f
.ends
