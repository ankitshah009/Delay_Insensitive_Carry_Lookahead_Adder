magic
tech scmos
timestamp 1179386234
<< checkpaint >>
rect -22 -25 62 105
<< ab >>
rect 0 0 40 80
<< pwell >>
rect -4 -7 44 36
<< nwell >>
rect -4 36 44 87
<< polysilicon >>
rect 9 64 15 65
rect 9 60 10 64
rect 14 60 15 64
rect 9 59 15 60
rect 9 56 11 59
rect 19 56 21 61
rect 29 56 31 61
rect 9 30 11 42
rect 19 39 21 42
rect 16 38 23 39
rect 16 34 18 38
rect 22 34 23 38
rect 16 33 23 34
rect 16 30 18 33
rect 29 31 31 42
rect 28 30 34 31
rect 28 26 29 30
rect 33 26 34 30
rect 28 25 34 26
rect 28 22 30 25
rect 9 14 11 18
rect 16 14 18 18
rect 28 10 30 15
<< ndiffusion >>
rect 2 29 9 30
rect 2 25 3 29
rect 7 25 9 29
rect 2 24 9 25
rect 4 18 9 24
rect 11 18 16 30
rect 18 22 26 30
rect 18 18 28 22
rect 20 15 28 18
rect 30 21 38 22
rect 30 17 33 21
rect 37 17 38 21
rect 30 15 38 17
rect 20 12 26 15
rect 20 8 21 12
rect 25 8 26 12
rect 20 7 26 8
<< pdiffusion >>
rect 2 72 8 73
rect 2 68 3 72
rect 7 68 8 72
rect 2 67 8 68
rect 21 68 27 69
rect 2 56 7 67
rect 21 64 22 68
rect 26 64 27 68
rect 21 63 27 64
rect 23 56 27 63
rect 2 42 9 56
rect 11 54 19 56
rect 11 50 13 54
rect 17 50 19 54
rect 11 47 19 50
rect 11 43 13 47
rect 17 43 19 47
rect 11 42 19 43
rect 21 42 29 56
rect 31 55 38 56
rect 31 51 33 55
rect 37 51 38 55
rect 31 50 38 51
rect 31 42 36 50
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect -2 72 42 78
rect -2 68 3 72
rect 7 68 42 72
rect 9 63 10 64
rect 2 60 10 63
rect 14 60 15 64
rect 22 63 26 64
rect 2 58 15 60
rect 2 41 6 58
rect 12 50 13 54
rect 17 50 18 54
rect 12 47 18 50
rect 26 51 33 55
rect 37 51 38 55
rect 10 43 13 47
rect 17 43 23 47
rect 10 42 23 43
rect 10 31 14 42
rect 26 39 30 51
rect 2 29 14 31
rect 2 25 3 29
rect 7 25 14 29
rect 18 38 30 39
rect 22 35 30 38
rect 18 21 22 34
rect 34 31 38 47
rect 26 30 38 31
rect 26 26 29 30
rect 33 26 38 30
rect 26 25 38 26
rect 18 17 33 21
rect 37 17 38 21
rect -2 8 21 12
rect 25 8 42 12
rect -2 2 42 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
<< ntransistor >>
rect 9 18 11 30
rect 16 18 18 30
rect 28 15 30 22
<< ptransistor >>
rect 9 42 11 56
rect 19 42 21 56
rect 29 42 31 56
<< polycontact >>
rect 10 60 14 64
rect 18 34 22 38
rect 29 26 33 30
<< ndcontact >>
rect 3 25 7 29
rect 33 17 37 21
rect 21 8 25 12
<< pdcontact >>
rect 3 68 7 72
rect 22 64 26 68
rect 13 50 17 54
rect 13 43 17 47
rect 33 51 37 55
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
<< psubstratepdiff >>
rect 0 2 40 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 40 2
rect 0 -3 40 -2
<< nsubstratendiff >>
rect 0 82 40 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 40 82
rect 0 77 40 78
<< labels >>
rlabel ptransistor 20 47 20 47 6 an
rlabel ndcontact 4 28 4 28 6 z
rlabel metal1 4 52 4 52 6 b
rlabel metal1 12 36 12 36 6 z
rlabel metal1 12 60 12 60 6 b
rlabel metal1 20 6 20 6 6 vss
rlabel metal1 20 28 20 28 6 an
rlabel metal1 28 28 28 28 6 a
rlabel metal1 20 44 20 44 6 z
rlabel metal1 20 74 20 74 6 vdd
rlabel metal1 28 19 28 19 6 an
rlabel metal1 36 36 36 36 6 a
rlabel metal1 32 53 32 53 6 an
<< end >>
