.subckt xor2v2x05 a b vdd vss z
*   SPICE3 file   created from xor2v2x05.ext -      technology: scmos
m00 z      bn     an     vdd p w=16u  l=2.3636u ad=64p      pd=24u      as=92p      ps=46u
m01 bn     an     z      vdd p w=16u  l=2.3636u ad=64p      pd=24u      as=64p      ps=24u
m02 vdd    b      bn     vdd p w=16u  l=2.3636u ad=110p     pd=36u      as=64p      ps=24u
m03 an     a      vdd    vdd p w=16u  l=2.3636u ad=92p      pd=46u      as=110p     ps=36u
m04 w1     bn     z      vss n w=11u  l=2.3636u ad=27.5p    pd=16u      as=53.3704p ps=27.7037u
m05 vss    an     w1     vss n w=11u  l=2.3636u ad=99.4783p pd=44u      as=27.5p    ps=16u
m06 bn     b      vss    vss n w=6u   l=2.3636u ad=24.8571p pd=13.7143u as=54.2609p ps=24u
m07 z      a      bn     vss n w=8u   l=2.3636u ad=38.8148p pd=20.1481u as=33.1429p ps=18.2857u
m08 an     b      z      vss n w=8u   l=2.3636u ad=33.1429p pd=18.2857u as=38.8148p ps=20.1481u
m09 vss    a      an     vss n w=6u   l=2.3636u ad=54.2609p pd=24u      as=24.8571p ps=13.7143u
C0  z      b      0.009f
C1  an     bn     0.524f
C2  a      vdd    0.018f
C3  bn     b      0.041f
C4  an     vdd    0.274f
C5  b      vdd    0.084f
C6  vss    z      0.274f
C7  a      an     0.083f
C8  vss    bn     0.093f
C9  vss    vdd    0.003f
C10 z      bn     0.497f
C11 a      b      0.186f
C12 an     b      0.123f
C13 z      vdd    0.042f
C14 bn     vdd    0.047f
C15 vss    a      0.028f
C16 w1     z      0.010f
C17 vss    an     0.090f
C18 w1     bn     0.005f
C19 a      z      0.003f
C20 z      an     0.327f
C21 a      bn     0.015f
C22 vss    b      0.029f
C24 a      vss    0.040f
C25 z      vss    0.021f
C26 an     vss    0.039f
C27 bn     vss    0.029f
C28 b      vss    0.061f
.ends
