magic
tech scmos
timestamp 1179386646
<< checkpaint >>
rect -22 -25 78 105
<< ab >>
rect 0 0 56 80
<< pwell >>
rect -4 -7 60 36
<< nwell >>
rect -4 36 60 87
<< polysilicon >>
rect 9 66 11 71
rect 19 66 21 71
rect 29 66 31 71
rect 39 66 41 71
rect 9 39 11 49
rect 19 46 21 49
rect 29 46 31 49
rect 19 45 25 46
rect 19 41 20 45
rect 24 41 25 45
rect 19 40 25 41
rect 29 45 35 46
rect 29 41 30 45
rect 34 41 35 45
rect 29 40 35 41
rect 9 38 15 39
rect 9 34 10 38
rect 14 36 15 38
rect 14 34 17 36
rect 9 33 17 34
rect 15 30 17 33
rect 22 30 24 40
rect 29 30 31 40
rect 39 39 41 49
rect 39 38 47 39
rect 39 35 42 38
rect 36 34 42 35
rect 46 34 47 38
rect 36 33 47 34
rect 36 30 38 33
rect 15 6 17 10
rect 22 6 24 10
rect 29 6 31 10
rect 36 6 38 10
<< ndiffusion >>
rect 10 22 15 30
rect 8 21 15 22
rect 8 17 9 21
rect 13 17 15 21
rect 8 16 15 17
rect 10 10 15 16
rect 17 10 22 30
rect 24 10 29 30
rect 31 10 36 30
rect 38 12 47 30
rect 38 10 41 12
rect 40 8 41 10
rect 45 8 47 12
rect 40 7 47 8
<< pdiffusion >>
rect 43 72 49 73
rect 43 68 44 72
rect 48 68 49 72
rect 43 66 49 68
rect 2 65 9 66
rect 2 61 3 65
rect 7 61 9 65
rect 2 49 9 61
rect 11 62 19 66
rect 11 58 13 62
rect 17 58 19 62
rect 11 55 19 58
rect 11 51 13 55
rect 17 51 19 55
rect 11 49 19 51
rect 21 65 29 66
rect 21 61 23 65
rect 27 61 29 65
rect 21 49 29 61
rect 31 62 39 66
rect 31 58 33 62
rect 37 58 39 62
rect 31 55 39 58
rect 31 51 33 55
rect 37 51 39 55
rect 31 49 39 51
rect 41 49 49 66
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect -2 72 58 78
rect -2 68 44 72
rect 48 68 58 72
rect 3 65 7 68
rect 23 65 27 68
rect 3 60 7 61
rect 13 62 17 63
rect 23 60 27 61
rect 33 62 38 63
rect 13 55 17 58
rect 37 58 38 62
rect 33 55 38 58
rect 2 51 13 55
rect 17 51 33 55
rect 37 51 38 55
rect 2 49 14 51
rect 2 21 6 49
rect 42 47 46 63
rect 18 45 24 47
rect 18 41 20 45
rect 29 41 30 45
rect 34 43 46 47
rect 10 38 14 39
rect 10 29 14 34
rect 18 37 24 41
rect 18 33 30 37
rect 34 33 38 43
rect 42 38 46 39
rect 10 25 22 29
rect 2 17 9 21
rect 13 17 14 21
rect 18 17 22 25
rect 26 17 30 33
rect 42 23 46 34
rect 34 17 46 23
rect -2 8 41 12
rect 45 8 58 12
rect -2 2 58 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
<< ntransistor >>
rect 15 10 17 30
rect 22 10 24 30
rect 29 10 31 30
rect 36 10 38 30
<< ptransistor >>
rect 9 49 11 66
rect 19 49 21 66
rect 29 49 31 66
rect 39 49 41 66
<< polycontact >>
rect 20 41 24 45
rect 30 41 34 45
rect 10 34 14 38
rect 42 34 46 38
<< ndcontact >>
rect 9 17 13 21
rect 41 8 45 12
<< pdcontact >>
rect 44 68 48 72
rect 3 61 7 65
rect 13 58 17 62
rect 13 51 17 55
rect 23 61 27 65
rect 33 58 37 62
rect 33 51 37 55
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
<< psubstratepdiff >>
rect 0 2 56 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 56 2
rect 0 -3 56 -2
<< nsubstratendiff >>
rect 0 82 56 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 56 82
rect 0 77 56 78
<< labels >>
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 32 12 32 6 d
rlabel metal1 12 52 12 52 6 z
rlabel metal1 28 6 28 6 6 vss
rlabel metal1 20 20 20 20 6 d
rlabel metal1 28 24 28 24 6 c
rlabel metal1 20 40 20 40 6 c
rlabel metal1 28 74 28 74 6 vdd
rlabel metal1 36 20 36 20 6 a
rlabel metal1 44 28 44 28 6 a
rlabel metal1 36 40 36 40 6 b
rlabel pdcontact 36 60 36 60 6 z
rlabel metal1 44 56 44 56 6 b
<< end >>
