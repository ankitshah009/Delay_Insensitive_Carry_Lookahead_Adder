magic
tech scmos
timestamp 1179386043
<< checkpaint >>
rect -22 -25 46 105
<< ab >>
rect 0 0 24 80
<< pwell >>
rect -4 -7 28 36
<< nwell >>
rect -4 36 28 87
<< polysilicon >>
rect 9 70 11 74
rect 9 39 11 42
rect 9 38 15 39
rect 9 34 10 38
rect 14 34 15 38
rect 9 33 15 34
rect 9 30 11 33
rect 9 11 11 16
<< ndiffusion >>
rect 2 28 9 30
rect 2 24 3 28
rect 7 24 9 28
rect 2 21 9 24
rect 2 17 3 21
rect 7 17 9 21
rect 2 16 9 17
rect 11 16 20 30
rect 13 12 20 16
rect 13 8 14 12
rect 18 8 20 12
rect 13 7 20 8
<< pdiffusion >>
rect 13 72 20 73
rect 13 70 14 72
rect 4 57 9 70
rect 2 56 9 57
rect 2 52 3 56
rect 7 52 9 56
rect 2 49 9 52
rect 2 45 3 49
rect 7 45 9 49
rect 2 44 9 45
rect 4 42 9 44
rect 11 68 14 70
rect 18 68 20 72
rect 11 42 20 68
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect -2 72 26 78
rect -2 68 14 72
rect 18 68 26 72
rect 2 57 14 63
rect 2 56 7 57
rect 2 52 3 56
rect 2 49 7 52
rect 2 45 3 49
rect 2 44 7 45
rect 2 29 6 44
rect 18 39 22 63
rect 10 38 22 39
rect 14 34 22 38
rect 10 33 22 34
rect 2 28 7 29
rect 2 24 3 28
rect 2 23 7 24
rect 2 21 14 23
rect 2 17 3 21
rect 7 17 14 21
rect 18 17 22 33
rect -2 8 14 12
rect 18 8 26 12
rect -2 2 26 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
<< ntransistor >>
rect 9 16 11 30
<< ptransistor >>
rect 9 42 11 70
<< polycontact >>
rect 10 34 14 38
<< ndcontact >>
rect 3 24 7 28
rect 3 17 7 21
rect 14 8 18 12
<< pdcontact >>
rect 3 52 7 56
rect 3 45 7 49
rect 14 68 18 72
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
<< psubstratepdiff >>
rect 0 2 24 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 24 2
rect 0 -3 24 -2
<< nsubstratendiff >>
rect 0 82 24 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 24 82
rect 0 77 24 78
<< labels >>
rlabel metal1 4 40 4 40 6 z
rlabel metal1 12 6 12 6 6 vss
rlabel metal1 12 20 12 20 6 z
rlabel polycontact 12 36 12 36 6 a
rlabel metal1 12 60 12 60 6 z
rlabel metal1 12 74 12 74 6 vdd
rlabel metal1 20 40 20 40 6 a
<< end >>
