magic
tech scmos
timestamp 1179385212
<< checkpaint >>
rect -22 -22 78 94
<< ab >>
rect 0 0 56 72
<< pwell >>
rect -4 -4 60 32
<< nwell >>
rect -4 32 60 76
<< polysilicon >>
rect 12 66 14 70
rect 19 66 21 70
rect 29 66 31 70
rect 39 66 41 70
rect 12 28 14 39
rect 19 36 21 39
rect 29 36 31 39
rect 39 36 41 39
rect 19 35 25 36
rect 19 31 20 35
rect 24 31 25 35
rect 19 30 25 31
rect 29 35 35 36
rect 29 31 30 35
rect 34 31 35 35
rect 29 30 35 31
rect 39 35 47 36
rect 39 31 42 35
rect 46 31 47 35
rect 39 30 47 31
rect 9 27 15 28
rect 9 23 10 27
rect 14 23 15 27
rect 9 22 15 23
rect 10 19 12 22
rect 20 19 22 30
rect 32 22 34 30
rect 39 22 41 30
rect 10 8 12 13
rect 20 8 22 13
rect 32 8 34 13
rect 39 8 41 13
<< ndiffusion >>
rect 24 19 32 22
rect 2 13 10 19
rect 12 18 20 19
rect 12 14 14 18
rect 18 14 20 18
rect 12 13 20 14
rect 22 13 32 19
rect 34 13 39 22
rect 41 19 46 22
rect 41 18 48 19
rect 41 14 43 18
rect 47 14 48 18
rect 41 13 48 14
rect 2 8 8 13
rect 24 8 30 13
rect 2 4 3 8
rect 7 4 8 8
rect 2 3 8 4
rect 24 4 25 8
rect 29 4 30 8
rect 24 3 30 4
<< pdiffusion >>
rect 7 60 12 66
rect 5 59 12 60
rect 5 55 6 59
rect 10 55 12 59
rect 5 51 12 55
rect 5 47 6 51
rect 10 47 12 51
rect 5 46 12 47
rect 7 39 12 46
rect 14 39 19 66
rect 21 58 29 66
rect 21 54 23 58
rect 27 54 29 58
rect 21 39 29 54
rect 31 65 39 66
rect 31 61 33 65
rect 37 61 39 65
rect 31 39 39 61
rect 41 59 46 66
rect 41 58 48 59
rect 41 54 43 58
rect 47 54 48 58
rect 41 53 48 54
rect 41 39 46 53
<< metal1 >>
rect -2 65 58 72
rect -2 64 33 65
rect 32 61 33 64
rect 37 64 58 65
rect 37 61 38 64
rect 2 18 6 59
rect 10 55 11 59
rect 22 54 23 58
rect 27 54 43 58
rect 47 54 48 58
rect 10 47 11 51
rect 18 45 30 51
rect 34 45 46 51
rect 10 27 14 43
rect 18 37 24 45
rect 20 35 24 37
rect 42 35 46 45
rect 29 31 30 35
rect 34 31 38 35
rect 20 30 24 31
rect 33 26 38 31
rect 42 30 46 31
rect 14 23 23 26
rect 10 22 23 23
rect 33 22 47 26
rect 2 14 14 18
rect 18 14 43 18
rect 47 14 48 18
rect -2 4 3 8
rect 7 4 25 8
rect 29 4 48 8
rect 52 4 58 8
rect -2 0 58 4
<< ntransistor >>
rect 10 13 12 19
rect 20 13 22 19
rect 32 13 34 22
rect 39 13 41 22
<< ptransistor >>
rect 12 39 14 66
rect 19 39 21 66
rect 29 39 31 66
rect 39 39 41 66
<< polycontact >>
rect 20 31 24 35
rect 30 31 34 35
rect 42 31 46 35
rect 10 23 14 27
<< ndcontact >>
rect 14 14 18 18
rect 43 14 47 18
rect 3 4 7 8
rect 25 4 29 8
<< pdcontact >>
rect 6 55 10 59
rect 6 47 10 51
rect 23 54 27 58
rect 33 61 37 65
rect 43 54 47 58
<< psubstratepcontact >>
rect 48 4 52 8
<< psubstratepdiff >>
rect 47 8 53 9
rect 47 4 48 8
rect 52 4 53 8
rect 47 3 53 4
<< labels >>
rlabel metal1 4 40 4 40 6 z
rlabel metal1 20 16 20 16 6 z
rlabel metal1 12 16 12 16 6 z
rlabel metal1 20 24 20 24 6 c
rlabel metal1 12 36 12 36 6 c
rlabel metal1 20 44 20 44 6 b
rlabel metal1 28 4 28 4 6 vss
rlabel metal1 36 16 36 16 6 z
rlabel metal1 28 16 28 16 6 z
rlabel metal1 36 28 36 28 6 a1
rlabel metal1 28 48 28 48 6 b
rlabel metal1 36 48 36 48 6 a2
rlabel metal1 28 68 28 68 6 vdd
rlabel ndcontact 44 16 44 16 6 z
rlabel metal1 44 24 44 24 6 a1
rlabel metal1 44 44 44 44 6 a2
rlabel metal1 35 56 35 56 6 n1
<< end >>
