magic
tech scmos
timestamp 1179384971
<< checkpaint >>
rect -22 -25 62 105
<< ab >>
rect 0 0 40 80
<< pwell >>
rect -4 -7 44 36
<< nwell >>
rect -4 36 44 87
<< polysilicon >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 9 39 11 42
rect 19 39 21 51
rect 29 47 31 51
rect 29 46 35 47
rect 29 42 30 46
rect 34 42 35 46
rect 29 41 35 42
rect 9 38 15 39
rect 9 34 10 38
rect 14 34 15 38
rect 9 33 15 34
rect 19 38 25 39
rect 19 34 20 38
rect 24 34 25 38
rect 19 33 25 34
rect 9 30 11 33
rect 22 30 24 33
rect 29 30 31 41
rect 9 11 11 16
rect 22 12 24 17
rect 29 12 31 17
<< ndiffusion >>
rect 2 29 9 30
rect 2 25 3 29
rect 7 25 9 29
rect 2 21 9 25
rect 2 17 3 21
rect 7 17 9 21
rect 2 16 9 17
rect 11 17 22 30
rect 24 17 29 30
rect 31 23 36 30
rect 31 22 38 23
rect 31 18 33 22
rect 37 18 38 22
rect 31 17 38 18
rect 11 16 20 17
rect 13 12 20 16
rect 13 8 14 12
rect 18 8 20 12
rect 13 7 20 8
<< pdiffusion >>
rect 4 63 9 70
rect 2 62 9 63
rect 2 58 3 62
rect 7 58 9 62
rect 2 55 9 58
rect 2 51 3 55
rect 7 51 9 55
rect 2 50 9 51
rect 4 42 9 50
rect 11 69 19 70
rect 11 65 13 69
rect 17 65 19 69
rect 11 62 19 65
rect 11 58 13 62
rect 17 58 19 62
rect 11 51 19 58
rect 21 63 29 70
rect 21 59 23 63
rect 27 59 29 63
rect 21 56 29 59
rect 21 52 23 56
rect 27 52 29 56
rect 21 51 29 52
rect 31 69 38 70
rect 31 65 33 69
rect 37 65 38 69
rect 31 62 38 65
rect 31 58 33 62
rect 37 58 38 62
rect 31 51 38 58
rect 11 42 17 51
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect -2 69 42 78
rect -2 68 13 69
rect 12 65 13 68
rect 17 68 33 69
rect 17 65 18 68
rect 2 62 7 63
rect 2 58 3 62
rect 12 62 18 65
rect 32 65 33 68
rect 37 68 42 69
rect 37 65 38 68
rect 12 58 13 62
rect 17 58 18 62
rect 23 63 27 64
rect 2 55 7 58
rect 2 51 3 55
rect 23 56 27 59
rect 32 62 38 65
rect 32 58 33 62
rect 37 58 38 62
rect 2 50 7 51
rect 14 52 23 54
rect 14 50 27 52
rect 2 30 6 50
rect 14 46 18 50
rect 10 42 18 46
rect 25 42 30 46
rect 34 42 38 55
rect 10 38 14 42
rect 17 34 20 38
rect 24 34 31 38
rect 10 30 14 34
rect 2 29 7 30
rect 2 25 3 29
rect 10 26 22 30
rect 2 23 7 25
rect 2 21 14 23
rect 2 17 3 21
rect 7 17 14 21
rect 18 22 22 26
rect 26 25 31 34
rect 18 18 33 22
rect 37 18 38 22
rect -2 8 14 12
rect 18 8 42 12
rect -2 2 42 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
<< ntransistor >>
rect 9 16 11 30
rect 22 17 24 30
rect 29 17 31 30
<< ptransistor >>
rect 9 42 11 70
rect 19 51 21 70
rect 29 51 31 70
<< polycontact >>
rect 30 42 34 46
rect 10 34 14 38
rect 20 34 24 38
<< ndcontact >>
rect 3 25 7 29
rect 3 17 7 21
rect 33 18 37 22
rect 14 8 18 12
<< pdcontact >>
rect 3 58 7 62
rect 3 51 7 55
rect 13 65 17 69
rect 13 58 17 62
rect 23 59 27 63
rect 23 52 27 56
rect 33 65 37 69
rect 33 58 37 62
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
<< psubstratepdiff >>
rect 0 2 40 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 40 2
rect 0 -3 40 -2
<< nsubstratendiff >>
rect 0 82 40 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 40 82
rect 0 77 40 78
<< labels >>
rlabel polycontact 12 36 12 36 6 zn
rlabel metal1 4 40 4 40 6 z
rlabel metal1 12 20 12 20 6 z
rlabel polycontact 12 36 12 36 6 zn
rlabel metal1 20 6 20 6 6 vss
rlabel metal1 20 36 20 36 6 a
rlabel metal1 28 32 28 32 6 a
rlabel metal1 28 44 28 44 6 b
rlabel metal1 25 57 25 57 6 zn
rlabel metal1 20 74 20 74 6 vdd
rlabel metal1 28 20 28 20 6 zn
rlabel metal1 36 52 36 52 6 b
<< end >>
