magic
tech scmos
timestamp 1179387142
<< checkpaint >>
rect -22 -22 86 94
<< ab >>
rect 0 0 64 72
<< pwell >>
rect -4 -4 68 32
<< nwell >>
rect -4 32 68 76
<< polysilicon >>
rect 39 65 41 70
rect 46 65 48 70
rect 29 58 31 63
rect 9 50 11 55
rect 29 43 31 50
rect 29 42 35 43
rect 29 38 30 42
rect 34 38 35 42
rect 9 35 11 38
rect 29 37 35 38
rect 9 34 18 35
rect 9 30 13 34
rect 17 30 18 34
rect 9 29 18 30
rect 9 26 11 29
rect 29 26 31 37
rect 39 35 41 50
rect 46 43 48 50
rect 46 42 57 43
rect 46 41 52 42
rect 51 38 52 41
rect 56 38 57 42
rect 51 37 57 38
rect 39 34 47 35
rect 39 30 42 34
rect 46 30 47 34
rect 39 29 47 30
rect 39 26 41 29
rect 9 15 11 20
rect 51 19 53 37
rect 29 14 31 19
rect 39 14 41 19
rect 51 7 53 12
<< ndiffusion >>
rect 2 25 9 26
rect 2 21 3 25
rect 7 21 9 25
rect 2 20 9 21
rect 11 25 18 26
rect 11 21 13 25
rect 17 21 18 25
rect 11 20 18 21
rect 22 25 29 26
rect 22 21 23 25
rect 27 21 29 25
rect 22 19 29 21
rect 31 24 39 26
rect 31 20 33 24
rect 37 20 39 24
rect 31 19 39 20
rect 41 19 49 26
rect 43 12 51 19
rect 53 17 60 19
rect 53 13 55 17
rect 59 13 60 17
rect 53 12 60 13
rect 43 8 49 12
rect 43 4 44 8
rect 48 4 49 8
rect 43 3 49 4
<< pdiffusion >>
rect 13 59 27 60
rect 13 55 14 59
rect 18 58 27 59
rect 34 58 39 65
rect 18 55 29 58
rect 13 51 29 55
rect 13 50 14 51
rect 4 44 9 50
rect 2 43 9 44
rect 2 39 3 43
rect 7 39 9 43
rect 2 38 9 39
rect 11 47 14 50
rect 18 50 29 51
rect 31 57 39 58
rect 31 53 33 57
rect 37 53 39 57
rect 31 50 39 53
rect 41 50 46 65
rect 48 64 56 65
rect 48 60 50 64
rect 54 60 56 64
rect 48 57 56 60
rect 48 53 50 57
rect 54 53 56 57
rect 48 50 56 53
rect 18 47 27 50
rect 11 38 27 47
<< metal1 >>
rect -2 68 66 72
rect -2 64 4 68
rect 8 64 66 68
rect 13 59 19 64
rect 13 55 14 59
rect 18 55 19 59
rect 50 57 54 60
rect 13 51 19 55
rect 13 47 14 51
rect 18 47 19 51
rect 23 53 33 57
rect 37 53 38 57
rect 2 39 3 43
rect 7 39 15 43
rect 2 38 15 39
rect 2 26 6 38
rect 23 34 27 53
rect 50 52 54 53
rect 42 46 46 51
rect 34 43 46 46
rect 30 42 46 43
rect 50 42 62 43
rect 34 38 38 42
rect 30 37 38 38
rect 50 38 52 42
rect 56 38 62 42
rect 50 37 62 38
rect 12 30 13 34
rect 17 30 27 34
rect 2 25 7 26
rect 2 21 3 25
rect 2 20 7 21
rect 13 25 17 26
rect 2 13 6 20
rect 13 8 17 21
rect 23 25 27 30
rect 42 34 46 35
rect 42 27 46 30
rect 58 29 62 37
rect 23 20 27 21
rect 33 24 37 25
rect 42 21 54 27
rect 33 17 37 20
rect 33 13 55 17
rect 59 13 60 17
rect -2 4 4 8
rect 8 4 12 8
rect 16 4 44 8
rect 48 4 66 8
rect -2 0 66 4
<< ntransistor >>
rect 9 20 11 26
rect 29 19 31 26
rect 39 19 41 26
rect 51 12 53 19
<< ptransistor >>
rect 9 38 11 50
rect 29 50 31 58
rect 39 50 41 65
rect 46 50 48 65
<< polycontact >>
rect 30 38 34 42
rect 13 30 17 34
rect 52 38 56 42
rect 42 30 46 34
<< ndcontact >>
rect 3 21 7 25
rect 13 21 17 25
rect 23 21 27 25
rect 33 20 37 24
rect 55 13 59 17
rect 44 4 48 8
<< pdcontact >>
rect 14 55 18 59
rect 3 39 7 43
rect 14 47 18 51
rect 33 53 37 57
rect 50 60 54 64
rect 50 53 54 57
<< psubstratepcontact >>
rect 4 4 8 8
rect 12 4 16 8
<< nsubstratencontact >>
rect 4 64 8 68
<< psubstratepdiff >>
rect 3 8 17 9
rect 3 4 4 8
rect 8 4 12 8
rect 16 4 17 8
rect 3 3 17 4
<< nsubstratendiff >>
rect 3 68 9 69
rect 3 64 4 68
rect 8 64 9 68
rect 3 57 9 64
<< labels >>
rlabel polysilicon 13 32 13 32 6 zn
rlabel metal1 4 28 4 28 6 z
rlabel metal1 12 40 12 40 6 z
rlabel metal1 19 32 19 32 6 zn
rlabel metal1 25 38 25 38 6 zn
rlabel metal1 32 4 32 4 6 vss
rlabel metal1 35 19 35 19 6 n1
rlabel metal1 44 28 44 28 6 a2
rlabel metal1 36 40 36 40 6 b
rlabel metal1 44 48 44 48 6 b
rlabel metal1 30 55 30 55 6 zn
rlabel metal1 32 68 32 68 6 vdd
rlabel metal1 46 15 46 15 6 n1
rlabel metal1 52 24 52 24 6 a2
rlabel metal1 60 36 60 36 6 a1
rlabel metal1 52 40 52 40 6 a1
<< end >>
