magic
tech scmos
timestamp 1185038996
<< checkpaint >>
rect -22 -24 102 124
<< ab >>
rect 0 0 80 100
<< pwell >>
rect -2 -4 82 49
<< nwell >>
rect -2 49 82 104
<< polysilicon >>
rect 45 95 47 98
rect 57 95 59 98
rect 11 83 13 86
rect 23 83 25 86
rect 35 83 37 86
rect 11 43 13 63
rect 23 53 25 63
rect 17 52 25 53
rect 17 48 18 52
rect 22 48 25 52
rect 17 47 25 48
rect 7 42 15 43
rect 7 38 8 42
rect 12 38 15 42
rect 7 37 15 38
rect 13 35 15 37
rect 21 35 23 47
rect 35 43 37 63
rect 67 82 73 83
rect 67 78 68 82
rect 72 78 73 82
rect 67 77 73 78
rect 67 75 69 77
rect 45 43 47 55
rect 57 43 59 55
rect 27 42 37 43
rect 27 38 28 42
rect 32 41 37 42
rect 43 42 63 43
rect 32 38 33 41
rect 27 37 33 38
rect 43 38 58 42
rect 62 38 63 42
rect 43 37 63 38
rect 29 35 31 37
rect 43 25 45 37
rect 55 25 57 37
rect 67 25 69 55
rect 13 12 15 15
rect 21 12 23 15
rect 29 12 31 15
rect 67 12 69 15
rect 43 2 45 5
rect 55 2 57 5
<< ndiffusion >>
rect 5 22 13 35
rect 5 18 6 22
rect 10 18 13 22
rect 5 15 13 18
rect 15 15 21 35
rect 23 15 29 35
rect 31 25 41 35
rect 31 15 43 25
rect 33 12 43 15
rect 33 8 36 12
rect 40 8 43 12
rect 33 5 43 8
rect 45 22 55 25
rect 45 18 48 22
rect 52 18 55 22
rect 45 5 55 18
rect 57 15 67 25
rect 69 22 77 25
rect 69 18 72 22
rect 76 18 77 22
rect 69 15 77 18
rect 57 12 65 15
rect 57 8 60 12
rect 64 8 65 12
rect 57 5 65 8
<< pdiffusion >>
rect 37 94 45 95
rect 15 92 21 93
rect 15 88 16 92
rect 20 88 21 92
rect 37 90 38 94
rect 42 90 45 94
rect 37 89 45 90
rect 15 83 21 88
rect 39 83 45 89
rect 3 82 11 83
rect 3 78 4 82
rect 8 78 11 82
rect 3 63 11 78
rect 13 63 23 83
rect 25 82 35 83
rect 25 78 28 82
rect 32 78 35 82
rect 25 63 35 78
rect 37 63 45 83
rect 39 55 45 63
rect 47 72 57 95
rect 47 68 50 72
rect 54 68 57 72
rect 47 62 57 68
rect 47 58 50 62
rect 54 58 57 62
rect 47 55 57 58
rect 59 94 67 95
rect 59 90 62 94
rect 66 90 67 94
rect 59 89 67 90
rect 59 75 65 89
rect 59 55 67 75
rect 69 72 77 75
rect 69 68 72 72
rect 76 68 77 72
rect 69 62 77 68
rect 69 58 72 62
rect 76 58 77 62
rect 69 55 77 58
<< metal1 >>
rect -2 94 82 101
rect -2 92 38 94
rect -2 88 16 92
rect 20 90 38 92
rect 42 90 62 94
rect 66 90 82 94
rect 20 88 82 90
rect -2 87 82 88
rect 3 82 9 83
rect 27 82 33 83
rect 67 82 73 83
rect 3 78 4 82
rect 8 78 28 82
rect 32 78 68 82
rect 72 78 73 82
rect 3 77 9 78
rect 27 77 33 78
rect 7 42 13 72
rect 7 38 8 42
rect 12 38 13 42
rect 7 28 13 38
rect 17 52 23 72
rect 17 48 18 52
rect 22 48 23 52
rect 17 28 23 48
rect 27 42 33 72
rect 27 38 28 42
rect 32 38 33 42
rect 27 28 33 38
rect 5 22 11 23
rect 38 22 42 78
rect 67 77 73 78
rect 5 18 6 22
rect 10 18 42 22
rect 47 72 55 73
rect 47 68 50 72
rect 54 68 55 72
rect 47 67 55 68
rect 71 72 77 73
rect 71 68 72 72
rect 76 68 77 72
rect 71 67 77 68
rect 47 63 53 67
rect 72 63 76 67
rect 47 62 55 63
rect 47 58 50 62
rect 54 58 55 62
rect 47 57 55 58
rect 71 62 77 63
rect 71 58 72 62
rect 76 58 77 62
rect 71 57 77 58
rect 47 22 53 57
rect 57 42 63 43
rect 72 42 76 57
rect 57 38 58 42
rect 62 38 76 42
rect 57 37 63 38
rect 72 23 76 38
rect 47 18 48 22
rect 52 18 53 22
rect 5 17 11 18
rect 47 17 53 18
rect 71 22 77 23
rect 71 18 72 22
rect 76 18 77 22
rect 71 17 77 18
rect -2 12 82 13
rect -2 8 36 12
rect 40 8 60 12
rect 64 8 82 12
rect -2 4 4 8
rect 8 4 12 8
rect 16 4 20 8
rect 24 4 82 8
rect -2 -1 82 4
<< ntransistor >>
rect 13 15 15 35
rect 21 15 23 35
rect 29 15 31 35
rect 43 5 45 25
rect 55 5 57 25
rect 67 15 69 25
<< ptransistor >>
rect 11 63 13 83
rect 23 63 25 83
rect 35 63 37 83
rect 45 55 47 95
rect 57 55 59 95
rect 67 55 69 75
<< polycontact >>
rect 18 48 22 52
rect 8 38 12 42
rect 68 78 72 82
rect 28 38 32 42
rect 58 38 62 42
<< ndcontact >>
rect 6 18 10 22
rect 36 8 40 12
rect 48 18 52 22
rect 72 18 76 22
rect 60 8 64 12
<< pdcontact >>
rect 16 88 20 92
rect 38 90 42 94
rect 4 78 8 82
rect 28 78 32 82
rect 50 68 54 72
rect 50 58 54 62
rect 62 90 66 94
rect 72 68 76 72
rect 72 58 76 62
<< psubstratepcontact >>
rect 4 4 8 8
rect 12 4 16 8
rect 20 4 24 8
<< psubstratepdiff >>
rect 3 8 25 9
rect 3 4 4 8
rect 8 4 12 8
rect 16 4 20 8
rect 24 4 25 8
rect 3 3 25 4
<< labels >>
rlabel metal1 10 50 10 50 6 i0
rlabel metal1 10 50 10 50 6 i0
rlabel metal1 30 50 30 50 6 i1
rlabel metal1 30 50 30 50 6 i1
rlabel polycontact 20 50 20 50 6 i2
rlabel polycontact 20 50 20 50 6 i2
rlabel metal1 40 6 40 6 6 vss
rlabel metal1 40 6 40 6 6 vss
rlabel metal1 50 45 50 45 6 nq
rlabel metal1 50 45 50 45 6 nq
rlabel metal1 40 94 40 94 6 vdd
rlabel metal1 40 94 40 94 6 vdd
<< end >>
