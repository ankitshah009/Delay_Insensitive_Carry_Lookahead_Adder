magic
tech scmos
timestamp 1180600636
<< checkpaint >>
rect -22 -22 62 122
<< ab >>
rect 0 0 40 100
<< pwell >>
rect -4 -4 44 48
<< nwell >>
rect -4 48 44 104
<< polysilicon >>
rect 23 94 25 98
rect 11 68 13 72
rect 11 53 13 56
rect 11 52 19 53
rect 11 48 14 52
rect 18 48 19 52
rect 11 47 19 48
rect 3 42 9 43
rect 23 42 25 55
rect 3 38 4 42
rect 8 38 25 42
rect 3 37 9 38
rect 11 32 19 33
rect 11 28 14 32
rect 18 28 19 32
rect 11 27 19 28
rect 11 24 13 27
rect 23 25 25 38
rect 11 14 13 18
rect 23 2 25 6
<< ndiffusion >>
rect 3 24 9 25
rect 18 24 23 25
rect 3 20 4 24
rect 8 20 11 24
rect 3 18 11 20
rect 13 18 23 24
rect 15 12 23 18
rect 15 8 16 12
rect 20 8 23 12
rect 15 6 23 8
rect 25 22 33 25
rect 25 18 28 22
rect 32 18 33 22
rect 25 6 33 18
<< pdiffusion >>
rect 15 92 23 94
rect 15 88 16 92
rect 20 88 23 92
rect 15 68 23 88
rect 3 62 11 68
rect 3 58 4 62
rect 8 58 11 62
rect 3 56 11 58
rect 13 56 23 68
rect 18 55 23 56
rect 25 82 33 94
rect 25 78 28 82
rect 32 78 33 82
rect 25 72 33 78
rect 25 68 28 72
rect 32 68 33 72
rect 25 62 33 68
rect 25 58 28 62
rect 32 58 33 62
rect 25 55 33 58
<< metal1 >>
rect -2 96 42 100
rect -2 92 4 96
rect 8 92 42 96
rect -2 88 16 92
rect 20 88 42 92
rect 4 86 8 88
rect 4 81 8 82
rect 4 62 8 63
rect 4 42 8 58
rect 13 48 14 52
rect 4 24 8 38
rect 13 28 14 32
rect 4 19 8 20
rect 18 17 22 83
rect 28 82 32 83
rect 28 72 32 78
rect 28 62 32 68
rect 28 22 32 58
rect 28 17 32 18
rect -2 8 16 12
rect 20 8 42 12
rect -2 0 42 8
<< ntransistor >>
rect 11 18 13 24
rect 23 6 25 25
<< ptransistor >>
rect 11 56 13 68
rect 23 55 25 94
<< polycontact >>
rect 14 48 18 52
rect 4 38 8 42
rect 14 28 18 32
<< ndcontact >>
rect 4 20 8 24
rect 16 8 20 12
rect 28 18 32 22
<< pdcontact >>
rect 16 88 20 92
rect 4 58 8 62
rect 28 78 32 82
rect 28 68 32 72
rect 28 58 32 62
<< nsubstratencontact >>
rect 4 92 8 96
rect 4 82 8 86
<< nsubstratendiff >>
rect 3 96 9 97
rect 3 92 4 96
rect 8 92 9 96
rect 3 86 9 92
rect 3 82 4 86
rect 8 82 9 86
rect 3 81 9 82
<< labels >>
rlabel metal1 20 6 20 6 6 vss
rlabel metal1 20 50 20 50 6 i
rlabel metal1 20 94 20 94 6 vdd
rlabel metal1 30 50 30 50 6 q
<< end >>
