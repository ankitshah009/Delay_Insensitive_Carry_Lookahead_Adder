magic
tech scmos
timestamp 1179386753
<< checkpaint >>
rect -22 -25 86 105
<< ab >>
rect 0 0 64 80
<< pwell >>
rect -4 -7 68 36
<< nwell >>
rect -4 36 68 87
<< polysilicon >>
rect 9 70 11 74
rect 16 70 18 74
rect 26 70 28 74
rect 33 70 35 74
rect 43 70 45 74
rect 50 70 52 74
rect 9 33 11 42
rect 16 39 18 42
rect 26 39 28 42
rect 16 38 28 39
rect 16 37 23 38
rect 22 34 23 37
rect 27 34 28 38
rect 22 33 28 34
rect 33 39 35 42
rect 43 39 45 42
rect 50 39 52 42
rect 33 38 45 39
rect 33 34 34 38
rect 38 37 45 38
rect 49 38 55 39
rect 38 34 39 37
rect 33 33 39 34
rect 49 34 50 38
rect 54 34 55 38
rect 49 33 55 34
rect 9 32 15 33
rect 9 28 10 32
rect 14 28 15 32
rect 23 28 25 33
rect 35 28 37 33
rect 49 29 51 33
rect 9 27 15 28
rect 13 24 15 27
rect 45 27 51 29
rect 45 24 47 27
rect 35 12 37 17
rect 45 12 47 17
rect 13 6 15 11
rect 23 6 25 11
<< ndiffusion >>
rect 18 24 23 28
rect 4 12 13 24
rect 4 8 6 12
rect 10 11 13 12
rect 15 22 23 24
rect 15 18 17 22
rect 21 18 23 22
rect 15 11 23 18
rect 25 17 35 28
rect 37 24 42 28
rect 37 22 45 24
rect 37 18 39 22
rect 43 18 45 22
rect 37 17 45 18
rect 47 22 55 24
rect 47 18 49 22
rect 53 18 55 22
rect 47 17 55 18
rect 25 12 33 17
rect 25 11 28 12
rect 10 8 11 11
rect 4 7 11 8
rect 27 8 28 11
rect 32 8 33 12
rect 27 7 33 8
<< pdiffusion >>
rect 4 55 9 70
rect 2 54 9 55
rect 2 50 3 54
rect 7 50 9 54
rect 2 47 9 50
rect 2 43 3 47
rect 7 43 9 47
rect 2 42 9 43
rect 11 42 16 70
rect 18 69 26 70
rect 18 65 20 69
rect 24 65 26 69
rect 18 62 26 65
rect 18 58 20 62
rect 24 58 26 62
rect 18 42 26 58
rect 28 42 33 70
rect 35 62 43 70
rect 35 58 37 62
rect 41 58 43 62
rect 35 55 43 58
rect 35 51 37 55
rect 41 51 43 55
rect 35 42 43 51
rect 45 42 50 70
rect 52 69 60 70
rect 52 65 54 69
rect 58 65 60 69
rect 52 62 60 65
rect 52 58 54 62
rect 58 58 60 62
rect 52 42 60 58
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect -2 69 66 78
rect -2 68 20 69
rect 19 65 20 68
rect 24 68 54 69
rect 24 65 25 68
rect 19 62 25 65
rect 53 65 54 68
rect 58 68 66 69
rect 58 65 59 68
rect 19 58 20 62
rect 24 58 25 62
rect 37 62 41 63
rect 53 62 59 65
rect 53 58 54 62
rect 58 58 59 62
rect 37 55 41 58
rect 2 50 3 54
rect 7 51 37 54
rect 7 50 41 51
rect 2 47 7 50
rect 2 43 3 47
rect 2 42 7 43
rect 22 42 55 46
rect 2 22 6 42
rect 22 38 28 42
rect 49 38 55 42
rect 22 34 23 38
rect 27 34 28 38
rect 33 34 34 38
rect 38 34 39 38
rect 49 34 50 38
rect 54 34 55 38
rect 10 32 14 33
rect 33 30 39 34
rect 14 28 39 30
rect 10 26 39 28
rect 49 22 53 23
rect 2 18 17 22
rect 21 18 39 22
rect 43 18 44 22
rect 49 12 53 18
rect -2 8 6 12
rect 10 8 28 12
rect 32 8 66 12
rect -2 2 66 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
<< ntransistor >>
rect 13 11 15 24
rect 23 11 25 28
rect 35 17 37 28
rect 45 17 47 24
<< ptransistor >>
rect 9 42 11 70
rect 16 42 18 70
rect 26 42 28 70
rect 33 42 35 70
rect 43 42 45 70
rect 50 42 52 70
<< polycontact >>
rect 23 34 27 38
rect 34 34 38 38
rect 50 34 54 38
rect 10 28 14 32
<< ndcontact >>
rect 6 8 10 12
rect 17 18 21 22
rect 39 18 43 22
rect 49 18 53 22
rect 28 8 32 12
<< pdcontact >>
rect 3 50 7 54
rect 3 43 7 47
rect 20 65 24 69
rect 20 58 24 62
rect 37 58 41 62
rect 37 51 41 55
rect 54 65 58 69
rect 54 58 58 62
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
<< psubstratepdiff >>
rect 0 2 64 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 64 2
rect 0 -3 64 -2
<< nsubstratendiff >>
rect 0 82 64 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 64 82
rect 0 77 64 78
<< labels >>
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 20 12 20 6 z
rlabel metal1 20 28 20 28 6 b
rlabel ndcontact 20 20 20 20 6 z
rlabel metal1 20 52 20 52 6 z
rlabel metal1 12 52 12 52 6 z
rlabel metal1 32 6 32 6 6 vss
rlabel metal1 28 20 28 20 6 z
rlabel metal1 28 28 28 28 6 b
rlabel metal1 36 20 36 20 6 z
rlabel metal1 36 32 36 32 6 b
rlabel metal1 28 44 28 44 6 a
rlabel metal1 36 44 36 44 6 a
rlabel metal1 36 52 36 52 6 z
rlabel metal1 28 52 28 52 6 z
rlabel metal1 32 74 32 74 6 vdd
rlabel metal1 44 44 44 44 6 a
rlabel metal1 52 40 52 40 6 a
<< end >>
