magic
tech scmos
timestamp 1179386434
<< checkpaint >>
rect -22 -22 134 94
<< ab >>
rect 0 0 112 72
<< pwell >>
rect -4 -4 116 32
<< nwell >>
rect -4 32 116 76
<< polysilicon >>
rect 9 66 11 70
rect 19 66 21 70
rect 29 66 31 70
rect 39 66 41 70
rect 49 66 51 70
rect 59 66 61 70
rect 69 66 71 70
rect 79 66 81 70
rect 90 56 92 61
rect 100 56 102 61
rect 9 35 11 39
rect 19 35 21 39
rect 29 35 31 39
rect 39 35 41 39
rect 49 35 51 39
rect 59 35 61 39
rect 69 35 71 39
rect 9 34 15 35
rect 9 30 10 34
rect 14 30 15 34
rect 9 29 15 30
rect 19 34 33 35
rect 19 30 26 34
rect 30 30 33 34
rect 19 29 33 30
rect 12 26 14 29
rect 19 26 21 29
rect 31 26 33 29
rect 38 34 51 35
rect 38 30 42 34
rect 46 30 51 34
rect 38 29 51 30
rect 55 34 71 35
rect 55 30 58 34
rect 62 33 71 34
rect 79 35 81 39
rect 90 35 92 39
rect 100 35 102 39
rect 79 34 92 35
rect 79 33 82 34
rect 62 30 63 33
rect 55 29 63 30
rect 81 30 82 33
rect 86 33 92 34
rect 96 34 102 35
rect 86 30 87 33
rect 81 29 87 30
rect 96 30 97 34
rect 101 30 102 34
rect 96 29 102 30
rect 38 26 40 29
rect 48 26 50 29
rect 55 26 57 29
rect 12 7 14 12
rect 19 7 21 12
rect 31 2 33 7
rect 38 2 40 7
rect 48 2 50 7
rect 55 2 57 7
<< ndiffusion >>
rect 5 25 12 26
rect 5 21 6 25
rect 10 21 12 25
rect 5 18 12 21
rect 5 14 6 18
rect 10 14 12 18
rect 5 12 12 14
rect 14 12 19 26
rect 21 12 31 26
rect 23 8 31 12
rect 23 4 24 8
rect 28 7 31 8
rect 33 7 38 26
rect 40 18 48 26
rect 40 14 42 18
rect 46 14 48 18
rect 40 7 48 14
rect 50 7 55 26
rect 57 8 66 26
rect 57 7 60 8
rect 28 4 29 7
rect 23 3 29 4
rect 59 4 60 7
rect 64 4 66 8
rect 59 3 66 4
<< pdiffusion >>
rect 2 65 9 66
rect 2 61 3 65
rect 7 61 9 65
rect 2 58 9 61
rect 2 54 3 58
rect 7 54 9 58
rect 2 39 9 54
rect 11 57 19 66
rect 11 53 13 57
rect 17 53 19 57
rect 11 50 19 53
rect 11 46 13 50
rect 17 46 19 50
rect 11 39 19 46
rect 21 65 29 66
rect 21 61 23 65
rect 27 61 29 65
rect 21 58 29 61
rect 21 54 23 58
rect 27 54 29 58
rect 21 39 29 54
rect 31 58 39 66
rect 31 54 33 58
rect 37 54 39 58
rect 31 50 39 54
rect 31 46 33 50
rect 37 46 39 50
rect 31 39 39 46
rect 41 65 49 66
rect 41 61 43 65
rect 47 61 49 65
rect 41 58 49 61
rect 41 54 43 58
rect 47 54 49 58
rect 41 39 49 54
rect 51 57 59 66
rect 51 53 53 57
rect 57 53 59 57
rect 51 50 59 53
rect 51 46 53 50
rect 57 46 59 50
rect 51 39 59 46
rect 61 65 69 66
rect 61 61 63 65
rect 67 61 69 65
rect 61 58 69 61
rect 61 54 63 58
rect 67 54 69 58
rect 61 39 69 54
rect 71 58 79 66
rect 71 54 73 58
rect 77 54 79 58
rect 71 50 79 54
rect 71 46 73 50
rect 77 46 79 50
rect 71 39 79 46
rect 81 65 88 66
rect 81 61 83 65
rect 87 61 88 65
rect 81 58 88 61
rect 81 54 83 58
rect 87 56 88 58
rect 87 54 90 56
rect 81 39 90 54
rect 92 50 100 56
rect 92 46 94 50
rect 98 46 100 50
rect 92 39 100 46
rect 102 55 110 56
rect 102 51 104 55
rect 108 51 110 55
rect 102 47 110 51
rect 102 43 104 47
rect 108 43 110 47
rect 102 39 110 43
<< metal1 >>
rect -2 68 114 72
rect -2 65 96 68
rect -2 64 3 65
rect 2 61 3 64
rect 7 64 23 65
rect 7 61 8 64
rect 2 58 8 61
rect 22 61 23 64
rect 27 64 43 65
rect 27 61 28 64
rect 22 58 28 61
rect 42 61 43 64
rect 47 64 63 65
rect 47 61 48 64
rect 2 54 3 58
rect 7 54 8 58
rect 13 57 17 58
rect 22 54 23 58
rect 27 54 28 58
rect 33 58 38 59
rect 37 54 38 58
rect 42 58 48 61
rect 62 61 63 64
rect 67 64 83 65
rect 67 61 68 64
rect 62 58 68 61
rect 82 61 83 64
rect 87 64 96 65
rect 100 64 104 68
rect 108 64 114 68
rect 87 61 88 64
rect 42 54 43 58
rect 47 54 48 58
rect 53 57 57 58
rect 13 50 17 53
rect 33 50 38 54
rect 62 54 63 58
rect 67 54 68 58
rect 73 58 78 59
rect 77 54 78 58
rect 82 58 88 61
rect 82 54 83 58
rect 87 54 88 58
rect 104 55 108 64
rect 53 50 57 53
rect 73 50 78 54
rect 2 46 13 50
rect 17 46 33 50
rect 37 46 53 50
rect 57 46 73 50
rect 77 46 94 50
rect 98 46 99 50
rect 104 47 108 51
rect 2 21 6 46
rect 104 42 108 43
rect 25 38 97 42
rect 10 34 20 35
rect 14 30 20 34
rect 25 34 31 38
rect 57 34 63 38
rect 25 30 26 34
rect 30 30 31 34
rect 41 30 42 34
rect 46 30 47 34
rect 57 30 58 34
rect 62 30 63 34
rect 81 30 82 34
rect 86 30 87 34
rect 93 30 97 38
rect 101 30 103 34
rect 10 29 20 30
rect 16 26 20 29
rect 41 26 47 30
rect 81 26 87 30
rect 10 21 11 25
rect 16 22 87 26
rect 5 18 11 21
rect 5 14 6 18
rect 10 14 42 18
rect 46 14 47 18
rect -2 4 24 8
rect 28 4 60 8
rect 64 4 82 8
rect 86 4 90 8
rect 94 4 114 8
rect -2 0 114 4
<< ntransistor >>
rect 12 12 14 26
rect 19 12 21 26
rect 31 7 33 26
rect 38 7 40 26
rect 48 7 50 26
rect 55 7 57 26
<< ptransistor >>
rect 9 39 11 66
rect 19 39 21 66
rect 29 39 31 66
rect 39 39 41 66
rect 49 39 51 66
rect 59 39 61 66
rect 69 39 71 66
rect 79 39 81 66
rect 90 39 92 56
rect 100 39 102 56
<< polycontact >>
rect 10 30 14 34
rect 26 30 30 34
rect 42 30 46 34
rect 58 30 62 34
rect 82 30 86 34
rect 97 30 101 34
<< ndcontact >>
rect 6 21 10 25
rect 6 14 10 18
rect 24 4 28 8
rect 42 14 46 18
rect 60 4 64 8
<< pdcontact >>
rect 3 61 7 65
rect 3 54 7 58
rect 13 53 17 57
rect 13 46 17 50
rect 23 61 27 65
rect 23 54 27 58
rect 33 54 37 58
rect 33 46 37 50
rect 43 61 47 65
rect 43 54 47 58
rect 53 53 57 57
rect 53 46 57 50
rect 63 61 67 65
rect 63 54 67 58
rect 73 54 77 58
rect 73 46 77 50
rect 83 61 87 65
rect 83 54 87 58
rect 94 46 98 50
rect 104 51 108 55
rect 104 43 108 47
<< psubstratepcontact >>
rect 82 4 86 8
rect 90 4 94 8
<< nsubstratencontact >>
rect 96 64 100 68
rect 104 64 108 68
<< psubstratepdiff >>
rect 81 8 95 24
rect 81 4 82 8
rect 86 4 90 8
rect 94 4 95 8
rect 81 3 95 4
<< nsubstratendiff >>
rect 95 68 109 69
rect 95 64 96 68
rect 100 64 104 68
rect 108 64 109 68
rect 95 63 109 64
<< labels >>
rlabel metal1 12 16 12 16 6 z
rlabel polycontact 12 32 12 32 6 b
rlabel metal1 4 32 4 32 6 z
rlabel metal1 12 48 12 48 6 z
rlabel metal1 28 16 28 16 6 z
rlabel metal1 36 16 36 16 6 z
rlabel metal1 20 16 20 16 6 z
rlabel metal1 20 24 20 24 6 b
rlabel metal1 28 24 28 24 6 b
rlabel metal1 36 24 36 24 6 b
rlabel polycontact 28 32 28 32 6 a
rlabel metal1 36 40 36 40 6 a
rlabel metal1 28 36 28 36 6 a
rlabel metal1 20 48 20 48 6 z
rlabel metal1 36 52 36 52 6 z
rlabel metal1 28 48 28 48 6 z
rlabel metal1 56 4 56 4 6 vss
rlabel ndcontact 44 16 44 16 6 z
rlabel metal1 52 24 52 24 6 b
rlabel metal1 60 24 60 24 6 b
rlabel metal1 44 28 44 28 6 b
rlabel metal1 44 40 44 40 6 a
rlabel metal1 52 40 52 40 6 a
rlabel metal1 60 36 60 36 6 a
rlabel metal1 44 48 44 48 6 z
rlabel metal1 52 48 52 48 6 z
rlabel metal1 60 48 60 48 6 z
rlabel metal1 56 68 56 68 6 vdd
rlabel metal1 68 24 68 24 6 b
rlabel metal1 76 24 76 24 6 b
rlabel metal1 84 28 84 28 6 b
rlabel metal1 68 40 68 40 6 a
rlabel metal1 76 40 76 40 6 a
rlabel metal1 84 40 84 40 6 a
rlabel metal1 68 48 68 48 6 z
rlabel metal1 76 52 76 52 6 z
rlabel metal1 84 48 84 48 6 z
rlabel polycontact 100 32 100 32 6 a
rlabel metal1 92 40 92 40 6 a
rlabel metal1 92 48 92 48 6 z
<< end >>
