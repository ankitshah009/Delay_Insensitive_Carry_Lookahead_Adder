magic
tech scmos
timestamp 1185039085
<< checkpaint >>
rect -22 -24 112 124
<< ab >>
rect 0 0 90 100
<< pwell >>
rect -2 -4 92 49
<< nwell >>
rect -2 49 92 104
<< polysilicon >>
rect 23 95 25 98
rect 35 95 37 98
rect 47 95 49 98
rect 59 95 61 98
rect 11 85 13 88
rect 11 53 13 65
rect 71 85 73 88
rect 23 53 25 55
rect 11 52 25 53
rect 11 51 18 52
rect 17 48 18 51
rect 22 51 25 52
rect 35 53 37 55
rect 35 52 43 53
rect 35 51 38 52
rect 22 48 23 51
rect 17 47 23 48
rect 37 48 38 51
rect 42 48 43 52
rect 37 47 43 48
rect 3 42 9 43
rect 3 38 4 42
rect 8 41 9 42
rect 47 41 49 55
rect 59 43 61 55
rect 71 53 73 65
rect 67 52 73 53
rect 67 48 68 52
rect 72 48 73 52
rect 67 47 73 48
rect 8 39 49 41
rect 8 38 9 39
rect 3 37 9 38
rect 17 32 23 33
rect 17 29 18 32
rect 11 28 18 29
rect 22 29 23 32
rect 37 32 43 33
rect 37 29 38 32
rect 22 28 25 29
rect 11 27 25 28
rect 11 25 13 27
rect 23 25 25 27
rect 35 28 38 29
rect 42 28 43 32
rect 35 27 43 28
rect 35 25 37 27
rect 47 25 49 39
rect 57 42 63 43
rect 57 38 58 42
rect 62 41 63 42
rect 77 42 83 43
rect 77 41 78 42
rect 62 39 78 41
rect 62 38 63 39
rect 57 37 63 38
rect 77 38 78 39
rect 82 38 83 42
rect 77 37 83 38
rect 67 32 73 33
rect 67 29 68 32
rect 59 28 68 29
rect 72 28 73 32
rect 59 27 73 28
rect 59 25 61 27
rect 71 25 73 27
rect 11 12 13 15
rect 71 12 73 15
rect 23 2 25 5
rect 35 2 37 5
rect 47 2 49 5
rect 59 2 61 5
<< ndiffusion >>
rect 3 22 11 25
rect 3 18 4 22
rect 8 18 11 22
rect 3 15 11 18
rect 13 15 23 25
rect 15 12 23 15
rect 15 8 16 12
rect 20 8 23 12
rect 15 5 23 8
rect 25 5 35 25
rect 37 22 47 25
rect 37 18 40 22
rect 44 18 47 22
rect 37 5 47 18
rect 49 5 59 25
rect 61 15 71 25
rect 73 22 83 25
rect 73 18 78 22
rect 82 18 83 22
rect 73 15 83 18
rect 61 12 69 15
rect 61 8 64 12
rect 68 8 69 12
rect 61 5 69 8
<< pdiffusion >>
rect 15 92 23 95
rect 15 88 16 92
rect 20 88 23 92
rect 15 85 23 88
rect 3 82 11 85
rect 3 78 4 82
rect 8 78 11 82
rect 3 72 11 78
rect 3 68 4 72
rect 8 68 11 72
rect 3 65 11 68
rect 13 65 23 85
rect 15 55 23 65
rect 25 82 35 95
rect 25 78 28 82
rect 32 78 35 82
rect 25 55 35 78
rect 37 72 47 95
rect 37 68 40 72
rect 44 68 47 72
rect 37 55 47 68
rect 49 82 59 95
rect 49 78 52 82
rect 56 78 59 82
rect 49 72 59 78
rect 49 68 52 72
rect 56 68 59 72
rect 49 62 59 68
rect 49 58 52 62
rect 56 58 59 62
rect 49 55 59 58
rect 61 92 69 95
rect 61 88 64 92
rect 68 88 69 92
rect 61 85 69 88
rect 61 65 71 85
rect 73 82 83 85
rect 73 78 78 82
rect 82 78 83 82
rect 73 72 83 78
rect 73 68 78 72
rect 82 68 83 72
rect 73 65 83 68
rect 61 55 69 65
<< metal1 >>
rect -2 96 92 101
rect -2 92 76 96
rect 80 92 92 96
rect -2 88 16 92
rect 20 88 64 92
rect 68 88 92 92
rect -2 87 92 88
rect 3 82 9 83
rect 27 82 33 83
rect 51 82 57 83
rect 77 82 83 83
rect 3 78 4 82
rect 8 78 9 82
rect 3 77 9 78
rect 4 73 8 77
rect 3 72 9 73
rect 3 68 4 72
rect 8 68 9 72
rect 3 67 9 68
rect 4 43 8 67
rect 17 52 23 82
rect 27 78 28 82
rect 32 78 52 82
rect 56 78 57 82
rect 27 77 33 78
rect 51 77 57 78
rect 52 73 56 77
rect 17 48 18 52
rect 22 48 23 52
rect 3 42 9 43
rect 3 38 4 42
rect 8 38 9 42
rect 3 37 9 38
rect 4 23 8 37
rect 17 32 23 48
rect 17 28 18 32
rect 22 28 23 32
rect 3 22 9 23
rect 3 18 4 22
rect 8 18 9 22
rect 17 18 23 28
rect 27 72 45 73
rect 27 68 40 72
rect 44 68 45 72
rect 27 67 45 68
rect 51 72 57 73
rect 51 68 52 72
rect 56 68 57 72
rect 51 67 57 68
rect 27 23 33 67
rect 52 63 56 67
rect 51 62 57 63
rect 51 58 52 62
rect 56 58 57 62
rect 51 57 57 58
rect 37 52 43 53
rect 67 52 73 82
rect 77 78 78 82
rect 82 78 83 82
rect 77 77 83 78
rect 78 73 82 77
rect 77 72 83 73
rect 77 68 78 72
rect 82 68 83 72
rect 77 67 83 68
rect 37 48 38 52
rect 42 48 68 52
rect 72 48 73 52
rect 37 47 43 48
rect 57 42 63 43
rect 48 38 58 42
rect 62 38 63 42
rect 37 32 43 33
rect 48 32 52 38
rect 57 37 63 38
rect 37 28 38 32
rect 42 28 52 32
rect 67 32 73 48
rect 78 43 82 67
rect 77 42 83 43
rect 77 38 78 42
rect 82 38 83 42
rect 77 37 83 38
rect 67 28 68 32
rect 72 28 73 32
rect 37 27 43 28
rect 27 22 45 23
rect 27 18 40 22
rect 44 18 45 22
rect 67 18 73 28
rect 78 23 82 37
rect 77 22 83 23
rect 77 18 78 22
rect 82 18 83 22
rect 3 17 9 18
rect 27 17 45 18
rect 77 17 83 18
rect -2 12 92 13
rect -2 8 16 12
rect 20 8 64 12
rect 68 8 92 12
rect -2 4 76 8
rect 80 4 92 8
rect -2 -1 92 4
<< ntransistor >>
rect 11 15 13 25
rect 23 5 25 25
rect 35 5 37 25
rect 47 5 49 25
rect 59 5 61 25
rect 71 15 73 25
<< ptransistor >>
rect 11 65 13 85
rect 23 55 25 95
rect 35 55 37 95
rect 47 55 49 95
rect 59 55 61 95
rect 71 65 73 85
<< polycontact >>
rect 18 48 22 52
rect 38 48 42 52
rect 4 38 8 42
rect 68 48 72 52
rect 18 28 22 32
rect 38 28 42 32
rect 58 38 62 42
rect 78 38 82 42
rect 68 28 72 32
<< ndcontact >>
rect 4 18 8 22
rect 16 8 20 12
rect 40 18 44 22
rect 78 18 82 22
rect 64 8 68 12
<< pdcontact >>
rect 16 88 20 92
rect 4 78 8 82
rect 4 68 8 72
rect 28 78 32 82
rect 40 68 44 72
rect 52 78 56 82
rect 52 68 56 72
rect 52 58 56 62
rect 64 88 68 92
rect 78 78 82 82
rect 78 68 82 72
<< psubstratepcontact >>
rect 76 4 80 8
<< nsubstratencontact >>
rect 76 92 80 96
<< psubstratepdiff >>
rect 75 8 87 9
rect 75 4 76 8
rect 80 4 87 8
rect 75 3 87 4
<< nsubstratendiff >>
rect 75 96 87 97
rect 75 92 76 96
rect 80 92 87 96
rect 75 91 87 92
<< labels >>
rlabel metal1 30 45 30 45 6 nq
rlabel metal1 30 45 30 45 6 nq
rlabel polycontact 20 50 20 50 6 i0
rlabel polycontact 20 50 20 50 6 i0
rlabel metal1 45 6 45 6 6 vss
rlabel metal1 45 6 45 6 6 vss
rlabel metal1 45 94 45 94 6 vdd
rlabel metal1 45 94 45 94 6 vdd
rlabel polycontact 70 50 70 50 6 i1
rlabel polycontact 70 50 70 50 6 i1
<< end >>
