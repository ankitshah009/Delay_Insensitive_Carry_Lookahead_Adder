magic
tech scmos
timestamp 1179387714
<< checkpaint >>
rect -22 -25 126 105
<< ab >>
rect 0 0 104 80
<< pwell >>
rect -4 -7 108 36
<< nwell >>
rect -4 36 108 87
<< polysilicon >>
rect 63 70 65 74
rect 73 70 75 74
rect 83 70 85 74
rect 93 70 95 74
rect 9 65 21 67
rect 9 62 11 65
rect 19 62 21 65
rect 29 65 50 67
rect 29 62 31 65
rect 39 62 41 65
rect 48 63 50 65
rect 48 62 54 63
rect 48 58 49 62
rect 53 58 54 62
rect 48 57 54 58
rect 63 47 65 50
rect 73 47 75 50
rect 83 47 85 50
rect 93 47 95 50
rect 55 46 79 47
rect 55 45 74 46
rect 9 38 11 42
rect 19 39 21 42
rect 18 38 24 39
rect 29 38 31 42
rect 18 34 19 38
rect 23 34 24 38
rect 39 35 41 42
rect 11 30 13 34
rect 18 33 24 34
rect 18 30 20 33
rect 28 30 30 34
rect 35 33 41 35
rect 35 30 37 33
rect 55 30 57 45
rect 73 42 74 45
rect 78 42 79 46
rect 73 41 79 42
rect 83 46 95 47
rect 83 42 90 46
rect 94 42 95 46
rect 83 41 95 42
rect 63 38 69 39
rect 63 34 64 38
rect 68 34 69 38
rect 63 33 69 34
rect 65 30 67 33
rect 75 30 77 41
rect 85 30 87 41
rect 11 8 13 17
rect 18 14 20 17
rect 28 14 30 17
rect 18 12 30 14
rect 35 8 37 17
rect 55 15 57 20
rect 85 15 87 20
rect 11 6 37 8
rect 65 6 67 10
rect 75 6 77 10
<< ndiffusion >>
rect 3 22 11 30
rect 3 18 5 22
rect 9 18 11 22
rect 3 17 11 18
rect 13 17 18 30
rect 20 29 28 30
rect 20 25 22 29
rect 26 25 28 29
rect 20 22 28 25
rect 20 18 22 22
rect 26 18 28 22
rect 20 17 28 18
rect 30 17 35 30
rect 37 22 55 30
rect 37 18 39 22
rect 43 20 55 22
rect 57 29 65 30
rect 57 25 59 29
rect 63 25 65 29
rect 57 20 65 25
rect 43 18 53 20
rect 37 17 53 18
rect 60 10 65 20
rect 67 29 75 30
rect 67 25 69 29
rect 73 25 75 29
rect 67 22 75 25
rect 67 18 69 22
rect 73 18 75 22
rect 67 10 75 18
rect 77 29 85 30
rect 77 25 79 29
rect 83 25 85 29
rect 77 20 85 25
rect 87 20 96 30
rect 77 10 82 20
rect 89 16 90 20
rect 94 16 96 20
rect 89 15 96 16
<< pdiffusion >>
rect 56 69 63 70
rect 56 65 57 69
rect 61 65 63 69
rect 4 55 9 62
rect 2 54 9 55
rect 2 50 3 54
rect 7 50 9 54
rect 2 47 9 50
rect 2 43 3 47
rect 7 43 9 47
rect 2 42 9 43
rect 11 61 19 62
rect 11 57 13 61
rect 17 57 19 61
rect 11 54 19 57
rect 11 50 13 54
rect 17 50 19 54
rect 11 42 19 50
rect 21 54 29 62
rect 21 50 23 54
rect 27 50 29 54
rect 21 47 29 50
rect 21 43 23 47
rect 27 43 29 47
rect 21 42 29 43
rect 31 47 39 62
rect 31 43 33 47
rect 37 43 39 47
rect 31 42 39 43
rect 41 55 46 62
rect 41 54 48 55
rect 41 50 43 54
rect 47 50 48 54
rect 56 50 63 65
rect 65 55 73 70
rect 65 51 67 55
rect 71 51 73 55
rect 65 50 73 51
rect 75 69 83 70
rect 75 65 77 69
rect 81 65 83 69
rect 75 50 83 65
rect 85 62 93 70
rect 85 58 87 62
rect 91 58 93 62
rect 85 50 93 58
rect 95 69 102 70
rect 95 65 97 69
rect 101 65 102 69
rect 95 50 102 65
rect 41 49 48 50
rect 41 42 46 49
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect -2 69 106 78
rect -2 68 57 69
rect 56 65 57 68
rect 61 68 77 69
rect 61 65 62 68
rect 76 65 77 68
rect 81 68 97 69
rect 81 65 82 68
rect 96 65 97 68
rect 101 68 106 69
rect 101 65 102 68
rect 12 61 49 62
rect 12 57 13 61
rect 17 58 49 61
rect 53 58 87 62
rect 91 58 102 62
rect 17 57 18 58
rect 2 54 7 55
rect 2 50 3 54
rect 12 54 18 57
rect 66 54 67 55
rect 12 50 13 54
rect 17 50 18 54
rect 22 50 23 54
rect 27 50 43 54
rect 47 50 48 54
rect 54 51 67 54
rect 71 51 72 55
rect 54 50 72 51
rect 2 47 7 50
rect 2 43 3 47
rect 22 47 27 50
rect 22 46 23 47
rect 7 43 23 46
rect 2 42 27 43
rect 32 43 33 47
rect 37 43 38 47
rect 32 42 38 43
rect 54 42 58 50
rect 82 46 86 55
rect 73 42 74 46
rect 78 42 86 46
rect 90 46 94 47
rect 2 30 6 42
rect 32 38 58 42
rect 90 38 94 42
rect 18 34 19 38
rect 23 34 38 38
rect 2 29 50 30
rect 2 26 22 29
rect 26 26 50 29
rect 22 22 26 25
rect 4 18 5 22
rect 9 18 10 22
rect 4 12 10 18
rect 22 17 26 18
rect 39 22 43 23
rect 46 22 50 26
rect 54 29 58 38
rect 63 34 64 38
rect 68 34 94 38
rect 69 29 74 30
rect 98 29 102 58
rect 54 25 59 29
rect 63 25 64 29
rect 73 25 74 29
rect 78 25 79 29
rect 83 25 102 29
rect 69 22 74 25
rect 46 18 69 22
rect 73 18 74 22
rect 90 20 94 21
rect 39 12 43 18
rect 90 12 94 16
rect -2 2 106 12
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
<< ntransistor >>
rect 11 17 13 30
rect 18 17 20 30
rect 28 17 30 30
rect 35 17 37 30
rect 55 20 57 30
rect 65 10 67 30
rect 75 10 77 30
rect 85 20 87 30
<< ptransistor >>
rect 9 42 11 62
rect 19 42 21 62
rect 29 42 31 62
rect 39 42 41 62
rect 63 50 65 70
rect 73 50 75 70
rect 83 50 85 70
rect 93 50 95 70
<< polycontact >>
rect 49 58 53 62
rect 19 34 23 38
rect 74 42 78 46
rect 90 42 94 46
rect 64 34 68 38
<< ndcontact >>
rect 5 18 9 22
rect 22 25 26 29
rect 22 18 26 22
rect 39 18 43 22
rect 59 25 63 29
rect 69 25 73 29
rect 69 18 73 22
rect 79 25 83 29
rect 90 16 94 20
<< pdcontact >>
rect 57 65 61 69
rect 3 50 7 54
rect 3 43 7 47
rect 13 57 17 61
rect 13 50 17 54
rect 23 50 27 54
rect 23 43 27 47
rect 33 43 37 47
rect 43 50 47 54
rect 67 51 71 55
rect 77 65 81 69
rect 87 58 91 62
rect 97 65 101 69
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
rect 90 -2 94 2
rect 98 -2 102 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
rect 90 78 94 82
rect 98 78 102 82
<< psubstratepdiff >>
rect 0 2 104 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 104 2
rect 0 -3 104 -2
<< nsubstratendiff >>
rect 0 82 104 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 104 82
rect 0 77 104 78
<< labels >>
rlabel ptransistor 20 50 20 50 6 bn
rlabel polycontact 51 60 51 60 6 an
rlabel metal1 12 28 12 28 6 z
rlabel pdcontact 4 44 4 44 6 z
rlabel metal1 12 44 12 44 6 z
rlabel metal1 15 56 15 56 6 an
rlabel metal1 20 28 20 28 6 z
rlabel metal1 28 28 28 28 6 z
rlabel metal1 36 28 36 28 6 z
rlabel metal1 20 44 20 44 6 z
rlabel metal1 28 36 28 36 6 bn
rlabel metal1 28 52 28 52 6 z
rlabel metal1 36 52 36 52 6 z
rlabel metal1 52 6 52 6 6 vss
rlabel metal1 44 28 44 28 6 z
rlabel metal1 60 20 60 20 6 z
rlabel metal1 52 20 52 20 6 z
rlabel metal1 45 40 45 40 6 bn
rlabel pdcontact 44 52 44 52 6 z
rlabel metal1 52 74 52 74 6 vdd
rlabel metal1 59 27 59 27 6 bn
rlabel metal1 68 20 68 20 6 z
rlabel metal1 76 36 76 36 6 a
rlabel metal1 68 36 68 36 6 a
rlabel polycontact 76 44 76 44 6 b
rlabel metal1 63 52 63 52 6 bn
rlabel metal1 90 27 90 27 6 an
rlabel metal1 84 36 84 36 6 a
rlabel polycontact 92 44 92 44 6 a
rlabel metal1 84 52 84 52 6 b
rlabel metal1 57 60 57 60 6 an
<< end >>
