magic
tech scmos
timestamp 1179386809
<< checkpaint >>
rect -22 -25 78 105
<< ab >>
rect 0 0 56 80
<< pwell >>
rect -4 -7 60 36
<< nwell >>
rect -4 36 60 87
<< polysilicon >>
rect 12 69 14 74
rect 19 69 21 74
rect 29 69 31 74
rect 36 69 38 74
rect 12 39 14 42
rect 19 39 21 42
rect 29 39 31 42
rect 36 39 38 42
rect 9 38 15 39
rect 9 34 10 38
rect 14 34 15 38
rect 9 33 15 34
rect 19 38 32 39
rect 19 34 27 38
rect 31 34 32 38
rect 19 33 32 34
rect 36 38 49 39
rect 36 34 44 38
rect 48 34 49 38
rect 36 33 49 34
rect 9 23 11 33
rect 19 23 21 33
rect 29 23 31 33
rect 39 30 41 33
rect 39 12 41 17
rect 9 6 11 10
rect 19 6 21 10
rect 29 6 31 10
<< ndiffusion >>
rect 34 23 39 30
rect 2 15 9 23
rect 2 11 3 15
rect 7 11 9 15
rect 2 10 9 11
rect 11 22 19 23
rect 11 18 13 22
rect 17 18 19 22
rect 11 10 19 18
rect 21 15 29 23
rect 21 11 23 15
rect 27 11 29 15
rect 21 10 29 11
rect 31 22 39 23
rect 31 18 33 22
rect 37 18 39 22
rect 31 17 39 18
rect 41 22 49 30
rect 41 18 43 22
rect 47 18 49 22
rect 41 17 49 18
rect 31 10 36 17
<< pdiffusion >>
rect 4 68 12 69
rect 4 64 6 68
rect 10 64 12 68
rect 4 60 12 64
rect 4 56 6 60
rect 10 56 12 60
rect 4 42 12 56
rect 14 42 19 69
rect 21 54 29 69
rect 21 50 23 54
rect 27 50 29 54
rect 21 47 29 50
rect 21 43 23 47
rect 27 43 29 47
rect 21 42 29 43
rect 31 42 36 69
rect 38 63 43 69
rect 38 62 46 63
rect 38 58 40 62
rect 44 58 46 62
rect 38 55 46 58
rect 38 51 40 55
rect 44 51 46 55
rect 38 42 46 51
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect -2 68 58 78
rect 6 60 10 64
rect 6 55 10 56
rect 40 62 44 68
rect 40 55 44 58
rect 22 50 23 54
rect 27 50 31 54
rect 40 50 44 51
rect 22 47 28 50
rect 2 43 23 47
rect 27 43 28 47
rect 2 22 6 43
rect 33 42 47 46
rect 10 38 22 39
rect 33 38 39 42
rect 14 34 22 38
rect 26 34 27 38
rect 31 34 39 38
rect 43 34 44 38
rect 48 34 49 38
rect 10 33 22 34
rect 17 30 22 33
rect 43 30 49 34
rect 17 26 49 30
rect 43 22 47 23
rect 2 18 13 22
rect 17 18 33 22
rect 37 18 39 22
rect 2 12 3 15
rect -2 11 3 12
rect 7 12 8 15
rect 22 12 23 15
rect 7 11 23 12
rect 27 12 28 15
rect 43 12 47 18
rect 27 11 58 12
rect -2 2 58 11
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
<< ntransistor >>
rect 9 10 11 23
rect 19 10 21 23
rect 29 10 31 23
rect 39 17 41 30
<< ptransistor >>
rect 12 42 14 69
rect 19 42 21 69
rect 29 42 31 69
rect 36 42 38 69
<< polycontact >>
rect 10 34 14 38
rect 27 34 31 38
rect 44 34 48 38
<< ndcontact >>
rect 3 11 7 15
rect 13 18 17 22
rect 23 11 27 15
rect 33 18 37 22
rect 43 18 47 22
<< pdcontact >>
rect 6 64 10 68
rect 6 56 10 60
rect 23 50 27 54
rect 23 43 27 47
rect 40 58 44 62
rect 40 51 44 55
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
<< psubstratepdiff >>
rect 0 2 56 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 56 2
rect 0 -3 56 -2
<< nsubstratendiff >>
rect 0 82 56 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 56 82
rect 0 77 56 78
<< labels >>
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 20 12 20 6 z
rlabel metal1 28 6 28 6 6 vss
rlabel metal1 20 20 20 20 6 z
rlabel metal1 28 28 28 28 6 a
rlabel metal1 28 20 28 20 6 z
rlabel metal1 20 32 20 32 6 a
rlabel metal1 28 52 28 52 6 z
rlabel metal1 28 74 28 74 6 vdd
rlabel ndcontact 36 20 36 20 6 z
rlabel metal1 36 28 36 28 6 a
rlabel metal1 44 28 44 28 6 a
rlabel metal1 36 40 36 40 6 b
rlabel metal1 44 44 44 44 6 b
<< end >>
