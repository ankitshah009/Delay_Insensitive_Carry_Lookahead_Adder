magic
tech scmos
timestamp 1179387172
<< checkpaint >>
rect -22 -22 86 94
<< ab >>
rect 0 0 64 72
<< pwell >>
rect -4 -4 68 32
<< nwell >>
rect -4 32 68 76
<< polysilicon >>
rect 9 59 11 64
rect 19 59 21 64
rect 29 59 31 64
rect 36 59 38 64
rect 46 55 48 60
rect 53 55 55 60
rect 9 35 11 39
rect 19 35 21 39
rect 9 34 21 35
rect 9 30 16 34
rect 20 30 21 34
rect 29 30 31 39
rect 36 36 38 39
rect 46 36 48 39
rect 36 34 48 36
rect 53 36 55 39
rect 53 35 62 36
rect 53 34 57 35
rect 38 33 48 34
rect 9 29 21 30
rect 28 29 34 30
rect 9 26 11 29
rect 28 25 29 29
rect 33 25 34 29
rect 28 24 34 25
rect 38 29 41 33
rect 45 29 48 33
rect 56 31 57 34
rect 61 31 62 35
rect 56 30 62 31
rect 38 28 48 29
rect 28 21 30 24
rect 38 21 40 28
rect 28 6 30 11
rect 38 6 40 11
rect 9 2 11 6
<< ndiffusion >>
rect 2 25 9 26
rect 2 21 3 25
rect 7 21 9 25
rect 2 18 9 21
rect 2 14 3 18
rect 7 14 9 18
rect 2 13 9 14
rect 4 6 9 13
rect 11 21 26 26
rect 11 19 28 21
rect 11 15 13 19
rect 17 15 28 19
rect 11 11 28 15
rect 30 20 38 21
rect 30 16 32 20
rect 36 16 38 20
rect 30 11 38 16
rect 40 16 48 21
rect 40 12 42 16
rect 46 12 48 16
rect 40 11 48 12
rect 11 7 13 11
rect 17 7 21 11
rect 25 7 26 11
rect 11 6 26 7
<< pdiffusion >>
rect 2 58 9 59
rect 2 54 3 58
rect 7 54 9 58
rect 2 51 9 54
rect 2 47 3 51
rect 7 47 9 51
rect 2 39 9 47
rect 11 51 19 59
rect 11 47 13 51
rect 17 47 19 51
rect 11 44 19 47
rect 11 40 13 44
rect 17 40 19 44
rect 11 39 19 40
rect 21 58 29 59
rect 21 54 23 58
rect 27 54 29 58
rect 21 39 29 54
rect 31 39 36 59
rect 38 55 43 59
rect 38 50 46 55
rect 38 46 40 50
rect 44 46 46 50
rect 38 39 46 46
rect 48 39 53 55
rect 55 54 62 55
rect 55 50 57 54
rect 61 50 62 54
rect 55 39 62 50
<< metal1 >>
rect -2 68 66 72
rect -2 64 48 68
rect 52 64 56 68
rect 60 64 66 68
rect 2 58 8 64
rect 2 54 3 58
rect 7 54 8 58
rect 22 58 28 64
rect 22 54 23 58
rect 27 54 28 58
rect 57 54 61 64
rect 2 51 8 54
rect 2 47 3 51
rect 7 47 8 51
rect 13 51 17 52
rect 13 44 17 47
rect 2 40 13 43
rect 2 38 17 40
rect 21 46 40 50
rect 44 46 45 50
rect 57 49 61 50
rect 2 26 6 38
rect 21 34 25 46
rect 58 42 62 43
rect 15 30 16 34
rect 20 30 25 34
rect 2 25 7 26
rect 2 21 3 25
rect 2 18 7 21
rect 21 20 25 30
rect 29 38 62 42
rect 29 29 33 38
rect 56 35 62 38
rect 29 24 33 25
rect 41 33 47 34
rect 45 29 47 33
rect 56 31 57 35
rect 61 31 62 35
rect 58 29 62 31
rect 41 27 47 29
rect 41 21 54 27
rect 2 14 3 18
rect 2 13 7 14
rect 13 19 17 20
rect 21 16 32 20
rect 36 16 37 20
rect 42 16 46 17
rect 13 11 17 15
rect -2 7 13 8
rect 21 11 25 12
rect 17 7 21 8
rect 42 8 46 12
rect 25 7 56 8
rect -2 4 56 7
rect 60 4 66 8
rect -2 0 66 4
<< ntransistor >>
rect 9 6 11 26
rect 28 11 30 21
rect 38 11 40 21
<< ptransistor >>
rect 9 39 11 59
rect 19 39 21 59
rect 29 39 31 59
rect 36 39 38 59
rect 46 39 48 55
rect 53 39 55 55
<< polycontact >>
rect 16 30 20 34
rect 29 25 33 29
rect 41 29 45 33
rect 57 31 61 35
<< ndcontact >>
rect 3 21 7 25
rect 3 14 7 18
rect 13 15 17 19
rect 32 16 36 20
rect 42 12 46 16
rect 13 7 17 11
rect 21 7 25 11
<< pdcontact >>
rect 3 54 7 58
rect 3 47 7 51
rect 13 47 17 51
rect 13 40 17 44
rect 23 54 27 58
rect 40 46 44 50
rect 57 50 61 54
<< psubstratepcontact >>
rect 56 4 60 8
<< nsubstratencontact >>
rect 48 64 52 68
rect 56 64 60 68
<< psubstratepdiff >>
rect 55 8 61 26
rect 55 4 56 8
rect 60 4 61 8
rect 55 3 61 4
<< nsubstratendiff >>
rect 47 68 61 69
rect 47 64 48 68
rect 52 64 56 68
rect 60 64 61 68
rect 47 63 61 64
<< labels >>
rlabel polysilicon 15 32 15 32 6 zn
rlabel metal1 4 28 4 28 6 z
rlabel metal1 12 40 12 40 6 z
rlabel metal1 20 32 20 32 6 zn
rlabel metal1 32 4 32 4 6 vss
rlabel metal1 29 18 29 18 6 zn
rlabel metal1 44 28 44 28 6 b
rlabel metal1 44 40 44 40 6 a
rlabel metal1 36 40 36 40 6 a
rlabel metal1 33 48 33 48 6 zn
rlabel metal1 32 68 32 68 6 vdd
rlabel metal1 52 24 52 24 6 b
rlabel metal1 60 36 60 36 6 a
rlabel metal1 52 40 52 40 6 a
<< end >>
