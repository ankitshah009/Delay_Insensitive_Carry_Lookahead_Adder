magic
tech scmos
timestamp 1179387248
<< checkpaint >>
rect -22 -25 126 105
<< ab >>
rect 0 0 104 80
<< pwell >>
rect -4 -7 108 36
<< nwell >>
rect -4 36 108 87
<< polysilicon >>
rect 9 70 11 74
rect 19 70 21 74
rect 31 70 33 74
rect 38 70 40 74
rect 45 70 47 74
rect 55 70 57 74
rect 62 70 64 74
rect 69 70 71 74
rect 79 58 81 63
rect 86 58 88 63
rect 93 58 95 63
rect 9 39 11 42
rect 19 39 21 42
rect 31 39 33 42
rect 9 38 21 39
rect 9 34 16 38
rect 20 34 21 38
rect 9 33 21 34
rect 28 38 34 39
rect 28 34 29 38
rect 33 34 34 38
rect 28 33 34 34
rect 38 33 40 42
rect 45 39 47 42
rect 55 39 57 42
rect 45 37 57 39
rect 9 30 11 33
rect 19 30 21 33
rect 29 24 31 33
rect 38 32 47 33
rect 38 28 42 32
rect 46 28 47 32
rect 38 27 47 28
rect 39 24 41 27
rect 51 24 53 37
rect 62 31 64 42
rect 69 39 71 42
rect 79 39 81 42
rect 69 38 81 39
rect 69 37 74 38
rect 73 34 74 37
rect 78 37 81 38
rect 78 34 79 37
rect 73 33 79 34
rect 62 30 68 31
rect 62 26 63 30
rect 67 29 68 30
rect 86 29 88 42
rect 67 27 88 29
rect 93 39 95 42
rect 93 38 99 39
rect 93 34 94 38
rect 98 34 99 38
rect 93 33 99 34
rect 67 26 68 27
rect 62 25 68 26
rect 9 11 11 16
rect 19 11 21 16
rect 29 6 31 11
rect 39 6 41 11
rect 93 23 95 33
rect 86 21 95 23
rect 51 8 53 11
rect 86 8 88 21
rect 51 6 88 8
<< ndiffusion >>
rect 2 21 9 30
rect 2 17 3 21
rect 7 17 9 21
rect 2 16 9 17
rect 11 29 19 30
rect 11 25 13 29
rect 17 25 19 29
rect 11 22 19 25
rect 11 18 13 22
rect 17 18 19 22
rect 11 16 19 18
rect 21 24 27 30
rect 21 21 29 24
rect 21 17 23 21
rect 27 17 29 21
rect 21 16 29 17
rect 23 11 29 16
rect 31 21 39 24
rect 31 17 33 21
rect 37 17 39 21
rect 31 11 39 17
rect 41 12 51 24
rect 41 11 44 12
rect 43 8 44 11
rect 48 11 51 12
rect 53 22 58 24
rect 53 21 60 22
rect 53 17 55 21
rect 59 17 60 21
rect 53 16 60 17
rect 53 11 58 16
rect 48 8 49 11
rect 43 7 49 8
<< pdiffusion >>
rect 2 69 9 70
rect 2 65 3 69
rect 7 65 9 69
rect 2 62 9 65
rect 2 58 3 62
rect 7 58 9 62
rect 2 42 9 58
rect 11 54 19 70
rect 11 50 13 54
rect 17 50 19 54
rect 11 47 19 50
rect 11 43 13 47
rect 17 43 19 47
rect 11 42 19 43
rect 21 69 31 70
rect 21 65 24 69
rect 28 65 31 69
rect 21 62 31 65
rect 21 58 24 62
rect 28 58 31 62
rect 21 42 31 58
rect 33 42 38 70
rect 40 42 45 70
rect 47 61 55 70
rect 47 57 49 61
rect 53 57 55 61
rect 47 54 55 57
rect 47 50 49 54
rect 53 50 55 54
rect 47 42 55 50
rect 57 42 62 70
rect 64 42 69 70
rect 71 58 77 70
rect 71 57 79 58
rect 71 53 73 57
rect 77 53 79 57
rect 71 42 79 53
rect 81 42 86 58
rect 88 42 93 58
rect 95 55 100 58
rect 95 54 102 55
rect 95 50 97 54
rect 101 50 102 54
rect 95 47 102 50
rect 95 43 97 47
rect 101 43 102 47
rect 95 42 102 43
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect -2 69 106 78
rect -2 68 3 69
rect 2 65 3 68
rect 7 68 24 69
rect 7 65 8 68
rect 2 62 8 65
rect 2 58 3 62
rect 7 58 8 62
rect 23 65 24 68
rect 28 68 106 69
rect 28 65 29 68
rect 23 62 29 65
rect 23 58 24 62
rect 28 58 29 62
rect 49 61 53 62
rect 2 46 6 55
rect 13 54 17 55
rect 49 54 53 57
rect 73 57 77 68
rect 13 47 17 50
rect 2 43 13 46
rect 2 42 17 43
rect 21 50 49 54
rect 53 50 67 54
rect 73 52 77 53
rect 2 30 6 42
rect 21 38 25 50
rect 63 47 67 50
rect 96 50 97 54
rect 101 50 102 54
rect 96 47 102 50
rect 33 42 55 46
rect 63 43 97 47
rect 101 43 102 47
rect 33 39 38 42
rect 15 34 16 38
rect 20 34 25 38
rect 2 29 17 30
rect 2 25 13 29
rect 21 29 25 34
rect 29 38 38 39
rect 33 34 38 38
rect 51 38 55 42
rect 89 38 102 39
rect 51 34 74 38
rect 78 34 79 38
rect 89 34 94 38
rect 98 34 102 38
rect 29 33 38 34
rect 89 33 102 34
rect 42 32 46 33
rect 21 25 36 29
rect 46 28 63 30
rect 42 26 63 28
rect 67 26 71 30
rect 89 26 95 33
rect 13 22 17 25
rect 2 17 3 21
rect 7 17 8 21
rect 32 21 36 25
rect 13 17 17 18
rect 22 17 23 21
rect 27 17 28 21
rect 32 17 33 21
rect 37 17 55 21
rect 59 17 60 21
rect 65 18 71 26
rect 2 12 8 17
rect 22 12 28 17
rect -2 8 44 12
rect 48 8 106 12
rect -2 2 106 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
<< ntransistor >>
rect 9 16 11 30
rect 19 16 21 30
rect 29 11 31 24
rect 39 11 41 24
rect 51 11 53 24
<< ptransistor >>
rect 9 42 11 70
rect 19 42 21 70
rect 31 42 33 70
rect 38 42 40 70
rect 45 42 47 70
rect 55 42 57 70
rect 62 42 64 70
rect 69 42 71 70
rect 79 42 81 58
rect 86 42 88 58
rect 93 42 95 58
<< polycontact >>
rect 16 34 20 38
rect 29 34 33 38
rect 42 28 46 32
rect 74 34 78 38
rect 63 26 67 30
rect 94 34 98 38
<< ndcontact >>
rect 3 17 7 21
rect 13 25 17 29
rect 13 18 17 22
rect 23 17 27 21
rect 33 17 37 21
rect 44 8 48 12
rect 55 17 59 21
<< pdcontact >>
rect 3 65 7 69
rect 3 58 7 62
rect 13 50 17 54
rect 13 43 17 47
rect 24 65 28 69
rect 24 58 28 62
rect 49 57 53 61
rect 49 50 53 54
rect 73 53 77 57
rect 97 50 101 54
rect 97 43 101 47
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
rect 90 -2 94 2
rect 98 -2 102 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
rect 90 78 94 82
rect 98 78 102 82
<< psubstratepdiff >>
rect 0 2 104 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 104 2
rect 0 -3 104 -2
<< nsubstratendiff >>
rect 0 82 104 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 104 82
rect 0 77 104 78
<< labels >>
rlabel polysilicon 15 36 15 36 6 zn
rlabel metal1 12 28 12 28 6 z
rlabel metal1 4 40 4 40 6 z
rlabel metal1 12 44 12 44 6 z
rlabel metal1 20 36 20 36 6 zn
rlabel metal1 36 40 36 40 6 a
rlabel metal1 52 6 52 6 6 vss
rlabel metal1 46 19 46 19 6 zn
rlabel metal1 52 28 52 28 6 b
rlabel metal1 60 28 60 28 6 b
rlabel metal1 44 44 44 44 6 a
rlabel metal1 52 44 52 44 6 a
rlabel metal1 60 36 60 36 6 a
rlabel metal1 51 56 51 56 6 zn
rlabel metal1 52 74 52 74 6 vdd
rlabel metal1 68 24 68 24 6 b
rlabel metal1 68 36 68 36 6 a
rlabel polycontact 76 36 76 36 6 a
rlabel metal1 44 52 44 52 6 zn
rlabel metal1 92 32 92 32 6 c
rlabel metal1 82 45 82 45 6 zn
rlabel metal1 100 36 100 36 6 c
rlabel metal1 99 48 99 48 6 zn
<< end >>
