magic
tech scmos
timestamp 1179387575
<< checkpaint >>
rect -22 -22 118 94
<< ab >>
rect 0 0 96 72
<< pwell >>
rect -4 -4 100 32
<< nwell >>
rect -4 32 100 76
<< polysilicon >>
rect 12 66 14 70
rect 19 66 21 70
rect 31 66 33 70
rect 38 66 40 70
rect 48 66 50 70
rect 58 66 60 70
rect 68 66 70 70
rect 75 66 77 70
rect 85 66 87 70
rect 12 35 14 38
rect 9 34 15 35
rect 9 30 10 34
rect 14 30 15 34
rect 9 29 15 30
rect 9 26 11 29
rect 19 26 21 38
rect 31 35 33 46
rect 38 43 40 46
rect 48 43 50 46
rect 58 43 60 46
rect 68 43 70 46
rect 38 41 43 43
rect 48 42 61 43
rect 48 41 56 42
rect 41 37 43 41
rect 55 38 56 41
rect 60 38 61 42
rect 55 37 61 38
rect 65 41 70 43
rect 41 35 51 37
rect 31 34 37 35
rect 31 30 32 34
rect 36 31 37 34
rect 49 31 51 35
rect 65 31 67 41
rect 75 35 77 46
rect 85 35 87 38
rect 36 30 44 31
rect 31 29 44 30
rect 49 29 67 31
rect 71 34 77 35
rect 71 30 72 34
rect 76 30 77 34
rect 71 29 77 30
rect 81 34 87 35
rect 81 30 82 34
rect 86 30 87 34
rect 81 29 87 30
rect 42 26 44 29
rect 52 26 54 29
rect 61 26 67 29
rect 28 17 34 18
rect 28 13 29 17
rect 33 13 34 17
rect 28 12 34 13
rect 61 22 62 26
rect 66 22 67 26
rect 84 24 86 29
rect 61 21 67 22
rect 9 7 11 12
rect 19 9 21 12
rect 28 9 30 12
rect 19 7 30 9
rect 42 9 44 14
rect 52 9 54 14
rect 84 6 86 11
<< ndiffusion >>
rect 4 18 9 26
rect 2 17 9 18
rect 2 13 3 17
rect 7 13 9 17
rect 2 12 9 13
rect 11 25 19 26
rect 11 21 13 25
rect 17 21 19 25
rect 11 12 19 21
rect 21 25 28 26
rect 21 21 23 25
rect 27 21 28 25
rect 21 20 28 21
rect 21 12 26 20
rect 36 14 42 26
rect 44 25 52 26
rect 44 21 46 25
rect 50 21 52 25
rect 44 14 52 21
rect 54 18 59 26
rect 77 23 84 24
rect 77 19 78 23
rect 82 19 84 23
rect 77 18 84 19
rect 54 14 62 18
rect 36 10 40 14
rect 34 8 40 10
rect 34 4 35 8
rect 39 4 40 8
rect 34 3 40 4
rect 56 8 62 14
rect 56 4 57 8
rect 61 4 62 8
rect 56 3 62 4
rect 79 11 84 18
rect 86 16 94 24
rect 86 12 88 16
rect 92 12 94 16
rect 86 11 94 12
<< pdiffusion >>
rect 7 58 12 66
rect 5 57 12 58
rect 5 53 6 57
rect 10 53 12 57
rect 5 50 12 53
rect 5 46 6 50
rect 10 46 12 50
rect 5 45 12 46
rect 7 38 12 45
rect 14 38 19 66
rect 21 65 31 66
rect 21 61 24 65
rect 28 61 31 65
rect 21 46 31 61
rect 33 46 38 66
rect 40 51 48 66
rect 40 47 42 51
rect 46 47 48 51
rect 40 46 48 47
rect 50 58 58 66
rect 50 54 52 58
rect 56 54 58 58
rect 50 46 58 54
rect 60 58 68 66
rect 60 54 62 58
rect 66 54 68 58
rect 60 51 68 54
rect 60 47 62 51
rect 66 47 68 51
rect 60 46 68 47
rect 70 46 75 66
rect 77 65 85 66
rect 77 61 79 65
rect 83 61 85 65
rect 77 58 85 61
rect 77 54 79 58
rect 83 54 85 58
rect 77 46 85 54
rect 21 38 26 46
rect 80 38 85 46
rect 87 59 92 66
rect 87 58 94 59
rect 87 54 89 58
rect 93 54 94 58
rect 87 51 94 54
rect 87 47 89 51
rect 93 47 94 51
rect 87 46 94 47
rect 87 38 92 46
<< metal1 >>
rect -2 65 98 72
rect -2 64 24 65
rect 23 61 24 64
rect 28 64 79 65
rect 28 61 29 64
rect 78 61 79 64
rect 83 64 98 65
rect 83 61 84 64
rect 62 58 67 59
rect 6 57 10 58
rect 6 51 10 53
rect 2 50 10 51
rect 25 54 52 58
rect 56 54 57 58
rect 66 54 67 58
rect 78 58 84 61
rect 78 54 79 58
rect 83 54 84 58
rect 89 58 94 59
rect 93 54 94 58
rect 25 50 31 54
rect 62 51 67 54
rect 2 25 6 50
rect 10 46 31 50
rect 34 47 42 51
rect 46 47 62 51
rect 66 47 67 51
rect 89 51 94 54
rect 34 42 38 47
rect 22 38 38 42
rect 22 34 26 38
rect 42 34 46 43
rect 73 42 79 50
rect 93 47 94 51
rect 89 46 94 47
rect 55 38 56 42
rect 60 38 86 42
rect 82 34 86 38
rect 9 30 10 34
rect 14 30 26 34
rect 31 30 32 34
rect 36 30 72 34
rect 76 30 77 34
rect 22 25 26 30
rect 82 29 86 30
rect 2 21 13 25
rect 17 21 18 25
rect 22 21 23 25
rect 27 21 46 25
rect 50 21 51 25
rect 57 22 62 26
rect 66 22 71 26
rect 90 25 94 46
rect 78 23 94 25
rect 82 21 94 23
rect 78 17 82 19
rect 2 13 3 17
rect 7 13 29 17
rect 33 13 82 17
rect 88 16 92 17
rect 88 8 92 12
rect -2 4 35 8
rect 39 4 57 8
rect 61 4 68 8
rect 72 4 98 8
rect -2 0 98 4
<< ntransistor >>
rect 9 12 11 26
rect 19 12 21 26
rect 42 14 44 26
rect 52 14 54 26
rect 84 11 86 24
<< ptransistor >>
rect 12 38 14 66
rect 19 38 21 66
rect 31 46 33 66
rect 38 46 40 66
rect 48 46 50 66
rect 58 46 60 66
rect 68 46 70 66
rect 75 46 77 66
rect 85 38 87 66
<< polycontact >>
rect 10 30 14 34
rect 56 38 60 42
rect 32 30 36 34
rect 72 30 76 34
rect 82 30 86 34
rect 29 13 33 17
rect 62 22 66 26
<< ndcontact >>
rect 3 13 7 17
rect 13 21 17 25
rect 23 21 27 25
rect 46 21 50 25
rect 78 19 82 23
rect 35 4 39 8
rect 57 4 61 8
rect 88 12 92 16
<< pdcontact >>
rect 6 53 10 57
rect 6 46 10 50
rect 24 61 28 65
rect 42 47 46 51
rect 52 54 56 58
rect 62 54 66 58
rect 62 47 66 51
rect 79 61 83 65
rect 79 54 83 58
rect 89 54 93 58
rect 89 47 93 51
<< psubstratepcontact >>
rect 68 4 72 8
<< psubstratepdiff >>
rect 67 8 73 18
rect 67 4 68 8
rect 72 4 73 8
rect 67 3 73 4
<< labels >>
rlabel ptransistor 13 49 13 49 6 an
rlabel polycontact 31 15 31 15 6 bn
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 48 12 48 6 z
rlabel metal1 17 32 17 32 6 an
rlabel metal1 20 48 20 48 6 z
rlabel metal1 28 52 28 52 6 z
rlabel metal1 48 4 48 4 6 vss
rlabel metal1 36 23 36 23 6 an
rlabel metal1 52 32 52 32 6 a1
rlabel metal1 36 32 36 32 6 a1
rlabel metal1 44 36 44 36 6 a1
rlabel metal1 44 56 44 56 6 z
rlabel metal1 52 56 52 56 6 z
rlabel metal1 36 56 36 56 6 z
rlabel metal1 48 68 48 68 6 vdd
rlabel metal1 60 24 60 24 6 a2
rlabel metal1 68 24 68 24 6 a2
rlabel metal1 68 32 68 32 6 a1
rlabel metal1 60 32 60 32 6 a1
rlabel metal1 60 40 60 40 6 b
rlabel metal1 68 40 68 40 6 b
rlabel metal1 76 44 76 44 6 b
rlabel metal1 50 49 50 49 6 an
rlabel metal1 64 53 64 53 6 an
rlabel metal1 80 19 80 19 6 bn
rlabel metal1 42 15 42 15 6 bn
rlabel polycontact 84 32 84 32 6 b
rlabel metal1 92 40 92 40 6 bn
<< end >>
