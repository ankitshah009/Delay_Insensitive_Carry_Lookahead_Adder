magic
tech scmos
timestamp 1179387495
<< checkpaint >>
rect -22 -25 86 105
<< ab >>
rect 0 0 64 80
<< pwell >>
rect -4 -7 68 36
<< nwell >>
rect -4 36 68 87
<< polysilicon >>
rect 11 71 34 73
rect 11 65 13 71
rect 9 63 13 65
rect 22 63 24 67
rect 32 63 34 71
rect 42 70 44 74
rect 49 70 51 74
rect 9 60 11 63
rect 9 39 11 42
rect 22 39 24 45
rect 32 40 34 45
rect 42 39 44 42
rect 49 39 51 42
rect 9 38 18 39
rect 9 37 13 38
rect 12 34 13 37
rect 17 34 18 38
rect 12 33 18 34
rect 22 38 28 39
rect 22 34 23 38
rect 27 34 28 38
rect 22 33 28 34
rect 38 37 44 39
rect 48 38 54 39
rect 2 30 8 31
rect 2 26 3 30
rect 7 26 8 30
rect 15 26 17 33
rect 25 26 27 33
rect 38 31 40 37
rect 48 34 49 38
rect 53 34 54 38
rect 48 33 54 34
rect 48 31 50 33
rect 35 29 40 31
rect 45 29 50 31
rect 35 26 37 29
rect 45 26 47 29
rect 2 25 8 26
rect 4 9 6 25
rect 56 22 62 23
rect 56 18 57 22
rect 61 18 62 22
rect 56 17 62 18
rect 15 13 17 17
rect 25 13 27 17
rect 35 9 37 17
rect 45 13 47 17
rect 56 9 58 17
rect 4 7 58 9
<< ndiffusion >>
rect 10 23 15 26
rect 8 22 15 23
rect 8 18 9 22
rect 13 18 15 22
rect 8 17 15 18
rect 17 22 25 26
rect 17 18 19 22
rect 23 18 25 22
rect 17 17 25 18
rect 27 25 35 26
rect 27 21 29 25
rect 33 21 35 25
rect 27 17 35 21
rect 37 22 45 26
rect 37 18 39 22
rect 43 18 45 22
rect 37 17 45 18
rect 47 23 52 26
rect 47 22 54 23
rect 47 18 49 22
rect 53 18 54 22
rect 47 17 54 18
<< pdiffusion >>
rect 37 63 42 70
rect 15 62 22 63
rect 15 60 16 62
rect 4 55 9 60
rect 2 54 9 55
rect 2 50 3 54
rect 7 50 9 54
rect 2 47 9 50
rect 2 43 3 47
rect 7 43 9 47
rect 2 42 9 43
rect 11 58 16 60
rect 20 58 22 62
rect 11 45 22 58
rect 24 57 32 63
rect 24 53 26 57
rect 30 53 32 57
rect 24 50 32 53
rect 24 46 26 50
rect 30 46 32 50
rect 24 45 32 46
rect 34 54 42 63
rect 34 50 36 54
rect 40 50 42 54
rect 34 45 42 50
rect 11 42 16 45
rect 37 42 42 45
rect 44 42 49 70
rect 51 69 59 70
rect 51 65 53 69
rect 57 65 59 69
rect 51 62 59 65
rect 51 58 53 62
rect 57 58 59 62
rect 51 42 59 58
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect -2 69 66 78
rect -2 68 53 69
rect 15 62 21 68
rect 15 58 16 62
rect 20 58 21 62
rect 52 65 53 68
rect 57 68 66 69
rect 57 65 58 68
rect 52 62 58 65
rect 52 58 53 62
rect 57 58 58 62
rect 26 57 30 58
rect 2 54 7 55
rect 2 50 3 54
rect 2 47 7 50
rect 18 47 22 55
rect 2 43 3 47
rect 2 42 7 43
rect 10 43 22 47
rect 26 50 30 53
rect 35 50 36 54
rect 40 50 62 54
rect 2 31 6 42
rect 10 41 17 43
rect 26 42 38 46
rect 13 38 17 41
rect 34 38 38 42
rect 13 33 17 34
rect 21 34 23 38
rect 27 34 31 38
rect 34 34 49 38
rect 53 34 54 38
rect 2 30 7 31
rect 21 30 25 34
rect 2 26 3 30
rect 17 26 25 30
rect 34 29 38 34
rect 58 30 62 50
rect 2 22 7 26
rect 29 25 38 29
rect 41 26 62 30
rect 2 18 9 22
rect 13 18 14 22
rect 18 18 19 22
rect 23 18 24 22
rect 41 22 45 26
rect 29 20 33 21
rect 38 18 39 22
rect 43 18 45 22
rect 48 18 49 22
rect 53 18 57 22
rect 61 18 62 22
rect 18 12 24 18
rect -2 2 66 12
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
<< ntransistor >>
rect 15 17 17 26
rect 25 17 27 26
rect 35 17 37 26
rect 45 17 47 26
<< ptransistor >>
rect 9 42 11 60
rect 22 45 24 63
rect 32 45 34 63
rect 42 42 44 70
rect 49 42 51 70
<< polycontact >>
rect 13 34 17 38
rect 23 34 27 38
rect 3 26 7 30
rect 49 34 53 38
rect 57 18 61 22
<< ndcontact >>
rect 9 18 13 22
rect 19 18 23 22
rect 29 21 33 25
rect 39 18 43 22
rect 49 18 53 22
<< pdcontact >>
rect 3 50 7 54
rect 3 43 7 47
rect 16 58 20 62
rect 26 53 30 57
rect 26 46 30 50
rect 36 50 40 54
rect 53 65 57 69
rect 53 58 57 62
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
<< psubstratepdiff >>
rect 0 2 64 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 64 2
rect 0 -3 64 -2
<< nsubstratendiff >>
rect 0 82 64 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 64 82
rect 0 77 64 78
<< labels >>
rlabel polysilicon 5 19 5 19 6 bn
rlabel polycontact 59 20 59 20 6 bn
rlabel ptransistor 50 53 50 53 6 an
rlabel metal1 4 36 4 36 6 bn
rlabel metal1 8 20 8 20 6 bn
rlabel metal1 20 28 20 28 6 a
rlabel metal1 12 44 12 44 6 b
rlabel metal1 20 52 20 52 6 b
rlabel metal1 32 6 32 6 6 vss
rlabel ndcontact 31 24 31 24 6 an
rlabel metal1 28 36 28 36 6 a
rlabel metal1 28 50 28 50 6 an
rlabel metal1 32 74 32 74 6 vdd
rlabel metal1 44 28 44 28 6 z
rlabel metal1 44 52 44 52 6 z
rlabel metal1 52 28 52 28 6 z
rlabel metal1 55 20 55 20 6 bn
rlabel metal1 44 36 44 36 6 an
rlabel metal1 60 40 60 40 6 z
rlabel metal1 52 52 52 52 6 z
<< end >>
