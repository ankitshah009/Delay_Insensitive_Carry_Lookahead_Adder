magic
tech scmos
timestamp 1179387630
<< checkpaint >>
rect -22 -25 86 105
<< ab >>
rect 0 0 64 80
<< pwell >>
rect -4 -7 68 36
<< nwell >>
rect -4 36 68 87
<< polysilicon >>
rect 10 66 21 68
rect 10 64 12 66
rect 6 63 12 64
rect 19 63 21 66
rect 39 63 45 64
rect 53 63 55 68
rect 6 59 7 63
rect 11 59 12 63
rect 6 58 12 59
rect 33 55 35 60
rect 39 59 40 63
rect 44 59 45 63
rect 39 58 45 59
rect 43 55 45 58
rect 19 39 21 42
rect 33 39 35 42
rect 13 37 21 39
rect 25 38 35 39
rect 13 30 15 37
rect 25 34 26 38
rect 30 37 35 38
rect 30 34 31 37
rect 25 33 31 34
rect 26 24 28 33
rect 43 29 45 42
rect 53 39 55 42
rect 49 38 55 39
rect 49 34 50 38
rect 54 34 55 38
rect 49 33 55 34
rect 36 24 38 29
rect 43 27 48 29
rect 46 24 48 27
rect 53 24 55 33
rect 13 9 15 23
rect 26 13 28 17
rect 36 9 38 17
rect 46 10 48 15
rect 53 10 55 15
rect 13 7 38 9
<< ndiffusion >>
rect 6 29 13 30
rect 6 25 7 29
rect 11 25 13 29
rect 6 23 13 25
rect 15 24 24 30
rect 15 23 26 24
rect 17 22 26 23
rect 17 18 18 22
rect 22 18 26 22
rect 17 17 26 18
rect 28 22 36 24
rect 28 18 30 22
rect 34 18 36 22
rect 28 17 36 18
rect 38 22 46 24
rect 38 18 40 22
rect 44 18 46 22
rect 38 17 46 18
rect 41 15 46 17
rect 48 15 53 24
rect 55 20 62 24
rect 55 16 57 20
rect 61 16 62 20
rect 55 15 62 16
<< pdiffusion >>
rect 14 48 19 63
rect 12 47 19 48
rect 12 43 13 47
rect 17 43 19 47
rect 12 42 19 43
rect 21 62 31 63
rect 21 58 23 62
rect 27 58 31 62
rect 21 55 31 58
rect 48 55 53 63
rect 21 42 33 55
rect 35 47 43 55
rect 35 43 37 47
rect 41 43 43 47
rect 35 42 43 43
rect 45 54 53 55
rect 45 50 47 54
rect 51 50 53 54
rect 45 47 53 50
rect 45 43 47 47
rect 51 43 53 47
rect 45 42 53 43
rect 55 62 62 63
rect 55 58 57 62
rect 61 58 62 62
rect 55 55 62 58
rect 55 51 57 55
rect 61 51 62 55
rect 55 50 62 51
rect 55 42 60 50
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect -2 68 66 78
rect 2 59 7 63
rect 11 59 15 63
rect 2 58 15 59
rect 22 62 28 68
rect 22 58 23 62
rect 27 58 28 62
rect 32 59 40 63
rect 44 62 61 63
rect 44 59 57 62
rect 2 49 6 58
rect 32 54 36 59
rect 57 55 61 58
rect 13 50 36 54
rect 47 54 51 55
rect 57 50 61 51
rect 13 47 17 50
rect 47 47 51 50
rect 7 43 13 46
rect 7 42 17 43
rect 36 43 37 47
rect 41 43 42 47
rect 7 29 11 42
rect 36 38 42 43
rect 51 43 62 46
rect 47 42 62 43
rect 17 34 26 38
rect 30 34 31 38
rect 36 34 50 38
rect 54 34 55 38
rect 17 26 23 34
rect 36 30 40 34
rect 58 30 62 42
rect 30 26 40 30
rect 49 26 62 30
rect 7 24 11 25
rect 30 22 34 26
rect 49 22 53 26
rect 17 18 18 22
rect 22 18 23 22
rect 17 12 23 18
rect 39 18 40 22
rect 44 18 53 22
rect 57 20 61 21
rect 30 17 34 18
rect 57 12 61 16
rect -2 2 66 12
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
<< ntransistor >>
rect 13 23 15 30
rect 26 17 28 24
rect 36 17 38 24
rect 46 15 48 24
rect 53 15 55 24
<< ptransistor >>
rect 19 42 21 63
rect 33 42 35 55
rect 43 42 45 55
rect 53 42 55 63
<< polycontact >>
rect 7 59 11 63
rect 40 59 44 63
rect 26 34 30 38
rect 50 34 54 38
<< ndcontact >>
rect 7 25 11 29
rect 18 18 22 22
rect 30 18 34 22
rect 40 18 44 22
rect 57 16 61 20
<< pdcontact >>
rect 13 43 17 47
rect 23 58 27 62
rect 37 43 41 47
rect 47 50 51 54
rect 47 43 51 47
rect 57 58 61 62
rect 57 51 61 55
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
<< psubstratepdiff >>
rect 0 2 64 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 64 2
rect 0 -3 64 -2
<< nsubstratendiff >>
rect 0 82 64 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 64 82
rect 0 77 64 78
<< labels >>
rlabel polycontact 52 36 52 36 6 an
rlabel polycontact 42 61 42 61 6 bn
rlabel metal1 4 56 4 56 6 b
rlabel metal1 20 32 20 32 6 a
rlabel metal1 9 35 9 35 6 bn
rlabel metal1 15 48 15 48 6 bn
rlabel metal1 12 60 12 60 6 b
rlabel metal1 32 6 32 6 6 vss
rlabel metal1 32 23 32 23 6 an
rlabel polycontact 28 36 28 36 6 a
rlabel metal1 32 74 32 74 6 vdd
rlabel metal1 44 20 44 20 6 z
rlabel metal1 39 40 39 40 6 an
rlabel metal1 52 28 52 28 6 z
rlabel metal1 52 44 52 44 6 z
rlabel metal1 45 36 45 36 6 an
rlabel metal1 60 36 60 36 6 z
rlabel metal1 59 56 59 56 6 bn
rlabel metal1 46 61 46 61 6 bn
<< end >>
