magic
tech scmos
timestamp 1180600814
<< checkpaint >>
rect -22 -22 142 122
<< ab >>
rect 0 0 120 100
<< pwell >>
rect -4 -4 124 48
<< nwell >>
rect -4 48 124 104
<< polysilicon >>
rect 13 94 15 98
rect 25 94 27 98
rect 37 85 39 89
rect 49 85 51 89
rect 61 85 63 89
rect 73 85 75 89
rect 87 85 89 89
rect 97 85 99 89
rect 107 85 109 89
rect 13 43 15 55
rect 25 43 27 55
rect 37 43 39 63
rect 49 43 51 63
rect 61 43 63 63
rect 73 43 75 61
rect 13 42 33 43
rect 13 38 28 42
rect 32 38 33 42
rect 13 37 33 38
rect 37 42 43 43
rect 37 38 38 42
rect 42 38 43 42
rect 37 37 43 38
rect 47 42 53 43
rect 47 38 48 42
rect 52 38 53 42
rect 47 37 53 38
rect 57 42 63 43
rect 57 38 58 42
rect 62 38 63 42
rect 57 37 63 38
rect 67 42 75 43
rect 67 38 68 42
rect 72 38 75 42
rect 87 53 89 56
rect 97 53 99 56
rect 87 52 93 53
rect 87 48 88 52
rect 92 48 93 52
rect 87 47 93 48
rect 97 52 103 53
rect 97 48 98 52
rect 102 48 103 52
rect 97 47 103 48
rect 87 39 89 47
rect 97 39 99 47
rect 67 37 75 38
rect 83 37 89 39
rect 95 37 99 39
rect 107 43 109 55
rect 107 42 113 43
rect 107 38 108 42
rect 112 38 113 42
rect 107 37 113 38
rect 13 34 15 37
rect 25 34 27 37
rect 39 33 41 37
rect 49 33 51 37
rect 59 33 61 37
rect 71 29 73 37
rect 83 25 85 37
rect 95 25 97 37
rect 107 25 109 37
rect 13 10 15 14
rect 25 10 27 14
rect 39 13 41 17
rect 49 13 51 17
rect 59 13 61 17
rect 71 13 73 17
rect 83 13 85 17
rect 95 13 97 17
rect 107 13 109 17
<< ndiffusion >>
rect 5 32 13 34
rect 5 28 6 32
rect 10 28 13 32
rect 5 22 13 28
rect 5 18 6 22
rect 10 18 13 22
rect 5 14 13 18
rect 15 32 25 34
rect 15 28 18 32
rect 22 28 25 32
rect 15 14 25 28
rect 27 33 37 34
rect 27 17 39 33
rect 41 17 49 33
rect 51 17 59 33
rect 61 29 66 33
rect 61 22 71 29
rect 61 18 64 22
rect 68 18 71 22
rect 61 17 71 18
rect 73 25 80 29
rect 73 22 83 25
rect 73 18 76 22
rect 80 18 83 22
rect 73 17 83 18
rect 85 17 95 25
rect 97 22 107 25
rect 97 18 100 22
rect 104 18 107 22
rect 97 17 107 18
rect 109 22 117 25
rect 109 18 112 22
rect 116 18 117 22
rect 109 17 117 18
rect 27 14 37 17
rect 31 12 37 14
rect 31 8 32 12
rect 36 8 37 12
rect 87 12 93 17
rect 31 7 37 8
rect 87 8 88 12
rect 92 8 93 12
rect 87 7 93 8
<< pdiffusion >>
rect 5 92 13 94
rect 5 88 6 92
rect 10 88 13 92
rect 5 82 13 88
rect 5 78 6 82
rect 10 78 13 82
rect 5 72 13 78
rect 5 68 6 72
rect 10 68 13 72
rect 5 62 13 68
rect 5 58 6 62
rect 10 58 13 62
rect 5 55 13 58
rect 15 82 25 94
rect 15 78 18 82
rect 22 78 25 82
rect 15 72 25 78
rect 15 68 18 72
rect 22 68 25 72
rect 15 62 25 68
rect 15 58 18 62
rect 22 58 25 62
rect 15 55 25 58
rect 27 85 34 94
rect 53 92 59 93
rect 53 88 54 92
rect 58 88 59 92
rect 53 85 59 88
rect 27 82 37 85
rect 27 78 30 82
rect 34 78 37 82
rect 27 63 37 78
rect 39 82 49 85
rect 39 78 42 82
rect 46 78 49 82
rect 39 63 49 78
rect 51 63 61 85
rect 63 82 73 85
rect 63 78 66 82
rect 70 78 73 82
rect 63 63 73 78
rect 27 55 34 63
rect 66 61 73 63
rect 75 72 87 85
rect 75 68 78 72
rect 82 68 87 72
rect 75 62 87 68
rect 75 61 78 62
rect 77 58 78 61
rect 82 58 87 62
rect 77 56 87 58
rect 89 56 97 85
rect 99 56 107 85
rect 102 55 107 56
rect 109 82 117 85
rect 109 78 112 82
rect 116 78 117 82
rect 109 55 117 78
<< metal1 >>
rect -2 96 122 100
rect -2 92 66 96
rect 70 92 78 96
rect 82 92 90 96
rect 94 92 102 96
rect 106 92 122 96
rect -2 88 6 92
rect 10 88 54 92
rect 58 88 122 92
rect 6 82 10 88
rect 6 72 10 78
rect 6 62 10 68
rect 6 57 10 58
rect 18 82 22 83
rect 18 72 22 78
rect 30 82 34 88
rect 41 78 42 82
rect 46 78 66 82
rect 70 78 112 82
rect 116 78 117 82
rect 30 77 34 78
rect 18 62 22 68
rect 6 32 10 33
rect 6 22 10 28
rect 6 12 10 18
rect 18 32 22 58
rect 18 17 22 28
rect 28 42 32 43
rect 28 22 32 38
rect 38 42 42 73
rect 38 27 42 38
rect 48 42 52 73
rect 48 27 52 38
rect 58 42 62 73
rect 58 37 62 38
rect 68 42 72 73
rect 68 37 72 38
rect 78 72 82 73
rect 78 62 82 68
rect 78 32 82 58
rect 64 28 82 32
rect 88 52 92 73
rect 64 22 68 28
rect 88 27 92 48
rect 98 52 102 73
rect 98 27 102 48
rect 108 42 112 73
rect 108 27 112 38
rect 112 22 116 23
rect 28 18 64 22
rect 75 18 76 22
rect 80 18 100 22
rect 104 18 105 22
rect 64 17 68 18
rect 112 12 116 18
rect -2 8 32 12
rect 36 10 88 12
rect 36 8 44 10
rect -2 6 44 8
rect 48 6 54 10
rect 58 6 64 10
rect 68 6 75 10
rect 79 8 88 10
rect 92 10 122 12
rect 92 8 102 10
rect 79 6 102 8
rect 106 6 110 10
rect 114 6 122 10
rect -2 0 122 6
<< ntransistor >>
rect 13 14 15 34
rect 25 14 27 34
rect 39 17 41 33
rect 49 17 51 33
rect 59 17 61 33
rect 71 17 73 29
rect 83 17 85 25
rect 95 17 97 25
rect 107 17 109 25
<< ptransistor >>
rect 13 55 15 94
rect 25 55 27 94
rect 37 63 39 85
rect 49 63 51 85
rect 61 63 63 85
rect 73 61 75 85
rect 87 56 89 85
rect 97 56 99 85
rect 107 55 109 85
<< polycontact >>
rect 28 38 32 42
rect 38 38 42 42
rect 48 38 52 42
rect 58 38 62 42
rect 68 38 72 42
rect 88 48 92 52
rect 98 48 102 52
rect 108 38 112 42
<< ndcontact >>
rect 6 28 10 32
rect 6 18 10 22
rect 18 28 22 32
rect 64 18 68 22
rect 76 18 80 22
rect 100 18 104 22
rect 112 18 116 22
rect 32 8 36 12
rect 88 8 92 12
<< pdcontact >>
rect 6 88 10 92
rect 6 78 10 82
rect 6 68 10 72
rect 6 58 10 62
rect 18 78 22 82
rect 18 68 22 72
rect 18 58 22 62
rect 54 88 58 92
rect 30 78 34 82
rect 42 78 46 82
rect 66 78 70 82
rect 78 68 82 72
rect 78 58 82 62
rect 112 78 116 82
<< psubstratepcontact >>
rect 44 6 48 10
rect 54 6 58 10
rect 64 6 68 10
rect 75 6 79 10
rect 102 6 106 10
rect 110 6 114 10
<< nsubstratencontact >>
rect 66 92 70 96
rect 78 92 82 96
rect 90 92 94 96
rect 102 92 106 96
<< psubstratepdiff >>
rect 43 10 80 11
rect 43 6 44 10
rect 48 6 54 10
rect 58 6 64 10
rect 68 6 75 10
rect 79 6 80 10
rect 101 10 115 11
rect 43 5 80 6
rect 101 6 102 10
rect 106 6 110 10
rect 114 6 115 10
rect 101 5 115 6
<< nsubstratendiff >>
rect 65 96 107 97
rect 65 92 66 96
rect 70 92 78 96
rect 82 92 90 96
rect 94 92 102 96
rect 106 92 107 96
rect 65 91 107 92
<< labels >>
rlabel metal1 20 50 20 50 6 q
rlabel metal1 40 50 40 50 6 i0
rlabel metal1 60 6 60 6 6 vss
rlabel metal1 50 50 50 50 6 i1
rlabel metal1 60 55 60 55 6 i2
rlabel metal1 60 94 60 94 6 vdd
rlabel metal1 70 55 70 55 6 i6
rlabel polycontact 90 50 90 50 6 i3
rlabel polycontact 100 50 100 50 6 i4
rlabel metal1 110 50 110 50 6 i5
<< end >>
