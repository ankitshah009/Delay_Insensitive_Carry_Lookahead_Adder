.subckt nd3v0x2 a b c vdd vss z
*   SPICE3 file   created from nd3v0x2.ext -      technology: scmos
m00 z      b      vdd    vdd p w=14u  l=2.3636u ad=65.3333p pd=20u      as=116.667p ps=33.3333u
m01 vdd    b      z      vdd p w=14u  l=2.3636u ad=116.667p pd=33.3333u as=65.3333p ps=20u
m02 z      c      vdd    vdd p w=28u  l=2.3636u ad=130.667p pd=40u      as=233.333p ps=66.6667u
m03 vdd    a      z      vdd p w=28u  l=2.3636u ad=233.333p pd=66.6667u as=130.667p ps=40u
m04 w1     a      vss    vss n w=14u  l=2.3636u ad=35p      pd=19u      as=126p     ps=46u
m05 w2     b      w1     vss n w=14u  l=2.3636u ad=35p      pd=19u      as=35p      ps=19u
m06 z      c      w2     vss n w=14u  l=2.3636u ad=56p      pd=22u      as=35p      ps=19u
m07 w3     c      z      vss n w=14u  l=2.3636u ad=35p      pd=19u      as=56p      ps=22u
m08 w4     b      w3     vss n w=14u  l=2.3636u ad=35p      pd=19u      as=35p      ps=19u
m09 vss    a      w4     vss n w=14u  l=2.3636u ad=126p     pd=46u      as=35p      ps=19u
C0  z      a      0.296f
C1  vss    c      0.022f
C2  z      b      0.142f
C3  a      c      0.191f
C4  vss    vdd    0.005f
C5  c      b      0.136f
C6  a      vdd    0.046f
C7  w4     a      0.007f
C8  b      vdd    0.043f
C9  w2     a      0.008f
C10 w1     z      0.015f
C11 vss    a      0.106f
C12 z      c      0.102f
C13 vss    b      0.028f
C14 a      b      0.206f
C15 z      vdd    0.385f
C16 c      vdd    0.021f
C17 w3     a      0.007f
C18 w2     z      0.010f
C19 vss    z      0.240f
C21 z      vss    0.013f
C22 a      vss    0.033f
C23 c      vss    0.022f
C24 b      vss    0.047f
.ends
