.subckt nr2av0x3 a b vdd vss z
*   SPICE3 file   created from nr2av0x3.ext -      technology: scmos
m00 w1     b      z      vdd p w=25u  l=2.3636u ad=62.5p    pd=30u      as=117p     ps=43.3333u
m01 vdd    an     w1     vdd p w=25u  l=2.3636u ad=106.796p pd=33.9806u as=62.5p    ps=30u
m02 w2     an     vdd    vdd p w=25u  l=2.3636u ad=62.5p    pd=30u      as=106.796p ps=33.9806u
m03 z      b      w2     vdd p w=25u  l=2.3636u ad=117p     pd=43.3333u as=62.5p    ps=30u
m04 w3     b      z      vdd p w=25u  l=2.3636u ad=62.5p    pd=30u      as=117p     ps=43.3333u
m05 vdd    an     w3     vdd p w=25u  l=2.3636u ad=106.796p pd=33.9806u as=62.5p    ps=30u
m06 an     a      vdd    vdd p w=28u  l=2.3636u ad=166p     pd=70u      as=119.612p ps=38.0583u
m07 z      b      vss    vss n w=20u  l=2.3636u ad=80p      pd=28u      as=177.407p ps=62.963u
m08 vss    an     z      vss n w=20u  l=2.3636u ad=177.407p pd=62.963u  as=80p      ps=28u
m09 an     a      vss    vss n w=14u  l=2.3636u ad=98p      pd=42u      as=124.185p ps=44.0741u
C0  z      b      0.334f
C1  a      an     0.248f
C2  w1     vdd    0.005f
C3  an     b      0.324f
C4  a      vdd    0.023f
C5  vss    z      0.060f
C6  b      vdd    0.042f
C7  w3     a      0.002f
C8  vss    an     0.145f
C9  w2     z      0.010f
C10 vss    vdd    0.005f
C11 w2     vdd    0.005f
C12 z      an     0.066f
C13 a      b      0.068f
C14 z      vdd    0.261f
C15 an     vdd    0.043f
C16 vss    a      0.026f
C17 w3     z      0.003f
C18 w1     z      0.010f
C19 vss    b      0.263f
C20 w3     vdd    0.005f
C21 z      a      0.015f
C23 z      vss    0.006f
C24 a      vss    0.019f
C25 an     vss    0.053f
C26 b      vss    0.049f
.ends
