.subckt xaon21v0x1 a1 a2 b vdd vss z
*   SPICE3 file   created from xaon21v0x1.ext -      technology: scmos
m00 z      an     bn     vdd p w=28u  l=2.3636u ad=112p     pd=36u      as=132p     ps=57u
m01 an     bn     z      vdd p w=28u  l=2.3636u ad=125.831p pd=47.9036u as=112p     ps=36u
m02 vdd    a2     an     vdd p w=27u  l=2.3636u ad=193.554p pd=71.5663u as=121.337p ps=46.1928u
m03 vdd    a1     an     vdd p w=28u  l=2.3636u ad=200.723p pd=74.2169u as=125.831p ps=47.9036u
m04 bn     b      vdd    vdd p w=14u  l=2.3636u ad=66p      pd=28.5u    as=100.361p ps=37.1084u
m05 vdd    b      bn     vdd p w=14u  l=2.3636u ad=100.361p pd=37.1084u as=66p      ps=28.5u
m06 w1     an     vss    vss n w=13u  l=2.3636u ad=32.5p    pd=18u      as=123.825p ps=39u
m07 z      bn     w1     vss n w=13u  l=2.3636u ad=54.4375p pd=21.9375u as=32.5p    ps=18u
m08 an     b      z      vss n w=19u  l=2.3636u ad=78.8788p pd=31.0909u as=79.5625p ps=32.0625u
m09 w2     a2     an     vss n w=14u  l=2.3636u ad=35p      pd=19u      as=58.1212p ps=22.9091u
m10 vss    a1     w2     vss n w=14u  l=2.3636u ad=133.35p  pd=42u      as=35p      ps=19u
m11 bn     b      vss    vss n w=13u  l=2.3636u ad=77p      pd=40u      as=123.825p ps=39u
C0  vdd    a1     0.017f
C1  b      bn     0.185f
C2  vss    an     0.106f
C3  z      a2     0.027f
C4  vdd    bn     0.463f
C5  z      an     0.505f
C6  a1     a2     0.233f
C7  a1     an     0.038f
C8  a2     bn     0.227f
C9  vss    z      0.188f
C10 bn     an     0.860f
C11 b      vdd    0.124f
C12 vss    a1     0.178f
C13 z      a1     0.011f
C14 b      a2     0.049f
C15 vss    bn     0.066f
C16 w1     an     0.007f
C17 b      an     0.015f
C18 z      bn     0.270f
C19 vdd    a2     0.017f
C20 vdd    an     0.119f
C21 a1     bn     0.149f
C22 w1     z      0.010f
C23 vss    b      0.020f
C24 a2     an     0.168f
C25 w2     a2     0.021f
C26 b      z      0.007f
C27 b      a1     0.054f
C28 z      vdd    0.043f
C29 vss    a2     0.055f
C31 b      vss    0.047f
C32 z      vss    0.012f
C34 a1     vss    0.016f
C35 a2     vss    0.023f
C36 bn     vss    0.028f
C37 an     vss    0.018f
.ends
