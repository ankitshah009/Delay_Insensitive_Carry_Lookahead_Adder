.subckt iv1v0x12 a vdd vss z
*   SPICE3 file   created from iv1v0x12.ext -      technology: scmos
m00 z      a      vdd    vdd p w=28u  l=2.3636u ad=176p     pd=50u      as=196p     ps=70u
m01 vdd    a      z      vdd p w=28u  l=2.3636u ad=196p     pd=70u      as=176p     ps=50u
m02 z      a      vdd    vdd p w=28u  l=2.3636u ad=176p     pd=50u      as=196p     ps=70u
m03 vdd    a      z      vdd p w=28u  l=2.3636u ad=196p     pd=70u      as=176p     ps=50u
m04 z      a      vdd    vdd p w=28u  l=2.3636u ad=176p     pd=50u      as=196p     ps=70u
m05 vdd    a      z      vdd p w=28u  l=2.3636u ad=196p     pd=70u      as=176p     ps=50u
m06 z      a      vss    vss n w=20u  l=2.3636u ad=136p     pd=42u      as=140p     ps=54u
m07 vss    a      z      vss n w=20u  l=2.3636u ad=140p     pd=54u      as=136p     ps=42u
m08 z      a      vss    vss n w=20u  l=2.3636u ad=136p     pd=42u      as=140p     ps=54u
m09 vss    a      z      vss n w=20u  l=2.3636u ad=140p     pd=54u      as=136p     ps=42u
m10 z      a      vss    vss n w=20u  l=2.3636u ad=136p     pd=42u      as=140p     ps=54u
m11 vss    a      z      vss n w=20u  l=2.3636u ad=140p     pd=54u      as=136p     ps=42u
C0  z      vdd    0.377f
C1  vss    z      0.434f
C2  vss    vdd    0.019f
C3  z      a      0.792f
C4  a      vdd    0.488f
C5  vss    a      0.224f
C7  z      vss    0.014f
C8  a      vss    0.283f
.ends
