magic
tech scmos
timestamp 1179385640
<< checkpaint >>
rect -22 -25 110 105
<< ab >>
rect 0 0 88 80
<< pwell >>
rect -4 -7 92 36
<< nwell >>
rect -4 36 92 87
<< polysilicon >>
rect 9 69 11 74
rect 19 69 21 74
rect 39 69 41 74
rect 46 69 48 74
rect 56 69 58 74
rect 66 69 68 74
rect 76 69 78 74
rect 9 39 11 42
rect 19 39 21 42
rect 39 39 41 42
rect 46 39 48 42
rect 56 39 58 42
rect 66 39 68 42
rect 76 39 78 42
rect 5 38 11 39
rect 5 34 6 38
rect 10 34 11 38
rect 5 33 11 34
rect 17 38 23 39
rect 17 34 18 38
rect 22 34 23 38
rect 17 33 23 34
rect 32 38 42 39
rect 32 34 33 38
rect 37 34 42 38
rect 46 36 49 39
rect 32 33 42 34
rect 9 30 11 33
rect 19 30 21 33
rect 40 30 42 33
rect 47 30 49 36
rect 55 38 61 39
rect 55 34 56 38
rect 60 34 61 38
rect 55 33 61 34
rect 65 38 71 39
rect 65 34 66 38
rect 70 34 71 38
rect 65 33 71 34
rect 76 38 86 39
rect 76 34 81 38
rect 85 34 86 38
rect 76 33 86 34
rect 57 30 59 33
rect 67 30 69 33
rect 77 30 79 33
rect 9 11 11 16
rect 19 11 21 16
rect 40 13 42 18
rect 47 8 49 18
rect 57 12 59 16
rect 67 8 69 16
rect 77 11 79 16
rect 47 6 69 8
<< ndiffusion >>
rect 2 29 9 30
rect 2 25 3 29
rect 7 25 9 29
rect 2 22 9 25
rect 2 18 3 22
rect 7 18 9 22
rect 2 16 9 18
rect 11 21 19 30
rect 11 17 13 21
rect 17 17 19 21
rect 11 16 19 17
rect 21 22 26 30
rect 21 21 28 22
rect 21 17 23 21
rect 27 17 28 21
rect 21 16 28 17
rect 32 18 40 30
rect 42 18 47 30
rect 49 29 57 30
rect 49 25 51 29
rect 55 25 57 29
rect 49 18 57 25
rect 32 12 38 18
rect 32 8 33 12
rect 37 8 38 12
rect 32 7 38 8
rect 52 16 57 18
rect 59 21 67 30
rect 59 17 61 21
rect 65 17 67 21
rect 59 16 67 17
rect 69 21 77 30
rect 69 17 71 21
rect 75 17 77 21
rect 69 16 77 17
rect 79 29 86 30
rect 79 25 81 29
rect 85 25 86 29
rect 79 22 86 25
rect 79 18 81 22
rect 85 18 86 22
rect 79 16 86 18
<< pdiffusion >>
rect 4 63 9 69
rect 2 62 9 63
rect 2 58 3 62
rect 7 58 9 62
rect 2 55 9 58
rect 2 51 3 55
rect 7 51 9 55
rect 2 50 9 51
rect 4 42 9 50
rect 11 68 19 69
rect 11 64 13 68
rect 17 64 19 68
rect 11 61 19 64
rect 11 57 13 61
rect 17 57 19 61
rect 11 42 19 57
rect 21 63 26 69
rect 32 68 39 69
rect 32 64 33 68
rect 37 64 39 68
rect 21 62 28 63
rect 21 58 23 62
rect 27 58 28 62
rect 21 55 28 58
rect 21 51 23 55
rect 27 51 28 55
rect 21 50 28 51
rect 32 61 39 64
rect 32 57 33 61
rect 37 57 39 61
rect 21 42 26 50
rect 32 42 39 57
rect 41 42 46 69
rect 48 49 56 69
rect 48 45 50 49
rect 54 45 56 49
rect 48 42 56 45
rect 58 63 66 69
rect 58 59 60 63
rect 64 59 66 63
rect 58 42 66 59
rect 68 68 76 69
rect 68 64 70 68
rect 74 64 76 68
rect 68 61 76 64
rect 68 57 70 61
rect 74 57 76 61
rect 68 42 76 57
rect 78 63 83 69
rect 78 62 85 63
rect 78 58 80 62
rect 84 58 85 62
rect 78 55 85 58
rect 78 51 80 55
rect 84 51 85 55
rect 78 50 85 51
rect 78 42 83 50
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect -2 68 90 78
rect 12 64 13 68
rect 17 64 18 68
rect 3 62 7 63
rect 3 55 7 58
rect 12 61 18 64
rect 32 64 33 68
rect 37 64 38 68
rect 12 57 13 61
rect 17 57 18 61
rect 23 62 27 63
rect 23 55 27 58
rect 32 61 38 64
rect 69 64 70 68
rect 74 64 75 68
rect 32 57 33 61
rect 37 57 38 61
rect 42 59 60 63
rect 64 59 65 63
rect 69 61 75 64
rect 7 51 17 54
rect 3 50 17 51
rect 42 54 46 59
rect 69 57 70 61
rect 74 57 75 61
rect 80 62 84 63
rect 80 55 84 58
rect 27 51 46 54
rect 23 50 46 51
rect 13 47 17 50
rect 50 49 54 55
rect 2 39 6 47
rect 13 43 22 47
rect 2 38 14 39
rect 2 34 6 38
rect 10 34 14 38
rect 2 33 14 34
rect 18 38 22 43
rect 42 45 50 47
rect 42 43 54 45
rect 22 34 33 38
rect 37 34 38 38
rect 18 30 22 34
rect 3 29 22 30
rect 7 26 22 29
rect 42 29 46 43
rect 58 39 62 55
rect 50 38 62 39
rect 50 34 56 38
rect 60 34 62 38
rect 50 33 62 34
rect 66 51 80 54
rect 66 50 84 51
rect 66 38 70 50
rect 82 39 86 47
rect 66 30 70 34
rect 74 38 86 39
rect 74 34 81 38
rect 85 34 86 38
rect 74 33 86 34
rect 66 29 85 30
rect 42 25 51 29
rect 55 25 56 29
rect 66 26 81 29
rect 3 22 7 25
rect 81 22 85 25
rect 3 17 7 18
rect 12 17 13 21
rect 17 17 18 21
rect 22 17 23 21
rect 27 17 61 21
rect 65 17 66 21
rect 70 17 71 21
rect 75 17 76 21
rect 81 17 85 18
rect 12 12 18 17
rect 70 12 76 17
rect -2 8 33 12
rect 37 8 90 12
rect -2 2 90 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
<< ntransistor >>
rect 9 16 11 30
rect 19 16 21 30
rect 40 18 42 30
rect 47 18 49 30
rect 57 16 59 30
rect 67 16 69 30
rect 77 16 79 30
<< ptransistor >>
rect 9 42 11 69
rect 19 42 21 69
rect 39 42 41 69
rect 46 42 48 69
rect 56 42 58 69
rect 66 42 68 69
rect 76 42 78 69
<< polycontact >>
rect 6 34 10 38
rect 18 34 22 38
rect 33 34 37 38
rect 56 34 60 38
rect 66 34 70 38
rect 81 34 85 38
<< ndcontact >>
rect 3 25 7 29
rect 3 18 7 22
rect 13 17 17 21
rect 23 17 27 21
rect 51 25 55 29
rect 33 8 37 12
rect 61 17 65 21
rect 71 17 75 21
rect 81 25 85 29
rect 81 18 85 22
<< pdcontact >>
rect 3 58 7 62
rect 3 51 7 55
rect 13 64 17 68
rect 13 57 17 61
rect 33 64 37 68
rect 23 58 27 62
rect 23 51 27 55
rect 33 57 37 61
rect 50 45 54 49
rect 60 59 64 63
rect 70 64 74 68
rect 70 57 74 61
rect 80 58 84 62
rect 80 51 84 55
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
<< psubstratepdiff >>
rect 0 2 88 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 88 2
rect 0 -3 88 -2
<< nsubstratendiff >>
rect 0 82 88 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 88 82
rect 0 77 88 78
<< labels >>
rlabel polysilicon 20 42 20 42 6 an
rlabel polysilicon 37 36 37 36 6 an
rlabel polycontact 68 36 68 36 6 bn
rlabel metal1 5 23 5 23 6 an
rlabel metal1 4 40 4 40 6 a
rlabel metal1 12 36 12 36 6 a
rlabel metal1 5 56 5 56 6 an
rlabel metal1 25 56 25 56 6 n1
rlabel metal1 44 6 44 6 6 vss
rlabel metal1 28 36 28 36 6 an
rlabel metal1 44 36 44 36 6 z
rlabel metal1 44 74 44 74 6 vdd
rlabel metal1 44 19 44 19 6 n3
rlabel metal1 52 36 52 36 6 c
rlabel metal1 60 44 60 44 6 c
rlabel metal1 52 52 52 52 6 z
rlabel metal1 68 40 68 40 6 bn
rlabel metal1 53 61 53 61 6 n1
rlabel metal1 84 40 84 40 6 b
rlabel metal1 76 36 76 36 6 b
<< end >>
