magic
tech scmos
timestamp 1179387324
<< checkpaint >>
rect -22 -25 30 105
<< ab >>
rect 0 0 8 80
<< pwell >>
rect -4 -7 12 36
<< nwell >>
rect -4 36 12 87
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect -2 68 10 78
rect -2 2 10 12
rect -2 -2 2 2
rect 6 -2 10 2
<< psubstratepcontact >>
rect 2 -2 6 2
<< nsubstratencontact >>
rect 2 78 6 82
<< psubstratepdiff >>
rect 0 2 8 3
rect 0 -2 2 2
rect 6 -2 8 2
rect 0 -3 8 -2
<< nsubstratendiff >>
rect 0 82 8 83
rect 0 78 2 82
rect 6 78 8 82
rect 0 77 8 78
<< labels >>
rlabel metal1 4 6 4 6 6 vss
rlabel metal1 4 74 4 74 6 vdd
<< end >>
