magic
tech scmos
timestamp 1179386320
<< checkpaint >>
rect -22 -25 78 105
<< ab >>
rect 0 0 56 80
<< pwell >>
rect -4 -7 60 36
<< nwell >>
rect -4 36 60 87
<< polysilicon >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 62 31 67
rect 39 62 41 67
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 39 39 41 42
rect 9 38 15 39
rect 9 34 10 38
rect 14 34 15 38
rect 9 33 15 34
rect 19 38 31 39
rect 19 34 26 38
rect 30 34 31 38
rect 19 33 31 34
rect 12 30 14 33
rect 19 30 21 33
rect 29 30 31 33
rect 36 38 42 39
rect 36 34 37 38
rect 41 34 42 38
rect 36 33 42 34
rect 36 30 38 33
rect 12 6 14 10
rect 19 6 21 10
rect 29 6 31 10
rect 36 6 38 10
<< ndiffusion >>
rect 3 12 12 30
rect 3 8 5 12
rect 9 10 12 12
rect 14 10 19 30
rect 21 22 29 30
rect 21 18 23 22
rect 27 18 29 22
rect 21 10 29 18
rect 31 10 36 30
rect 38 22 46 30
rect 38 18 41 22
rect 45 18 46 22
rect 38 17 46 18
rect 38 10 43 17
rect 9 8 10 10
rect 3 7 10 8
<< pdiffusion >>
rect 2 69 9 70
rect 2 65 3 69
rect 7 65 9 69
rect 2 62 9 65
rect 2 58 3 62
rect 7 58 9 62
rect 2 42 9 58
rect 11 54 19 70
rect 11 50 13 54
rect 17 50 19 54
rect 11 47 19 50
rect 11 43 13 47
rect 17 43 19 47
rect 11 42 19 43
rect 21 62 27 70
rect 21 61 29 62
rect 21 57 23 61
rect 27 57 29 61
rect 21 42 29 57
rect 31 61 39 62
rect 31 57 33 61
rect 37 57 39 61
rect 31 54 39 57
rect 31 50 33 54
rect 37 50 39 54
rect 31 42 39 50
rect 41 61 49 62
rect 41 57 43 61
rect 47 57 49 61
rect 41 54 49 57
rect 41 50 43 54
rect 47 50 49 54
rect 41 42 49 50
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect -2 69 58 78
rect -2 68 3 69
rect 2 65 3 68
rect 7 68 58 69
rect 7 65 8 68
rect 2 62 8 65
rect 2 58 3 62
rect 7 58 8 62
rect 22 61 28 68
rect 22 57 23 61
rect 27 57 28 61
rect 33 61 38 63
rect 37 57 38 61
rect 33 54 38 57
rect 12 50 13 54
rect 17 50 33 54
rect 37 50 38 54
rect 42 61 48 68
rect 42 57 43 61
rect 47 57 48 61
rect 42 54 48 57
rect 42 50 43 54
rect 47 50 48 54
rect 12 47 18 50
rect 2 43 13 47
rect 17 43 18 47
rect 2 22 6 43
rect 25 42 39 46
rect 10 38 14 39
rect 25 38 31 42
rect 25 34 26 38
rect 30 34 31 38
rect 36 34 37 38
rect 41 34 42 38
rect 10 30 14 34
rect 36 30 42 34
rect 10 26 47 30
rect 2 18 23 22
rect 27 18 31 22
rect 40 18 41 22
rect 45 18 46 22
rect 40 12 46 18
rect -2 8 5 12
rect 9 8 58 12
rect -2 2 58 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
<< ntransistor >>
rect 12 10 14 30
rect 19 10 21 30
rect 29 10 31 30
rect 36 10 38 30
<< ptransistor >>
rect 9 42 11 70
rect 19 42 21 70
rect 29 42 31 62
rect 39 42 41 62
<< polycontact >>
rect 10 34 14 38
rect 26 34 30 38
rect 37 34 41 38
<< ndcontact >>
rect 5 8 9 12
rect 23 18 27 22
rect 41 18 45 22
<< pdcontact >>
rect 3 65 7 69
rect 3 58 7 62
rect 13 50 17 54
rect 13 43 17 47
rect 23 57 27 61
rect 33 57 37 61
rect 33 50 37 54
rect 43 57 47 61
rect 43 50 47 54
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
<< psubstratepdiff >>
rect 0 2 56 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 56 2
rect 0 -3 56 -2
<< nsubstratendiff >>
rect 0 82 56 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 56 82
rect 0 77 56 78
<< labels >>
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 20 12 20 6 z
rlabel polycontact 12 36 12 36 6 a
rlabel metal1 28 6 28 6 6 vss
rlabel metal1 20 20 20 20 6 z
rlabel metal1 20 28 20 28 6 a
rlabel metal1 28 28 28 28 6 a
rlabel metal1 28 20 28 20 6 z
rlabel metal1 28 40 28 40 6 b
rlabel metal1 28 52 28 52 6 z
rlabel metal1 20 52 20 52 6 z
rlabel metal1 28 74 28 74 6 vdd
rlabel metal1 36 28 36 28 6 a
rlabel metal1 44 28 44 28 6 a
rlabel metal1 36 44 36 44 6 b
rlabel pdcontact 36 60 36 60 6 z
<< end >>
