.subckt cgi2v0x2 a b c vdd vss z
*   SPICE3 file   created from cgi2v0x2.ext -      technology: scmos
m00 n1     a      vdd    vdd p w=28u  l=2.3636u ad=112p     pd=36u      as=158.667p ps=48.6667u
m01 z      c      n1     vdd p w=28u  l=2.3636u ad=112p     pd=36u      as=112p     ps=36u
m02 n1     c      z      vdd p w=28u  l=2.3636u ad=112p     pd=36u      as=112p     ps=36u
m03 vdd    a      n1     vdd p w=28u  l=2.3636u ad=158.667p pd=48.6667u as=112p     ps=36u
m04 w1     a      vdd    vdd p w=28u  l=2.3636u ad=70p      pd=33u      as=158.667p ps=48.6667u
m05 z      b      w1     vdd p w=28u  l=2.3636u ad=112p     pd=36u      as=70p      ps=33u
m06 w2     b      z      vdd p w=28u  l=2.3636u ad=70p      pd=33u      as=112p     ps=36u
m07 vdd    a      w2     vdd p w=28u  l=2.3636u ad=158.667p pd=48.6667u as=70p      ps=33u
m08 n1     b      vdd    vdd p w=28u  l=2.3636u ad=112p     pd=36u      as=158.667p ps=48.6667u
m09 vdd    b      n1     vdd p w=28u  l=2.3636u ad=158.667p pd=48.6667u as=112p     ps=36u
m10 n3     a      vss    vss n w=14u  l=2.3636u ad=56p      pd=22u      as=97.3333p ps=36u
m11 z      c      n3     vss n w=14u  l=2.3636u ad=57.5p    pd=23.5u    as=56p      ps=22u
m12 n3     c      z      vss n w=14u  l=2.3636u ad=56p      pd=22u      as=57.5p    ps=23.5u
m13 vss    a      n3     vss n w=14u  l=2.3636u ad=97.3333p pd=36u      as=56p      ps=22u
m14 w3     a      vss    vss n w=17u  l=2.3636u ad=42.5p    pd=22u      as=118.19p  ps=43.7143u
m15 z      b      w3     vss n w=17u  l=2.3636u ad=69.8214p pd=28.5357u as=42.5p    ps=22u
m16 w4     b      z      vss n w=11u  l=2.3636u ad=27.5p    pd=16u      as=45.1786p ps=18.4643u
m17 vss    a      w4     vss n w=11u  l=2.3636u ad=76.4762p pd=28.2857u as=27.5p    ps=16u
m18 n3     b      vss    vss n w=14u  l=2.3636u ad=56p      pd=22u      as=97.3333p ps=36u
m19 vss    b      n3     vss n w=14u  l=2.3636u ad=97.3333p pd=36u      as=56p      ps=22u
C0  w1     z      0.007f
C1  w2     n1     0.010f
C2  vss    z      0.160f
C3  n3     n1     0.069f
C4  z      n1     0.155f
C5  n3     c      0.043f
C6  vss    b      0.099f
C7  n1     b      0.062f
C8  w1     a      0.010f
C9  w2     vdd    0.005f
C10 z      c      0.248f
C11 vss    a      0.111f
C12 w4     n3     0.005f
C13 n1     a      0.588f
C14 z      vdd    0.092f
C15 b      c      0.026f
C16 b      vdd    0.044f
C17 c      a      0.368f
C18 n3     z      0.395f
C19 w4     b      0.008f
C20 a      vdd    0.309f
C21 w1     n1     0.010f
C22 vss    n1     0.003f
C23 n3     b      0.188f
C24 z      b      0.116f
C25 w2     a      0.016f
C26 n3     a      0.110f
C27 vss    c      0.024f
C28 w1     vdd    0.005f
C29 z      a      0.606f
C30 n1     c      0.048f
C31 vss    vdd    0.009f
C32 w3     n3     0.010f
C33 n1     vdd    0.597f
C34 b      a      0.448f
C35 w3     z      0.007f
C36 n3     vss    0.595f
C37 c      vdd    0.024f
C38 n3     vss    0.002f
C40 z      vss    0.005f
C41 b      vss    0.062f
C42 c      vss    0.035f
C43 a      vss    0.069f
.ends
