.subckt an4v0x1 a b c d vdd vss z
*   SPICE3 file   created from an4v0x1.ext -      technology: scmos
m00 vdd    zn     z      vdd p w=18u  l=2.3636u ad=113.4p   pd=42.1714u as=116p     ps=50u
m01 zn     a      vdd    vdd p w=13u  l=2.3636u ad=52p      pd=21u      as=81.9p    ps=30.4571u
m02 vdd    b      zn     vdd p w=13u  l=2.3636u ad=81.9p    pd=30.4571u as=52p      ps=21u
m03 zn     c      vdd    vdd p w=13u  l=2.3636u ad=52p      pd=21u      as=81.9p    ps=30.4571u
m04 vdd    d      zn     vdd p w=13u  l=2.3636u ad=81.9p    pd=30.4571u as=52p      ps=21u
m05 vss    zn     z      vss n w=9u   l=2.3636u ad=86.04p   pd=24.48u   as=57p      ps=32u
m06 w1     a      vss    vss n w=16u  l=2.3636u ad=40p      pd=21u      as=152.96p  ps=43.52u
m07 w2     b      w1     vss n w=16u  l=2.3636u ad=40p      pd=21u      as=40p      ps=21u
m08 w3     c      w2     vss n w=16u  l=2.3636u ad=40p      pd=21u      as=40p      ps=21u
m09 zn     d      w3     vss n w=16u  l=2.3636u ad=92p      pd=46u      as=40p      ps=21u
C0  z      zn     0.268f
C1  w3     a      0.005f
C2  vss    d      0.051f
C3  z      c      0.011f
C4  vss    b      0.017f
C5  zn     d      0.103f
C6  w1     a      0.005f
C7  vss    vdd    0.003f
C8  d      c      0.209f
C9  zn     b      0.140f
C10 z      a      0.020f
C11 w2     vss    0.003f
C12 d      a      0.101f
C13 c      b      0.192f
C14 zn     vdd    0.344f
C15 w2     zn     0.010f
C16 b      a      0.167f
C17 c      vdd    0.035f
C18 vss    zn     0.271f
C19 a      vdd    0.027f
C20 vss    c      0.017f
C21 z      d      0.007f
C22 w2     a      0.005f
C23 zn     c      0.102f
C24 z      b      0.017f
C25 vss    a      0.056f
C26 w3     vss    0.003f
C27 z      vdd    0.054f
C28 d      b      0.036f
C29 zn     a      0.319f
C30 w1     vss    0.003f
C31 w3     zn     0.010f
C32 c      a      0.055f
C33 d      vdd    0.029f
C34 vss    z      0.089f
C35 w1     zn     0.010f
C36 b      vdd    0.038f
C38 z      vss    0.013f
C39 zn     vss    0.023f
C40 d      vss    0.039f
C41 c      vss    0.025f
C42 b      vss    0.026f
C43 a      vss    0.027f
.ends
