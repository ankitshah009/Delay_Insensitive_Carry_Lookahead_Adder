.subckt no3_x4 i0 i1 i2 nq vdd vss
*   SPICE3 file   created from no3_x4.ext -      technology: scmos
m00 w1     i2     w2     vdd p w=38u  l=2.3636u ad=114p     pd=44u      as=304p     ps=92u
m01 w3     i1     w1     vdd p w=38u  l=2.3636u ad=114p     pd=44u      as=114p     ps=44u
m02 vdd    i0     w3     vdd p w=38u  l=2.3636u ad=248.397p pd=57u      as=114p     ps=44u
m03 nq     w4     vdd    vdd p w=39u  l=2.3636u ad=195p     pd=49u      as=254.934p ps=58.5u
m04 vdd    w4     nq     vdd p w=39u  l=2.3636u ad=254.934p pd=58.5u    as=195p     ps=49u
m05 w4     w2     vdd    vdd p w=20u  l=2.3636u ad=160p     pd=56u      as=130.735p ps=30u
m06 vss    i2     w2     vss n w=10u  l=2.3636u ad=58.718p  pd=23.3333u as=61p      ps=26u
m07 w2     i1     vss    vss n w=10u  l=2.3636u ad=61p      pd=26u      as=58.718p  ps=23.3333u
m08 vss    i0     w2     vss n w=10u  l=2.3636u ad=58.718p  pd=23.3333u as=61p      ps=26u
m09 nq     w4     vss    vss n w=19u  l=2.3636u ad=95p      pd=29u      as=111.564p ps=44.3333u
m10 vss    w4     nq     vss n w=19u  l=2.3636u ad=111.564p pd=44.3333u as=95p      ps=29u
m11 w4     w2     vss    vss n w=10u  l=2.3636u ad=80p      pd=36u      as=58.718p  ps=23.3333u
C0  vss    nq     0.058f
C1  vdd    i0     0.035f
C2  w2     i1     0.171f
C3  w4     i1     0.043f
C4  vdd    i2     0.013f
C5  nq     w2     0.401f
C6  i0     i2     0.121f
C7  w1     w2     0.012f
C8  nq     w4     0.106f
C9  vss    i0     0.011f
C10 w3     vdd    0.011f
C11 vss    i2     0.011f
C12 w2     vdd    0.460f
C13 nq     i1     0.054f
C14 vdd    w4     0.016f
C15 w2     i0     0.337f
C16 w1     i1     0.013f
C17 vdd    i1     0.013f
C18 w4     i0     0.123f
C19 w2     i2     0.135f
C20 vss    w2     0.238f
C21 i0     i1     0.303f
C22 w4     i2     0.025f
C23 vss    w4     0.051f
C24 w3     w2     0.012f
C25 nq     vdd    0.027f
C26 i1     i2     0.344f
C27 nq     i0     0.087f
C28 w1     vdd    0.011f
C29 vss    i1     0.011f
C30 w2     w4     0.288f
C31 nq     i2     0.039f
C32 w3     i1     0.013f
C34 nq     vss    0.012f
C35 w2     vss    0.041f
C37 w4     vss    0.071f
C38 i0     vss    0.034f
C39 i1     vss    0.029f
C40 i2     vss    0.030f
.ends
