.subckt nr2v0x1 a b vdd vss z
*   SPICE3 file   created from nr2v0x1.ext -      technology: scmos
m00 w1     a      vdd    vdd p w=28u  l=2.3636u ad=176p     pd=50u      as=196p     ps=70u
m01 z      b      w1     vdd p w=28u  l=2.3636u ad=196p     pd=70u      as=176p     ps=50u
m02 z      a      vss    vss n w=20u  l=2.3636u ad=136p     pd=42u      as=140p     ps=54u
m03 vss    b      z      vss n w=20u  l=2.3636u ad=140p     pd=54u      as=136p     ps=42u
C0  vss    z      0.079f
C1  z      b      0.222f
C2  vss    vdd    0.004f
C3  z      a      0.174f
C4  b      vdd    0.010f
C5  a      vdd    0.041f
C6  vss    b      0.047f
C7  vss    a      0.031f
C8  z      w1     0.023f
C9  b      a      0.100f
C10 z      vdd    0.021f
C11 w1     vdd    0.010f
C13 z      vss    0.006f
C14 b      vss    0.045f
C15 a      vss    0.045f
.ends
