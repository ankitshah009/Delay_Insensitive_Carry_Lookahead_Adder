.subckt mxi2v2x05 a0 a1 s vdd vss z
*   SPICE3 file   created from mxi2v2x05.ext -      technology: scmos
m00 sn     s      vdd    vdd p w=6u   l=2.3636u ad=42p      pd=26u      as=70.4p    ps=27.6u
m01 a0n    a0     vdd    vdd p w=12u  l=2.3636u ad=48p      pd=20u      as=140.8p   ps=55.2u
m02 z      s      a0n    vdd p w=12u  l=2.3636u ad=48p      pd=20u      as=48p      ps=20u
m03 a1n    sn     z      vdd p w=12u  l=2.3636u ad=48p      pd=20u      as=48p      ps=20u
m04 vdd    a1     a1n    vdd p w=12u  l=2.3636u ad=140.8p   pd=55.2u    as=48p      ps=20u
m05 a0n    a0     vss    vss n w=6u   l=2.3636u ad=24p      pd=14u      as=44.6667p ps=23.3333u
m06 z      sn     a0n    vss n w=6u   l=2.3636u ad=24p      pd=14u      as=24p      ps=14u
m07 a1n    s      z      vss n w=6u   l=2.3636u ad=24p      pd=14u      as=24p      ps=14u
m08 vss    a1     a1n    vss n w=6u   l=2.3636u ad=44.6667p pd=23.3333u as=24p      ps=14u
m09 sn     s      vss    vss n w=6u   l=2.3636u ad=42p      pd=26u      as=44.6667p ps=23.3333u
C0  s      vdd    0.064f
C1  vss    a0     0.023f
C2  z      a1     0.037f
C3  a1n    sn     0.057f
C4  a0n    sn     0.038f
C5  z      a0     0.038f
C6  a1n    s      0.018f
C7  vss    vdd    0.007f
C8  z      vdd    0.012f
C9  a0n    s      0.017f
C10 a1     a0     0.022f
C11 vss    a1n    0.068f
C12 a1     vdd    0.012f
C13 sn     s      0.332f
C14 vss    a0n    0.067f
C15 a1n    z      0.293f
C16 a0     vdd    0.075f
C17 z      a0n    0.172f
C18 a1n    a1     0.094f
C19 vss    sn     0.026f
C20 z      sn     0.065f
C21 a0n    a1     0.020f
C22 a1n    a0     0.016f
C23 vss    s      0.027f
C24 a1     sn     0.137f
C25 z      s      0.038f
C26 a1n    vdd    0.009f
C27 a0n    a0     0.078f
C28 a1     s      0.137f
C29 a0n    vdd    0.010f
C30 sn     a0     0.048f
C31 vss    z      0.061f
C32 sn     vdd    0.216f
C33 a0     s      0.042f
C34 a1n    a0n    0.068f
C35 vss    a1     0.085f
C37 a1n    vss    0.009f
C38 z      vss    0.009f
C39 a0n    vss    0.009f
C40 a1     vss    0.024f
C41 sn     vss    0.041f
C42 a0     vss    0.024f
C43 s      vss    0.070f
.ends
