magic
tech scmos
timestamp 1170759828
<< checkpaint >>
rect -22 -26 86 114
<< ab >>
rect 0 0 64 88
<< pwell >>
rect -4 -8 68 40
<< nwell >>
rect -4 40 68 96
<< polysilicon >>
rect 2 82 11 83
rect 2 78 6 82
rect 10 78 11 82
rect 2 77 11 78
rect 9 74 11 77
rect 21 77 30 83
rect 34 77 43 83
rect 21 74 23 77
rect 41 74 43 77
rect 53 77 62 83
rect 53 74 55 77
rect 9 43 11 46
rect 21 43 23 46
rect 41 43 43 46
rect 53 43 55 46
rect 2 37 14 43
rect 18 42 30 43
rect 18 38 22 42
rect 26 38 30 42
rect 18 37 30 38
rect 34 42 46 43
rect 34 38 38 42
rect 42 38 46 42
rect 34 37 46 38
rect 50 42 62 43
rect 50 38 54 42
rect 58 38 62 42
rect 50 37 62 38
rect 9 34 11 37
rect 21 34 23 37
rect 41 34 43 37
rect 53 34 55 37
rect 9 11 11 14
rect 2 5 11 11
rect 21 11 23 14
rect 41 11 43 14
rect 21 5 30 11
rect 34 5 43 11
rect 53 11 55 14
rect 53 5 62 11
<< ndiffusion >>
rect 2 14 9 34
rect 11 26 21 34
rect 11 22 14 26
rect 18 22 21 26
rect 11 19 21 22
rect 11 15 14 19
rect 18 15 21 19
rect 11 14 21 15
rect 23 26 30 34
rect 23 22 25 26
rect 29 22 30 26
rect 23 19 30 22
rect 23 15 25 19
rect 29 15 30 19
rect 23 14 30 15
rect 34 19 41 34
rect 34 15 35 19
rect 39 15 41 19
rect 34 14 41 15
rect 43 26 53 34
rect 43 22 46 26
rect 50 22 53 26
rect 43 19 53 22
rect 43 15 46 19
rect 50 15 53 19
rect 43 14 53 15
rect 55 32 62 34
rect 55 28 57 32
rect 61 28 62 32
rect 55 25 62 28
rect 55 21 57 25
rect 61 21 62 25
rect 55 14 62 21
rect 13 2 19 14
rect 45 2 51 14
<< pdiffusion >>
rect 13 74 19 86
rect 45 74 51 86
rect 2 46 9 74
rect 11 73 21 74
rect 11 69 14 73
rect 18 69 21 73
rect 11 66 21 69
rect 11 62 14 66
rect 18 62 21 66
rect 11 46 21 62
rect 23 73 30 74
rect 23 69 25 73
rect 29 69 30 73
rect 23 65 30 69
rect 23 61 25 65
rect 29 61 30 65
rect 23 46 30 61
rect 34 73 41 74
rect 34 69 35 73
rect 39 69 41 73
rect 34 65 41 69
rect 34 61 35 65
rect 39 61 41 65
rect 34 46 41 61
rect 43 58 53 74
rect 43 54 46 58
rect 50 54 53 58
rect 43 51 53 54
rect 43 47 46 51
rect 50 47 53 51
rect 43 46 53 47
rect 55 73 62 74
rect 55 69 57 73
rect 61 69 62 73
rect 55 46 62 69
<< metal1 >>
rect -2 86 2 90
rect 10 86 22 90
rect 30 86 34 90
rect 42 86 54 90
rect 62 86 66 90
rect 6 82 10 86
rect 6 77 10 78
rect 14 82 18 86
rect 14 73 18 78
rect 57 82 61 86
rect 57 73 61 78
rect 24 69 25 73
rect 29 69 35 73
rect 39 69 40 73
rect 14 66 18 69
rect 57 68 61 69
rect 14 61 18 62
rect 24 61 25 65
rect 29 61 35 65
rect 39 61 40 65
rect 46 58 50 63
rect 22 42 26 55
rect 22 33 26 38
rect 38 42 42 55
rect 38 33 42 38
rect 46 51 50 54
rect 46 33 50 47
rect 54 42 58 63
rect 54 37 58 38
rect 46 32 61 33
rect 46 29 57 32
rect 54 28 57 29
rect 14 26 18 27
rect 14 19 18 22
rect 24 22 25 26
rect 29 22 46 26
rect 50 22 51 26
rect 24 19 30 22
rect 45 19 51 22
rect 24 15 25 19
rect 29 15 30 19
rect 34 15 35 19
rect 39 15 40 19
rect 45 15 46 19
rect 50 15 51 19
rect 54 25 61 28
rect 54 21 57 25
rect 54 17 61 21
rect 14 10 18 15
rect 14 2 18 6
rect 34 10 40 15
rect 34 6 35 10
rect 39 6 40 10
rect 34 2 40 6
rect -2 -2 2 2
rect 10 -2 22 2
rect 30 -2 34 2
rect 42 -2 54 2
rect 62 -2 66 2
<< metal2 >>
rect -2 86 6 90
rect 10 86 22 90
rect 26 86 38 90
rect 42 86 54 90
rect 58 86 66 90
rect -2 82 66 86
rect -2 78 14 82
rect 18 78 57 82
rect 61 78 66 82
rect -2 76 66 78
rect -2 10 66 12
rect -2 6 14 10
rect 18 6 35 10
rect 39 6 66 10
rect -2 2 66 6
rect -2 -2 6 2
rect 10 -2 22 2
rect 26 -2 38 2
rect 42 -2 54 2
rect 58 -2 66 2
<< ntransistor >>
rect 9 14 11 34
rect 21 14 23 34
rect 41 14 43 34
rect 53 14 55 34
<< ptransistor >>
rect 9 46 11 74
rect 21 46 23 74
rect 41 46 43 74
rect 53 46 55 74
<< polycontact >>
rect 6 78 10 82
rect 22 38 26 42
rect 38 38 42 42
rect 54 38 58 42
<< ndcontact >>
rect 14 22 18 26
rect 14 15 18 19
rect 25 22 29 26
rect 25 15 29 19
rect 35 15 39 19
rect 46 22 50 26
rect 46 15 50 19
rect 57 28 61 32
rect 57 21 61 25
<< pdcontact >>
rect 14 69 18 73
rect 14 62 18 66
rect 25 69 29 73
rect 25 61 29 65
rect 35 69 39 73
rect 35 61 39 65
rect 46 54 50 58
rect 46 47 50 51
rect 57 69 61 73
<< m2contact >>
rect 6 86 10 90
rect 22 86 26 90
rect 38 86 42 90
rect 54 86 58 90
rect 14 78 18 82
rect 57 78 61 82
rect 14 6 18 10
rect 35 6 39 10
rect 6 -2 10 2
rect 22 -2 26 2
rect 38 -2 42 2
rect 54 -2 58 2
<< psubstratepcontact >>
rect 2 -2 6 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 58 -2 62 2
<< nsubstratencontact >>
rect 2 86 6 90
rect 26 86 30 90
rect 34 86 38 90
rect 58 86 62 90
<< psubstratepdiff >>
rect 0 2 7 3
rect 25 2 39 3
rect 57 2 64 3
rect 0 -2 2 2
rect 6 -2 7 2
rect 0 -3 7 -2
rect 25 -2 26 2
rect 30 -2 34 2
rect 38 -2 39 2
rect 25 -3 39 -2
rect 57 -2 58 2
rect 62 -2 64 2
rect 57 -3 64 -2
<< nsubstratendiff >>
rect 0 90 7 91
rect 0 86 2 90
rect 6 86 7 90
rect 25 90 39 91
rect 25 86 26 90
rect 30 86 34 90
rect 38 86 39 90
rect 57 90 64 91
rect 57 86 58 90
rect 62 86 64 90
rect 0 85 7 86
rect 25 85 39 86
rect 57 85 64 86
<< labels >>
rlabel metal1 24 44 24 44 6 a1
rlabel metal1 40 44 40 44 6 a2
rlabel metal1 56 24 56 24 6 z
rlabel pdcontact 48 48 48 48 6 z
rlabel metal1 56 52 56 52 6 b
rlabel metal2 32 6 32 6 6 vss
rlabel metal2 32 82 32 82 6 vdd
<< end >>
