.subckt vddtie vdd vss z
*   SPICE3 file   created from vddtie.ext -      technology: scmos
m00 z      vss    vdd    vdd p w=30u  l=2.3636u ad=270p     pd=78u      as=270p     ps=78u
m01 z      vss    vss    vss n w=23u  l=2.3636u ad=207p     pd=64u      as=207p     ps=64u
C0  z      vss    0.171f
C1  vss    vdd    0.008f
C2  z      vdd    0.113f
C3  z      vss    0.008f
.ends
