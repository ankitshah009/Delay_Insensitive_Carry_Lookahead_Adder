.subckt bf1v0x1 a vdd vss z
*   SPICE3 file   created from bf1v0x1.ext -      technology: scmos
m00 vdd    an     z      vdd p w=18u  l=2.3636u ad=144p     pd=47.6129u as=116p     ps=50u
m01 an     a      vdd    vdd p w=13u  l=2.3636u ad=77p      pd=40u      as=104p     ps=34.3871u
m02 vss    an     z      vss n w=9u   l=2.3636u ad=46.5882p pd=20.1176u as=57p      ps=32u
m03 an     a      vss    vss n w=8u   l=2.3636u ad=52p      pd=30u      as=41.4118p ps=17.8824u
C0  vss    a      0.003f
C1  vss    an     0.062f
C2  a      z      0.046f
C3  z      an     0.080f
C4  a      vdd    0.083f
C5  an     vdd    0.022f
C6  vss    z      0.035f
C7  a      an     0.079f
C8  vss    vdd    0.003f
C9  z      vdd    0.039f
C11 a      vss    0.021f
C12 z      vss    0.006f
C13 an     vss    0.026f
.ends
