magic
tech scmos
timestamp 1179385516
<< checkpaint >>
rect -22 -22 54 94
<< ab >>
rect 0 0 32 72
<< pwell >>
rect -4 -4 36 32
<< nwell >>
rect -4 32 36 76
<< polysilicon >>
rect 9 56 11 61
rect 21 60 27 61
rect 21 56 22 60
rect 26 56 27 60
rect 21 55 27 56
rect 21 52 23 55
rect 9 35 11 38
rect 9 34 16 35
rect 9 30 11 34
rect 15 30 16 34
rect 9 29 16 30
rect 9 26 11 29
rect 21 26 23 38
rect 9 12 11 17
rect 21 14 23 19
<< ndiffusion >>
rect 2 25 9 26
rect 2 21 3 25
rect 7 21 9 25
rect 2 20 9 21
rect 4 17 9 20
rect 11 23 21 26
rect 11 19 14 23
rect 18 19 21 23
rect 23 25 30 26
rect 23 21 25 25
rect 29 21 30 25
rect 23 19 30 21
rect 11 17 19 19
<< pdiffusion >>
rect 13 68 19 69
rect 13 64 14 68
rect 18 64 19 68
rect 13 56 19 64
rect 4 51 9 56
rect 2 50 9 51
rect 2 46 3 50
rect 7 46 9 50
rect 2 43 9 46
rect 2 39 3 43
rect 7 39 9 43
rect 2 38 9 39
rect 11 52 19 56
rect 11 38 21 52
rect 23 44 28 52
rect 23 43 30 44
rect 23 39 25 43
rect 29 39 30 43
rect 23 38 30 39
<< metal1 >>
rect -2 68 34 72
rect -2 64 4 68
rect 8 64 14 68
rect 18 64 24 68
rect 28 64 34 68
rect 21 59 22 60
rect 18 56 22 59
rect 26 59 27 60
rect 26 56 30 59
rect 18 53 30 56
rect 2 50 14 51
rect 2 46 3 50
rect 7 46 14 50
rect 2 45 14 46
rect 18 45 22 53
rect 2 43 7 45
rect 2 39 3 43
rect 2 38 7 39
rect 25 43 29 44
rect 2 25 6 38
rect 25 34 29 39
rect 10 30 11 34
rect 15 30 30 34
rect 24 25 30 30
rect 2 21 3 25
rect 7 21 8 25
rect 14 23 18 24
rect 24 21 25 25
rect 29 21 30 25
rect 14 8 18 19
rect -2 4 4 8
rect 8 4 24 8
rect 28 4 34 8
rect -2 0 34 4
<< ntransistor >>
rect 9 17 11 26
rect 21 19 23 26
<< ptransistor >>
rect 9 38 11 56
rect 21 38 23 52
<< polycontact >>
rect 22 56 26 60
rect 11 30 15 34
<< ndcontact >>
rect 3 21 7 25
rect 14 19 18 23
rect 25 21 29 25
<< pdcontact >>
rect 14 64 18 68
rect 3 46 7 50
rect 3 39 7 43
rect 25 39 29 43
<< psubstratepcontact >>
rect 4 4 8 8
rect 24 4 28 8
<< nsubstratencontact >>
rect 4 64 8 68
rect 24 64 28 68
<< psubstratepdiff >>
rect 3 8 29 9
rect 3 4 4 8
rect 8 4 24 8
rect 28 4 29 8
rect 3 3 29 4
<< nsubstratendiff >>
rect 3 68 9 69
rect 3 64 4 68
rect 8 64 9 68
rect 3 63 9 64
rect 23 68 29 69
rect 23 64 24 68
rect 28 64 29 68
rect 23 63 29 64
<< labels >>
rlabel polycontact 12 32 12 32 6 an
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 48 12 48 6 z
rlabel metal1 16 4 16 4 6 vss
rlabel metal1 20 52 20 52 6 a
rlabel metal1 16 68 16 68 6 vdd
rlabel metal1 20 32 20 32 6 an
rlabel metal1 27 32 27 32 6 an
rlabel metal1 28 56 28 56 6 a
<< end >>
