magic
tech scmos
timestamp 1179385843
<< checkpaint >>
rect -22 -22 62 94
<< ab >>
rect 0 0 40 72
<< pwell >>
rect -4 -4 44 32
<< nwell >>
rect -4 32 44 76
<< polysilicon >>
rect 9 65 11 70
rect 19 65 21 70
rect 29 65 31 70
rect 9 35 11 38
rect 19 35 21 38
rect 29 35 31 38
rect 9 34 31 35
rect 9 30 18 34
rect 22 30 26 34
rect 30 30 31 34
rect 9 29 31 30
rect 9 26 11 29
rect 19 26 21 29
rect 9 2 11 6
rect 19 2 21 6
<< ndiffusion >>
rect 2 18 9 26
rect 2 14 3 18
rect 7 14 9 18
rect 2 11 9 14
rect 2 7 3 11
rect 7 7 9 11
rect 2 6 9 7
rect 11 25 19 26
rect 11 21 13 25
rect 17 21 19 25
rect 11 18 19 21
rect 11 14 13 18
rect 17 14 19 18
rect 11 6 19 14
rect 21 25 29 26
rect 21 21 23 25
rect 27 21 29 25
rect 21 18 29 21
rect 21 14 23 18
rect 27 14 29 18
rect 21 13 29 14
rect 21 6 27 13
<< pdiffusion >>
rect 4 51 9 65
rect 2 50 9 51
rect 2 46 3 50
rect 7 46 9 50
rect 2 43 9 46
rect 2 39 3 43
rect 7 39 9 43
rect 2 38 9 39
rect 11 64 19 65
rect 11 60 13 64
rect 17 60 19 64
rect 11 56 19 60
rect 11 52 13 56
rect 17 52 19 56
rect 11 38 19 52
rect 21 50 29 65
rect 21 46 23 50
rect 27 46 29 50
rect 21 43 29 46
rect 21 39 23 43
rect 27 39 29 43
rect 21 38 29 39
rect 31 64 38 65
rect 31 60 33 64
rect 37 60 38 64
rect 31 56 38 60
rect 31 52 33 56
rect 37 52 38 56
rect 31 38 38 52
<< metal1 >>
rect -2 64 42 72
rect 13 56 17 60
rect 13 51 17 52
rect 33 56 37 60
rect 33 51 37 52
rect 2 50 7 51
rect 2 46 3 50
rect 2 43 7 46
rect 2 39 3 43
rect 23 50 27 51
rect 23 43 27 46
rect 7 39 23 42
rect 2 38 27 39
rect 2 26 6 38
rect 34 34 38 43
rect 17 30 18 34
rect 22 30 26 34
rect 30 30 38 34
rect 2 25 17 26
rect 2 22 13 25
rect 13 18 17 21
rect 2 14 3 18
rect 7 14 8 18
rect 2 11 8 14
rect 13 13 17 14
rect 22 21 23 25
rect 27 21 28 25
rect 34 21 38 30
rect 22 18 28 21
rect 22 14 23 18
rect 27 14 28 18
rect 2 8 3 11
rect -2 7 3 8
rect 7 8 8 11
rect 22 8 28 14
rect 7 7 32 8
rect -2 4 32 7
rect 36 4 42 8
rect -2 0 42 4
<< ntransistor >>
rect 9 6 11 26
rect 19 6 21 26
<< ptransistor >>
rect 9 38 11 65
rect 19 38 21 65
rect 29 38 31 65
<< polycontact >>
rect 18 30 22 34
rect 26 30 30 34
<< ndcontact >>
rect 3 14 7 18
rect 3 7 7 11
rect 13 21 17 25
rect 13 14 17 18
rect 23 21 27 25
rect 23 14 27 18
<< pdcontact >>
rect 3 46 7 50
rect 3 39 7 43
rect 13 60 17 64
rect 13 52 17 56
rect 23 46 27 50
rect 23 39 27 43
rect 33 60 37 64
rect 33 52 37 56
<< psubstratepcontact >>
rect 32 4 36 8
<< psubstratepdiff >>
rect 31 8 37 9
rect 31 4 32 8
rect 36 4 37 8
rect 31 3 37 4
<< labels >>
rlabel pdcontact 4 40 4 40 6 z
rlabel metal1 12 24 12 24 6 z
rlabel metal1 12 40 12 40 6 z
rlabel metal1 20 4 20 4 6 vss
rlabel polycontact 20 32 20 32 6 a
rlabel metal1 20 40 20 40 6 z
rlabel metal1 20 68 20 68 6 vdd
rlabel metal1 36 32 36 32 6 a
<< end >>
