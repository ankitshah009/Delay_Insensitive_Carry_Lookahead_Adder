.subckt cgi2cv0x1 a b c vdd vss z
*   SPICE3 file   created from cgi2cv0x1.ext -      technology: scmos
m00 vdd    a      n1     vdd p w=27u  l=2.3636u ad=121.5p   pd=36u      as=125.667p ps=46u
m01 w1     a      vdd    vdd p w=27u  l=2.3636u ad=67.5p    pd=32u      as=121.5p   ps=36u
m02 z      b      w1     vdd p w=27u  l=2.3636u ad=108p     pd=35u      as=67.5p    ps=32u
m03 n1     w2     z      vdd p w=27u  l=2.3636u ad=125.667p pd=46u      as=108p     ps=35u
m04 vdd    b      n1     vdd p w=27u  l=2.3636u ad=121.5p   pd=36u      as=125.667p ps=46u
m05 w2     c      vdd    vdd p w=27u  l=2.3636u ad=161p     pd=68u      as=121.5p   ps=36u
m06 vss    a      n3     vss n w=12u  l=2.3636u ad=73.5p    pd=27u      as=56p      ps=26u
m07 w3     a      vss    vss n w=12u  l=2.3636u ad=30p      pd=17u      as=73.5p    ps=27u
m08 z      b      w3     vss n w=12u  l=2.3636u ad=48p      pd=20u      as=30p      ps=17u
m09 n3     w2     z      vss n w=12u  l=2.3636u ad=56p      pd=26u      as=48p      ps=20u
m10 vss    b      n3     vss n w=12u  l=2.3636u ad=73.5p    pd=27u      as=56p      ps=26u
m11 w2     c      vss    vss n w=12u  l=2.3636u ad=72p      pd=38u      as=73.5p    ps=27u
C0  n1     b      0.081f
C1  vdd    a      0.022f
C2  c      w2     0.291f
C3  n3     vdd    0.005f
C4  c      a      0.010f
C5  w2     b      0.322f
C6  z      vdd    0.062f
C7  vss    n1     0.018f
C8  b      a      0.126f
C9  n3     b      0.014f
C10 vss    w2     0.131f
C11 w1     n1     0.023f
C12 z      c      0.033f
C13 w3     n3     0.006f
C14 vdd    c      0.068f
C15 z      b      0.120f
C16 vss    a      0.020f
C17 n3     vss    0.337f
C18 w3     z      0.008f
C19 vdd    b      0.032f
C20 n1     w2     0.024f
C21 vss    z      0.068f
C22 n1     a      0.042f
C23 c      b      0.252f
C24 vss    vdd    0.002f
C25 n3     n1     0.038f
C26 z      w1     0.007f
C27 w2     a      0.041f
C28 n3     w2     0.087f
C29 w1     vdd    0.004f
C30 z      n1     0.191f
C31 vss    c      0.014f
C32 vdd    n1     0.370f
C33 z      w2     0.068f
C34 vss    b      0.032f
C35 n3     a      0.041f
C36 n1     c      0.008f
C37 z      a      0.098f
C38 vdd    w2     0.044f
C39 n3     z      0.177f
C40 n3     vss    0.003f
C42 z      vss    0.003f
C44 c      vss    0.015f
C45 w2     vss    0.024f
C46 b      vss    0.040f
C47 a      vss    0.042f
.ends
