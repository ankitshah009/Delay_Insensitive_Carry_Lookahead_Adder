magic
tech scmos
timestamp 1179387646
<< checkpaint >>
rect -22 -25 134 105
<< ab >>
rect 0 0 112 80
<< pwell >>
rect -4 -7 116 36
<< nwell >>
rect -4 36 116 87
<< polysilicon >>
rect 9 70 11 74
rect 19 70 21 74
rect 61 70 63 74
rect 71 70 73 74
rect 29 63 31 68
rect 39 63 41 68
rect 48 47 54 48
rect 48 43 49 47
rect 53 43 54 47
rect 48 42 54 43
rect 81 63 83 68
rect 91 63 93 68
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 39 39 41 42
rect 48 39 50 42
rect 9 38 25 39
rect 9 37 20 38
rect 16 34 20 37
rect 24 34 25 38
rect 29 37 50 39
rect 61 39 63 42
rect 71 39 73 42
rect 81 39 83 42
rect 91 39 93 42
rect 61 38 73 39
rect 61 37 66 38
rect 16 33 25 34
rect 9 28 11 33
rect 16 31 28 33
rect 16 28 18 31
rect 26 28 28 31
rect 33 28 35 37
rect 65 34 66 37
rect 70 37 73 38
rect 78 38 103 39
rect 78 37 98 38
rect 70 34 71 37
rect 65 33 71 34
rect 78 33 80 37
rect 97 34 98 37
rect 102 34 103 38
rect 97 33 103 34
rect 65 28 67 33
rect 75 31 80 33
rect 75 28 77 31
rect 85 30 91 31
rect 9 8 11 16
rect 16 12 18 16
rect 26 12 28 16
rect 33 8 35 16
rect 9 6 35 8
rect 85 26 86 30
rect 90 27 91 30
rect 90 26 97 27
rect 85 25 97 26
rect 85 22 87 25
rect 95 22 97 25
rect 65 6 67 10
rect 75 6 77 10
rect 85 8 87 13
rect 95 8 97 13
<< ndiffusion >>
rect 2 21 9 28
rect 2 17 3 21
rect 7 17 9 21
rect 2 16 9 17
rect 11 16 16 28
rect 18 27 26 28
rect 18 23 20 27
rect 24 23 26 27
rect 18 16 26 23
rect 28 16 33 28
rect 35 16 44 28
rect 60 23 65 28
rect 58 22 65 23
rect 58 18 59 22
rect 63 18 65 22
rect 58 17 65 18
rect 37 12 44 16
rect 37 8 38 12
rect 42 8 44 12
rect 60 10 65 17
rect 67 27 75 28
rect 67 23 69 27
rect 73 23 75 27
rect 67 10 75 23
rect 77 22 83 28
rect 77 18 85 22
rect 77 14 79 18
rect 83 14 85 18
rect 77 13 85 14
rect 87 21 95 22
rect 87 17 89 21
rect 93 17 95 21
rect 87 13 95 17
rect 97 13 105 22
rect 77 10 83 13
rect 37 7 44 8
rect 99 12 105 13
rect 99 8 100 12
rect 104 8 105 12
rect 99 7 105 8
<< pdiffusion >>
rect 4 63 9 70
rect 2 62 9 63
rect 2 58 3 62
rect 7 58 9 62
rect 2 55 9 58
rect 2 51 3 55
rect 7 51 9 55
rect 2 50 9 51
rect 4 42 9 50
rect 11 54 19 70
rect 11 50 13 54
rect 17 50 19 54
rect 11 47 19 50
rect 11 43 13 47
rect 17 43 19 47
rect 11 42 19 43
rect 21 63 26 70
rect 54 69 61 70
rect 54 65 55 69
rect 59 65 61 69
rect 21 62 29 63
rect 21 58 23 62
rect 27 58 29 62
rect 21 42 29 58
rect 31 47 39 63
rect 31 43 33 47
rect 37 43 39 47
rect 31 42 39 43
rect 41 62 48 63
rect 41 58 43 62
rect 47 58 48 62
rect 41 57 48 58
rect 54 62 61 65
rect 54 58 55 62
rect 59 58 61 62
rect 54 57 61 58
rect 41 42 46 57
rect 56 42 61 57
rect 63 61 71 70
rect 63 57 65 61
rect 69 57 71 61
rect 63 54 71 57
rect 63 50 65 54
rect 69 50 71 54
rect 63 42 71 50
rect 73 63 79 70
rect 73 62 81 63
rect 73 58 75 62
rect 79 58 81 62
rect 73 42 81 58
rect 83 47 91 63
rect 83 43 85 47
rect 89 43 91 47
rect 83 42 91 43
rect 93 62 100 63
rect 93 58 95 62
rect 99 58 100 62
rect 93 42 100 58
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect -2 69 114 78
rect -2 68 55 69
rect 54 65 55 68
rect 59 68 114 69
rect 59 65 60 68
rect 54 62 60 65
rect 74 62 80 68
rect 2 58 3 62
rect 7 58 23 62
rect 27 58 43 62
rect 47 58 48 62
rect 54 58 55 62
rect 59 58 60 62
rect 65 61 69 62
rect 2 55 7 58
rect 2 51 3 55
rect 74 58 75 62
rect 79 58 80 62
rect 94 62 100 68
rect 94 58 95 62
rect 99 58 100 62
rect 65 54 69 57
rect 2 50 7 51
rect 12 50 13 54
rect 17 50 65 54
rect 69 50 110 54
rect 2 30 6 50
rect 12 47 17 50
rect 49 47 53 50
rect 12 43 13 47
rect 12 42 17 43
rect 32 43 33 47
rect 37 43 38 47
rect 32 38 38 43
rect 84 46 85 47
rect 49 42 53 43
rect 57 43 85 46
rect 89 43 90 47
rect 57 42 90 43
rect 57 38 61 42
rect 97 38 103 46
rect 19 34 20 38
rect 24 34 61 38
rect 65 34 66 38
rect 70 34 82 38
rect 89 34 98 38
rect 102 34 103 38
rect 57 30 61 34
rect 78 30 82 34
rect 2 27 24 30
rect 2 26 20 27
rect 57 27 73 30
rect 57 26 69 27
rect 20 22 24 23
rect 78 26 86 30
rect 90 26 91 30
rect 69 22 73 23
rect 3 21 7 22
rect 20 18 59 22
rect 63 18 64 22
rect 106 21 110 50
rect 79 18 83 19
rect 3 12 7 17
rect 88 17 89 21
rect 93 17 110 21
rect 79 12 83 14
rect -2 8 38 12
rect 42 8 100 12
rect 104 8 114 12
rect -2 2 114 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
<< ntransistor >>
rect 9 16 11 28
rect 16 16 18 28
rect 26 16 28 28
rect 33 16 35 28
rect 65 10 67 28
rect 75 10 77 28
rect 85 13 87 22
rect 95 13 97 22
<< ptransistor >>
rect 9 42 11 70
rect 19 42 21 70
rect 29 42 31 63
rect 39 42 41 63
rect 61 42 63 70
rect 71 42 73 70
rect 81 42 83 63
rect 91 42 93 63
<< polycontact >>
rect 49 43 53 47
rect 20 34 24 38
rect 66 34 70 38
rect 98 34 102 38
rect 86 26 90 30
<< ndcontact >>
rect 3 17 7 21
rect 20 23 24 27
rect 59 18 63 22
rect 38 8 42 12
rect 69 23 73 27
rect 79 14 83 18
rect 89 17 93 21
rect 100 8 104 12
<< pdcontact >>
rect 3 58 7 62
rect 3 51 7 55
rect 13 50 17 54
rect 13 43 17 47
rect 55 65 59 69
rect 23 58 27 62
rect 33 43 37 47
rect 43 58 47 62
rect 55 58 59 62
rect 65 57 69 61
rect 65 50 69 54
rect 75 58 79 62
rect 85 43 89 47
rect 95 58 99 62
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
rect 90 -2 94 2
rect 98 -2 102 2
rect 106 -2 110 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
rect 90 78 94 82
rect 98 78 102 82
rect 106 78 110 82
<< psubstratepdiff >>
rect 0 2 112 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 112 2
rect 0 -3 112 -2
<< nsubstratendiff >>
rect 0 82 112 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 112 82
rect 0 77 112 78
<< labels >>
rlabel polycontact 51 45 51 45 6 bn
rlabel metal1 12 28 12 28 6 z
rlabel metal1 4 44 4 44 6 z
rlabel metal1 14 48 14 48 6 bn
rlabel metal1 12 60 12 60 6 z
rlabel metal1 20 28 20 28 6 z
rlabel metal1 36 20 36 20 6 z
rlabel metal1 28 20 28 20 6 z
rlabel metal1 35 40 35 40 6 an
rlabel metal1 20 60 20 60 6 z
rlabel metal1 36 60 36 60 6 z
rlabel metal1 28 60 28 60 6 z
rlabel metal1 56 6 56 6 6 vss
rlabel metal1 44 20 44 20 6 z
rlabel ndcontact 60 20 60 20 6 z
rlabel metal1 52 20 52 20 6 z
rlabel metal1 40 36 40 36 6 an
rlabel metal1 51 48 51 48 6 bn
rlabel pdcontact 44 60 44 60 6 z
rlabel metal1 56 74 56 74 6 vdd
rlabel ndcontact 71 26 71 26 6 an
rlabel metal1 84 28 84 28 6 b
rlabel polycontact 68 36 68 36 6 b
rlabel metal1 73 44 73 44 6 an
rlabel metal1 76 36 76 36 6 b
rlabel metal1 67 56 67 56 6 bn
rlabel metal1 99 19 99 19 6 bn
rlabel metal1 92 36 92 36 6 a
rlabel metal1 100 40 100 40 6 a
rlabel metal1 61 52 61 52 6 bn
<< end >>
