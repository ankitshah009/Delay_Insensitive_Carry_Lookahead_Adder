magic
tech scmos
timestamp 1179385184
<< checkpaint >>
rect -22 -25 70 105
<< ab >>
rect 0 0 48 80
<< pwell >>
rect -4 -7 52 36
<< nwell >>
rect -4 36 52 87
<< polysilicon >>
rect 10 70 12 74
rect 17 70 19 74
rect 27 70 29 74
rect 37 70 39 74
rect 10 39 12 42
rect 2 38 12 39
rect 2 34 3 38
rect 7 34 12 38
rect 2 33 12 34
rect 17 39 19 42
rect 27 39 29 42
rect 37 39 39 42
rect 17 38 23 39
rect 17 34 18 38
rect 22 34 23 38
rect 17 33 23 34
rect 27 38 33 39
rect 27 34 28 38
rect 32 34 33 38
rect 27 33 33 34
rect 37 38 46 39
rect 37 34 41 38
rect 45 34 46 38
rect 37 33 46 34
rect 10 30 12 33
rect 20 30 22 33
rect 10 19 12 24
rect 20 20 22 24
rect 30 23 32 33
rect 37 23 39 33
rect 30 9 32 14
rect 37 9 39 14
<< ndiffusion >>
rect 2 24 10 30
rect 12 29 20 30
rect 12 25 14 29
rect 18 25 20 29
rect 12 24 20 25
rect 22 24 28 30
rect 2 15 8 24
rect 24 23 28 24
rect 24 18 30 23
rect 2 11 3 15
rect 7 11 8 15
rect 2 10 8 11
rect 22 15 30 18
rect 22 11 23 15
rect 27 14 30 15
rect 32 14 37 23
rect 39 22 46 23
rect 39 18 41 22
rect 45 18 46 22
rect 39 17 46 18
rect 39 14 44 17
rect 27 11 28 14
rect 22 10 28 11
<< pdiffusion >>
rect 5 55 10 70
rect 3 54 10 55
rect 3 50 4 54
rect 8 50 10 54
rect 3 47 10 50
rect 3 43 4 47
rect 8 43 10 47
rect 3 42 10 43
rect 12 42 17 70
rect 19 62 27 70
rect 19 58 21 62
rect 25 58 27 62
rect 19 42 27 58
rect 29 69 37 70
rect 29 65 31 69
rect 35 65 37 69
rect 29 42 37 65
rect 39 63 44 70
rect 39 62 46 63
rect 39 58 41 62
rect 45 58 46 62
rect 39 57 46 58
rect 39 42 44 57
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect -2 69 50 78
rect -2 68 31 69
rect 30 65 31 68
rect 35 68 50 69
rect 35 65 36 68
rect 2 55 6 63
rect 20 58 21 62
rect 25 58 41 62
rect 45 58 46 62
rect 2 54 8 55
rect 2 50 4 54
rect 2 47 8 50
rect 18 49 30 55
rect 34 49 46 55
rect 2 43 4 47
rect 8 43 14 47
rect 2 38 7 39
rect 2 34 3 38
rect 2 33 7 34
rect 2 22 6 33
rect 10 30 14 43
rect 18 38 22 49
rect 18 33 22 34
rect 26 38 34 39
rect 26 34 28 38
rect 32 34 34 38
rect 40 38 46 49
rect 40 34 41 38
rect 45 34 46 38
rect 26 33 34 34
rect 30 30 34 33
rect 10 29 24 30
rect 10 25 14 29
rect 18 25 24 29
rect 30 26 39 30
rect 20 22 24 25
rect 2 18 15 22
rect 20 18 41 22
rect 45 18 46 22
rect 2 12 3 15
rect -2 11 3 12
rect 7 12 8 15
rect 22 12 23 15
rect 7 11 23 12
rect 27 12 28 15
rect 27 11 50 12
rect -2 2 50 11
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
<< ntransistor >>
rect 10 24 12 30
rect 20 24 22 30
rect 30 14 32 23
rect 37 14 39 23
<< ptransistor >>
rect 10 42 12 70
rect 17 42 19 70
rect 27 42 29 70
rect 37 42 39 70
<< polycontact >>
rect 3 34 7 38
rect 18 34 22 38
rect 28 34 32 38
rect 41 34 45 38
<< ndcontact >>
rect 14 25 18 29
rect 3 11 7 15
rect 23 11 27 15
rect 41 18 45 22
<< pdcontact >>
rect 4 50 8 54
rect 4 43 8 47
rect 21 58 25 62
rect 31 65 35 69
rect 41 58 45 62
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
<< psubstratepdiff >>
rect 0 2 48 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 48 2
rect 0 -3 48 -2
<< nsubstratendiff >>
rect 0 82 48 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 48 82
rect 0 77 48 78
<< labels >>
rlabel metal1 4 32 4 32 6 c
rlabel metal1 4 56 4 56 6 z
rlabel metal1 12 20 12 20 6 c
rlabel metal1 12 36 12 36 6 z
rlabel metal1 24 6 24 6 6 vss
rlabel metal1 20 44 20 44 6 b
rlabel metal1 24 74 24 74 6 vdd
rlabel metal1 28 20 28 20 6 z
rlabel metal1 36 28 36 28 6 a1
rlabel metal1 36 20 36 20 6 z
rlabel metal1 28 36 28 36 6 a1
rlabel metal1 36 52 36 52 6 a2
rlabel metal1 28 52 28 52 6 b
rlabel metal1 44 48 44 48 6 a2
rlabel metal1 33 60 33 60 6 n1
<< end >>
