.subckt xor3v1x05 a b c vdd vss z
*   SPICE3 file   created from xor3v1x05.ext -      technology: scmos
m00 vdd    b      bn     vdd p w=19u  l=2.3636u ad=117.8p   pd=37.4571u as=107p     ps=52u
m01 an     a      vdd    vdd p w=19u  l=2.3636u ad=76p      pd=27u      as=117.8p   ps=37.4571u
m02 iz     bn     an     vdd p w=19u  l=2.3636u ad=76p      pd=27u      as=76p      ps=27u
m03 bn     an     iz     vdd p w=19u  l=2.3636u ad=107p     pd=52u      as=76p      ps=27u
m04 vdd    c      cn     vdd p w=16u  l=2.3636u ad=99.2p    pd=31.5429u as=93p      ps=46u
m05 zn     iz     vdd    vdd p w=16u  l=2.3636u ad=64p      pd=24u      as=99.2p    ps=31.5429u
m06 z      cn     zn     vdd p w=16u  l=2.3636u ad=64p      pd=24u      as=64p      ps=24u
m07 cn     zn     z      vdd p w=16u  l=2.3636u ad=93p      pd=46u      as=64p      ps=24u
m08 vss    b      bn     vss n w=9u   l=2.3636u ad=77.0625p pd=33.375u  as=57p      ps=32u
m09 an     a      vss    vss n w=9u   l=2.3636u ad=36p      pd=17u      as=77.0625p ps=33.375u
m10 iz     b      an     vss n w=9u   l=2.3636u ad=36p      pd=17u      as=36p      ps=17u
m11 w1     bn     iz     vss n w=9u   l=2.3636u ad=22.5p    pd=14u      as=36p      ps=17u
m12 vss    an     w1     vss n w=9u   l=2.3636u ad=77.0625p pd=33.375u  as=22.5p    ps=14u
m13 vss    c      cn     vss n w=7u   l=2.3636u ad=59.9375p pd=25.9583u as=49p      ps=28u
m14 zn     iz     vss    vss n w=7u   l=2.3636u ad=28p      pd=15u      as=59.9375p ps=25.9583u
m15 z      c      zn     vss n w=7u   l=2.3636u ad=28p      pd=15u      as=28p      ps=15u
m16 w2     cn     z      vss n w=7u   l=2.3636u ad=17.5p    pd=12u      as=28p      ps=15u
m17 vss    zn     w2     vss n w=7u   l=2.3636u ad=59.9375p pd=25.9583u as=17.5p    ps=12u
C0  vss    cn     0.138f
C1  z      zn     0.405f
C2  w1     iz     0.010f
C3  iz     vdd    0.041f
C4  an     a      0.077f
C5  c      b      0.006f
C6  zn     cn     0.570f
C7  z      iz     0.003f
C8  vss    c      0.031f
C9  bn     b      0.187f
C10 an     vdd    0.046f
C11 vss    bn     0.075f
C12 cn     iz     0.156f
C13 zn     c      0.054f
C14 a      vdd    0.014f
C15 iz     c      0.242f
C16 vss    b      0.019f
C17 cn     an     0.025f
C18 iz     bn     0.252f
C19 z      vdd    0.037f
C20 c      an     0.061f
C21 vss    zn     0.082f
C22 cn     vdd    0.368f
C23 an     bn     0.586f
C24 c      a      0.004f
C25 iz     b      0.003f
C26 vss    iz     0.197f
C27 z      cn     0.231f
C28 an     b      0.046f
C29 bn     a      0.245f
C30 c      vdd    0.025f
C31 zn     iz     0.052f
C32 z      c      0.007f
C33 vss    an     0.132f
C34 a      b      0.121f
C35 bn     vdd    0.248f
C36 cn     c      0.236f
C37 vss    a      0.066f
C38 zn     an     0.006f
C39 b      vdd    0.082f
C40 w2     z      0.010f
C41 cn     bn     0.012f
C42 iz     an     0.487f
C43 vss    z      0.146f
C44 c      bn     0.031f
C45 zn     vdd    0.048f
C46 iz     a      0.017f
C48 z      vss    0.014f
C49 zn     vss    0.041f
C50 cn     vss    0.038f
C51 iz     vss    0.045f
C52 c      vss    0.053f
C53 an     vss    0.037f
C54 bn     vss    0.040f
C55 a      vss    0.029f
C56 b      vss    0.052f
.ends
