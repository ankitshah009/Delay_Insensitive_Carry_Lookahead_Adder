.subckt iv1v1x8 a vdd vss z
*   SPICE3 file   created from iv1v1x8.ext -      technology: scmos
m00 z      a      vdd    vdd p w=28u  l=2.3636u ad=114.154p pd=38.7692u as=150.769p ps=52.7692u
m01 vdd    a      z      vdd p w=28u  l=2.3636u ad=150.769p pd=52.7692u as=114.154p ps=38.7692u
m02 z      a      vdd    vdd p w=28u  l=2.3636u ad=114.154p pd=38.7692u as=150.769p ps=52.7692u
m03 vdd    a      z      vdd p w=20u  l=2.3636u ad=107.692p pd=37.6923u as=81.5385p ps=27.6923u
m04 z      a      vss    vss n w=9u   l=2.3636u ad=37.4348p pd=14.6087u as=49.9565p ps=18.7826u
m05 vss    a      z      vss n w=20u  l=2.3636u ad=111.014p pd=41.7391u as=83.1884p ps=32.4638u
m06 z      a      vss    vss n w=20u  l=2.3636u ad=83.1884p pd=32.4638u as=111.014p ps=41.7391u
m07 vss    a      z      vss n w=20u  l=2.3636u ad=111.014p pd=41.7391u as=83.1884p ps=32.4638u
C0  vss    z      0.270f
C1  z      a      0.326f
C2  vss    vdd    0.014f
C3  a      vdd    0.082f
C4  vss    a      0.047f
C5  z      vdd    0.144f
C7  z      vss    0.004f
C8  a      vss    0.058f
.ends
