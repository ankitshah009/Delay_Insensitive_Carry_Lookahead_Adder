magic
tech scmos
timestamp 1179387421
<< checkpaint >>
rect -22 -25 174 105
<< ab >>
rect 0 0 152 80
<< pwell >>
rect -4 -7 156 36
<< nwell >>
rect -4 36 156 87
<< polysilicon >>
rect 9 70 11 74
rect 19 70 21 74
rect 51 70 53 74
rect 58 70 60 74
rect 68 70 70 74
rect 78 70 80 74
rect 88 70 90 74
rect 95 70 97 74
rect 111 70 113 74
rect 121 70 123 74
rect 131 70 133 74
rect 141 70 143 74
rect 35 46 41 47
rect 35 42 36 46
rect 40 42 41 46
rect 9 39 11 42
rect 19 39 21 42
rect 9 38 21 39
rect 9 34 16 38
rect 20 34 21 38
rect 35 39 41 42
rect 51 39 53 42
rect 35 37 53 39
rect 35 35 41 37
rect 9 33 21 34
rect 9 30 11 33
rect 19 30 21 33
rect 29 33 41 35
rect 29 30 31 33
rect 39 30 41 33
rect 58 30 60 42
rect 68 39 70 42
rect 78 39 80 42
rect 64 38 80 39
rect 64 34 65 38
rect 69 37 80 38
rect 88 39 90 42
rect 95 39 97 42
rect 111 39 113 42
rect 121 39 123 42
rect 131 39 133 42
rect 69 34 70 37
rect 88 36 91 39
rect 95 38 107 39
rect 95 37 102 38
rect 64 33 70 34
rect 54 29 60 30
rect 54 25 55 29
rect 59 26 60 29
rect 79 28 81 33
rect 89 30 91 36
rect 101 34 102 37
rect 106 34 107 38
rect 101 33 107 34
rect 111 38 117 39
rect 111 34 112 38
rect 116 34 117 38
rect 111 33 117 34
rect 121 38 133 39
rect 121 34 122 38
rect 126 34 133 38
rect 141 39 143 42
rect 141 38 150 39
rect 141 35 145 38
rect 121 33 133 34
rect 114 30 116 33
rect 121 30 123 33
rect 131 30 133 33
rect 138 34 145 35
rect 149 34 150 38
rect 138 33 150 34
rect 138 30 140 33
rect 59 25 70 26
rect 54 24 70 25
rect 9 11 11 16
rect 19 11 21 16
rect 29 11 31 16
rect 39 11 41 16
rect 68 8 70 24
rect 79 8 81 11
rect 89 8 91 11
rect 68 6 91 8
rect 114 7 116 12
rect 121 7 123 12
rect 131 7 133 12
rect 138 7 140 12
<< ndiffusion >>
rect 2 29 9 30
rect 2 25 3 29
rect 7 25 9 29
rect 2 22 9 25
rect 2 18 3 22
rect 7 18 9 22
rect 2 16 9 18
rect 11 21 19 30
rect 11 17 13 21
rect 17 17 19 21
rect 11 16 19 17
rect 21 29 29 30
rect 21 25 23 29
rect 27 25 29 29
rect 21 22 29 25
rect 21 18 23 22
rect 27 18 29 22
rect 21 16 29 18
rect 31 22 39 30
rect 31 18 33 22
rect 37 18 39 22
rect 31 16 39 18
rect 41 29 48 30
rect 41 25 43 29
rect 47 25 48 29
rect 41 24 48 25
rect 84 28 89 30
rect 41 16 46 24
rect 74 23 79 28
rect 72 22 79 23
rect 72 18 73 22
rect 77 18 79 22
rect 72 17 79 18
rect 74 11 79 17
rect 81 21 89 28
rect 81 17 83 21
rect 87 17 89 21
rect 81 11 89 17
rect 91 29 98 30
rect 91 25 93 29
rect 97 25 98 29
rect 91 24 98 25
rect 91 11 96 24
rect 105 12 114 30
rect 116 12 121 30
rect 123 21 131 30
rect 123 17 125 21
rect 129 17 131 21
rect 123 12 131 17
rect 133 12 138 30
rect 140 26 148 30
rect 140 22 142 26
rect 146 22 148 26
rect 140 18 148 22
rect 140 14 142 18
rect 146 14 148 18
rect 140 12 148 14
rect 105 8 107 12
rect 111 8 112 12
rect 105 7 112 8
<< pdiffusion >>
rect 99 70 109 72
rect 2 69 9 70
rect 2 65 3 69
rect 7 65 9 69
rect 2 61 9 65
rect 2 57 3 61
rect 7 57 9 61
rect 2 42 9 57
rect 11 55 19 70
rect 11 51 13 55
rect 17 51 19 55
rect 11 48 19 51
rect 11 44 13 48
rect 17 44 19 48
rect 11 42 19 44
rect 21 69 29 70
rect 21 65 23 69
rect 27 65 29 69
rect 21 62 29 65
rect 21 58 23 62
rect 27 58 29 62
rect 21 42 29 58
rect 43 69 51 70
rect 43 65 45 69
rect 49 65 51 69
rect 43 62 51 65
rect 43 58 45 62
rect 49 58 51 62
rect 43 42 51 58
rect 53 42 58 70
rect 60 47 68 70
rect 60 43 62 47
rect 66 43 68 47
rect 60 42 68 43
rect 70 62 78 70
rect 70 58 72 62
rect 76 58 78 62
rect 70 55 78 58
rect 70 51 72 55
rect 76 51 78 55
rect 70 42 78 51
rect 80 47 88 70
rect 80 43 82 47
rect 86 43 88 47
rect 80 42 88 43
rect 90 42 95 70
rect 97 66 102 70
rect 106 66 111 70
rect 97 63 111 66
rect 97 59 102 63
rect 106 59 111 63
rect 97 42 111 59
rect 113 62 121 70
rect 113 58 115 62
rect 119 58 121 62
rect 113 55 121 58
rect 113 51 115 55
rect 119 51 121 55
rect 113 42 121 51
rect 123 69 131 70
rect 123 65 125 69
rect 129 65 131 69
rect 123 62 131 65
rect 123 58 125 62
rect 129 58 131 62
rect 123 42 131 58
rect 133 62 141 70
rect 133 58 135 62
rect 139 58 141 62
rect 133 55 141 58
rect 133 51 135 55
rect 139 51 141 55
rect 133 42 141 51
rect 143 69 150 70
rect 143 65 145 69
rect 149 65 150 69
rect 143 62 150 65
rect 143 58 145 62
rect 149 58 150 62
rect 143 42 150 58
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect 118 78 122 82
rect 126 78 130 82
rect 134 78 138 82
rect 142 78 146 82
rect 150 78 154 82
rect -2 70 154 78
rect -2 69 102 70
rect -2 68 3 69
rect 7 68 23 69
rect 3 61 7 65
rect 22 65 23 68
rect 27 68 45 69
rect 27 65 28 68
rect 22 62 28 65
rect 22 58 23 62
rect 27 58 28 62
rect 44 65 45 68
rect 49 68 102 69
rect 49 65 50 68
rect 44 62 50 65
rect 101 66 102 68
rect 106 69 154 70
rect 106 68 125 69
rect 106 66 107 68
rect 101 63 107 66
rect 124 65 125 68
rect 129 68 145 69
rect 129 65 130 68
rect 44 58 45 62
rect 49 58 50 62
rect 72 62 76 63
rect 101 59 102 63
rect 106 59 107 63
rect 115 62 119 63
rect 3 56 7 57
rect 13 55 17 56
rect 72 55 76 58
rect 124 62 130 65
rect 144 65 145 68
rect 149 68 154 69
rect 149 65 150 68
rect 124 58 125 62
rect 129 58 130 62
rect 135 62 140 63
rect 139 58 140 62
rect 144 62 150 65
rect 144 58 145 62
rect 149 58 150 62
rect 115 55 119 58
rect 135 55 140 58
rect 13 48 17 51
rect 2 44 13 47
rect 2 43 17 44
rect 2 29 6 43
rect 26 38 30 55
rect 46 51 72 55
rect 76 51 115 55
rect 119 51 135 55
rect 139 51 140 55
rect 46 46 50 51
rect 35 42 36 46
rect 40 42 50 46
rect 57 43 62 47
rect 66 43 82 47
rect 86 43 87 47
rect 57 42 87 43
rect 15 34 16 38
rect 20 34 65 38
rect 69 34 71 38
rect 82 30 87 42
rect 102 38 106 51
rect 146 46 150 55
rect 111 42 150 46
rect 111 38 117 42
rect 145 38 150 42
rect 111 34 112 38
rect 116 34 117 38
rect 121 34 122 38
rect 126 34 127 38
rect 73 29 98 30
rect 2 25 3 29
rect 7 25 23 29
rect 27 25 43 29
rect 47 25 55 29
rect 59 25 60 29
rect 73 25 93 29
rect 97 25 98 29
rect 3 22 7 25
rect 23 22 27 25
rect 73 22 78 25
rect 3 17 7 18
rect 12 17 13 21
rect 17 17 18 21
rect 32 18 33 22
rect 37 18 73 22
rect 77 18 78 22
rect 102 21 106 34
rect 121 30 127 34
rect 149 34 150 38
rect 145 33 150 34
rect 121 26 135 30
rect 142 26 146 27
rect 23 17 27 18
rect 82 17 83 21
rect 87 17 125 21
rect 129 17 130 21
rect 142 18 146 22
rect 12 12 18 17
rect 142 12 146 14
rect -2 8 107 12
rect 111 8 154 12
rect -2 2 154 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 122 2
rect 126 -2 130 2
rect 134 -2 138 2
rect 142 -2 146 2
rect 150 -2 154 2
<< ntransistor >>
rect 9 16 11 30
rect 19 16 21 30
rect 29 16 31 30
rect 39 16 41 30
rect 79 11 81 28
rect 89 11 91 30
rect 114 12 116 30
rect 121 12 123 30
rect 131 12 133 30
rect 138 12 140 30
<< ptransistor >>
rect 9 42 11 70
rect 19 42 21 70
rect 51 42 53 70
rect 58 42 60 70
rect 68 42 70 70
rect 78 42 80 70
rect 88 42 90 70
rect 95 42 97 70
rect 111 42 113 70
rect 121 42 123 70
rect 131 42 133 70
rect 141 42 143 70
<< polycontact >>
rect 36 42 40 46
rect 16 34 20 38
rect 65 34 69 38
rect 55 25 59 29
rect 102 34 106 38
rect 112 34 116 38
rect 122 34 126 38
rect 145 34 149 38
<< ndcontact >>
rect 3 25 7 29
rect 3 18 7 22
rect 13 17 17 21
rect 23 25 27 29
rect 23 18 27 22
rect 33 18 37 22
rect 43 25 47 29
rect 73 18 77 22
rect 83 17 87 21
rect 93 25 97 29
rect 125 17 129 21
rect 142 22 146 26
rect 142 14 146 18
rect 107 8 111 12
<< pdcontact >>
rect 3 65 7 69
rect 3 57 7 61
rect 13 51 17 55
rect 13 44 17 48
rect 23 65 27 69
rect 23 58 27 62
rect 45 65 49 69
rect 45 58 49 62
rect 62 43 66 47
rect 72 58 76 62
rect 72 51 76 55
rect 82 43 86 47
rect 102 66 106 70
rect 102 59 106 63
rect 115 58 119 62
rect 115 51 119 55
rect 125 65 129 69
rect 125 58 129 62
rect 135 58 139 62
rect 135 51 139 55
rect 145 65 149 69
rect 145 58 149 62
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
rect 90 -2 94 2
rect 98 -2 102 2
rect 106 -2 110 2
rect 114 -2 118 2
rect 122 -2 126 2
rect 130 -2 134 2
rect 138 -2 142 2
rect 146 -2 150 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
rect 90 78 94 82
rect 98 78 102 82
rect 106 78 110 82
rect 114 78 118 82
rect 122 78 126 82
rect 130 78 134 82
rect 138 78 142 82
rect 146 78 150 82
<< psubstratepdiff >>
rect 0 2 152 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 122 2
rect 126 -2 130 2
rect 134 -2 138 2
rect 142 -2 146 2
rect 150 -2 152 2
rect 0 -3 152 -2
<< nsubstratendiff >>
rect 0 82 152 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect 118 78 122 82
rect 126 78 130 82
rect 134 78 138 82
rect 142 78 146 82
rect 150 78 152 82
rect 0 77 152 78
<< labels >>
rlabel polysilicon 38 40 38 40 6 an
rlabel polycontact 57 27 57 27 6 bn
rlabel polycontact 104 36 104 36 6 an
rlabel metal1 25 23 25 23 6 bn
rlabel metal1 5 23 5 23 6 bn
rlabel metal1 20 36 20 36 6 b
rlabel metal1 15 49 15 49 6 bn
rlabel ndcontact 36 20 36 20 6 z
rlabel metal1 44 20 44 20 6 z
rlabel metal1 52 20 52 20 6 z
rlabel metal1 28 44 28 44 6 b
rlabel metal1 42 44 42 44 6 an
rlabel metal1 36 36 36 36 6 b
rlabel metal1 44 36 44 36 6 b
rlabel metal1 52 36 52 36 6 b
rlabel metal1 76 6 76 6 6 vss
rlabel metal1 60 20 60 20 6 z
rlabel metal1 31 27 31 27 6 bn
rlabel metal1 68 20 68 20 6 z
rlabel metal1 76 28 76 28 6 z
rlabel metal1 60 36 60 36 6 b
rlabel metal1 60 44 60 44 6 z
rlabel polycontact 68 36 68 36 6 b
rlabel metal1 68 44 68 44 6 z
rlabel metal1 76 44 76 44 6 z
rlabel metal1 84 36 84 36 6 z
rlabel metal1 74 57 74 57 6 an
rlabel metal1 76 74 76 74 6 vdd
rlabel metal1 92 28 92 28 6 z
rlabel metal1 116 44 116 44 6 a1
rlabel polycontact 104 36 104 36 6 an
rlabel metal1 117 57 117 57 6 an
rlabel metal1 106 19 106 19 6 an
rlabel metal1 132 28 132 28 6 a2
rlabel metal1 124 32 124 32 6 a2
rlabel metal1 124 44 124 44 6 a1
rlabel metal1 148 44 148 44 6 a1
rlabel metal1 132 44 132 44 6 a1
rlabel metal1 140 44 140 44 6 a1
rlabel metal1 93 53 93 53 6 an
rlabel metal1 137 57 137 57 6 an
<< end >>
