magic
tech scmos
timestamp 1185094774
<< checkpaint >>
rect -22 -22 92 122
<< ab >>
rect 0 0 70 100
<< pwell >>
rect -4 -4 74 48
<< nwell >>
rect -4 48 74 104
<< polysilicon >>
rect 13 94 15 98
rect 21 94 23 98
rect 29 94 31 98
rect 41 94 43 98
rect 49 94 51 98
rect 57 94 59 98
rect 13 39 15 55
rect 21 46 23 55
rect 29 52 31 55
rect 41 52 43 55
rect 49 52 51 55
rect 57 52 59 55
rect 29 50 43 52
rect 21 45 33 46
rect 21 44 28 45
rect 27 41 28 44
rect 32 41 33 45
rect 27 40 33 41
rect 13 38 23 39
rect 13 37 18 38
rect 17 34 18 37
rect 22 34 23 38
rect 17 33 23 34
rect 17 22 19 33
rect 29 22 31 40
rect 41 33 43 50
rect 47 51 53 52
rect 47 47 48 51
rect 52 47 53 51
rect 47 46 53 47
rect 57 51 63 52
rect 57 47 58 51
rect 62 47 63 51
rect 57 46 63 47
rect 37 32 43 33
rect 37 28 38 32
rect 42 28 43 32
rect 37 27 43 28
rect 41 22 43 27
rect 17 2 19 7
rect 29 2 31 7
rect 41 2 43 7
<< ndiffusion >>
rect 9 21 17 22
rect 9 17 10 21
rect 14 17 17 21
rect 9 16 17 17
rect 12 7 17 16
rect 19 12 29 22
rect 19 8 22 12
rect 26 8 29 12
rect 19 7 29 8
rect 31 21 41 22
rect 31 17 34 21
rect 38 17 41 21
rect 31 7 41 17
rect 43 20 52 22
rect 43 16 46 20
rect 50 16 52 20
rect 43 12 52 16
rect 43 8 46 12
rect 50 8 52 12
rect 43 7 52 8
<< pdiffusion >>
rect 4 92 13 94
rect 4 88 6 92
rect 10 88 13 92
rect 4 82 13 88
rect 4 78 6 82
rect 10 78 13 82
rect 4 55 13 78
rect 15 55 21 94
rect 23 55 29 94
rect 31 82 41 94
rect 31 78 34 82
rect 38 78 41 82
rect 31 73 41 78
rect 31 69 34 73
rect 38 69 41 73
rect 31 55 41 69
rect 43 55 49 94
rect 51 55 57 94
rect 59 92 67 94
rect 59 88 62 92
rect 66 88 67 92
rect 59 82 67 88
rect 59 78 62 82
rect 66 78 67 82
rect 59 55 67 78
<< metal1 >>
rect -2 92 72 100
rect -2 88 6 92
rect 10 88 62 92
rect 66 88 72 92
rect 6 82 10 88
rect 6 77 10 78
rect 34 82 38 83
rect 34 73 38 78
rect 62 82 66 88
rect 62 77 66 78
rect 8 69 34 73
rect 8 68 38 69
rect 8 22 12 68
rect 17 58 63 62
rect 17 38 22 58
rect 17 34 18 38
rect 17 27 22 34
rect 28 51 53 53
rect 28 47 48 51
rect 52 47 53 51
rect 57 51 63 58
rect 57 47 58 51
rect 62 47 63 51
rect 28 45 32 47
rect 28 27 32 41
rect 58 33 62 43
rect 38 32 62 33
rect 42 28 62 32
rect 38 27 62 28
rect 8 21 39 22
rect 8 17 10 21
rect 14 17 34 21
rect 38 17 39 21
rect 46 20 50 21
rect 58 17 62 27
rect 46 12 50 16
rect -2 8 22 12
rect 26 8 46 12
rect 50 8 72 12
rect -2 4 60 8
rect 64 4 72 8
rect -2 0 72 4
<< ntransistor >>
rect 17 7 19 22
rect 29 7 31 22
rect 41 7 43 22
<< ptransistor >>
rect 13 55 15 94
rect 21 55 23 94
rect 29 55 31 94
rect 41 55 43 94
rect 49 55 51 94
rect 57 55 59 94
<< polycontact >>
rect 28 41 32 45
rect 18 34 22 38
rect 48 47 52 51
rect 58 47 62 51
rect 38 28 42 32
<< ndcontact >>
rect 10 17 14 21
rect 22 8 26 12
rect 34 17 38 21
rect 46 16 50 20
rect 46 8 50 12
<< pdcontact >>
rect 6 88 10 92
rect 6 78 10 82
rect 34 78 38 82
rect 34 69 38 73
rect 62 88 66 92
rect 62 78 66 82
<< psubstratepcontact >>
rect 60 4 64 8
<< psubstratepdiff >>
rect 59 8 65 9
rect 59 4 60 8
rect 64 4 65 8
rect 59 3 65 4
<< labels >>
rlabel metal1 20 20 20 20 6 z
rlabel metal1 10 45 10 45 6 z
rlabel metal1 20 45 20 45 6 a
rlabel metal1 20 70 20 70 6 z
rlabel metal1 35 6 35 6 6 vss
rlabel metal1 30 20 30 20 6 z
rlabel metal1 30 40 30 40 6 b
rlabel metal1 30 60 30 60 6 a
rlabel metal1 30 70 30 70 6 z
rlabel metal1 35 94 35 94 6 vdd
rlabel polycontact 40 30 40 30 6 c
rlabel metal1 50 30 50 30 6 c
rlabel metal1 40 50 40 50 6 b
rlabel polycontact 50 50 50 50 6 b
rlabel metal1 50 60 50 60 6 a
rlabel metal1 40 60 40 60 6 a
rlabel metal1 60 30 60 30 6 c
rlabel metal1 60 55 60 55 6 a
<< end >>
