magic
tech scmos
timestamp 1179387711
<< checkpaint >>
rect -22 -22 126 94
<< ab >>
rect 0 0 104 72
<< pwell >>
rect -4 -4 108 32
<< nwell >>
rect -4 32 108 76
<< polysilicon >>
rect 63 66 65 70
rect 73 66 75 70
rect 83 66 85 70
rect 93 66 95 70
rect 9 61 21 63
rect 9 58 11 61
rect 19 58 21 61
rect 29 61 50 63
rect 29 58 31 61
rect 39 58 41 61
rect 48 59 50 61
rect 48 58 54 59
rect 48 54 49 58
rect 53 54 54 58
rect 48 53 54 54
rect 63 43 65 46
rect 73 43 75 46
rect 83 43 85 46
rect 93 43 95 46
rect 55 42 79 43
rect 55 41 74 42
rect 9 34 11 38
rect 19 35 21 38
rect 18 34 24 35
rect 29 34 31 38
rect 18 30 19 34
rect 23 30 24 34
rect 39 31 41 38
rect 11 26 13 30
rect 18 29 24 30
rect 18 26 20 29
rect 28 26 30 30
rect 35 29 41 31
rect 35 26 37 29
rect 55 26 57 41
rect 73 38 74 41
rect 78 38 79 42
rect 73 37 79 38
rect 83 42 95 43
rect 83 38 90 42
rect 94 38 95 42
rect 83 37 95 38
rect 63 34 69 35
rect 63 30 64 34
rect 68 30 69 34
rect 63 29 69 30
rect 65 26 67 29
rect 75 26 77 37
rect 85 26 87 37
rect 11 4 13 13
rect 18 10 20 13
rect 28 10 30 13
rect 18 8 30 10
rect 35 4 37 13
rect 55 11 57 16
rect 11 2 37 4
rect 85 11 87 16
rect 65 2 67 6
rect 75 2 77 6
<< ndiffusion >>
rect 3 18 11 26
rect 3 14 5 18
rect 9 14 11 18
rect 3 13 11 14
rect 13 13 18 26
rect 20 25 28 26
rect 20 21 22 25
rect 26 21 28 25
rect 20 18 28 21
rect 20 14 22 18
rect 26 14 28 18
rect 20 13 28 14
rect 30 13 35 26
rect 37 18 55 26
rect 37 14 39 18
rect 43 16 55 18
rect 57 25 65 26
rect 57 21 59 25
rect 63 21 65 25
rect 57 16 65 21
rect 43 14 53 16
rect 37 13 53 14
rect 60 6 65 16
rect 67 25 75 26
rect 67 21 69 25
rect 73 21 75 25
rect 67 18 75 21
rect 67 14 69 18
rect 73 14 75 18
rect 67 6 75 14
rect 77 25 85 26
rect 77 21 79 25
rect 83 21 85 25
rect 77 16 85 21
rect 87 16 96 26
rect 77 6 82 16
rect 89 12 90 16
rect 94 12 96 16
rect 89 11 96 12
<< pdiffusion >>
rect 56 65 63 66
rect 56 61 57 65
rect 61 61 63 65
rect 4 51 9 58
rect 2 50 9 51
rect 2 46 3 50
rect 7 46 9 50
rect 2 43 9 46
rect 2 39 3 43
rect 7 39 9 43
rect 2 38 9 39
rect 11 57 19 58
rect 11 53 13 57
rect 17 53 19 57
rect 11 50 19 53
rect 11 46 13 50
rect 17 46 19 50
rect 11 38 19 46
rect 21 50 29 58
rect 21 46 23 50
rect 27 46 29 50
rect 21 43 29 46
rect 21 39 23 43
rect 27 39 29 43
rect 21 38 29 39
rect 31 43 39 58
rect 31 39 33 43
rect 37 39 39 43
rect 31 38 39 39
rect 41 51 46 58
rect 41 50 48 51
rect 41 46 43 50
rect 47 46 48 50
rect 56 46 63 61
rect 65 51 73 66
rect 65 47 67 51
rect 71 47 73 51
rect 65 46 73 47
rect 75 65 83 66
rect 75 61 77 65
rect 81 61 83 65
rect 75 46 83 61
rect 85 58 93 66
rect 85 54 87 58
rect 91 54 93 58
rect 85 46 93 54
rect 95 65 102 66
rect 95 61 97 65
rect 101 61 102 65
rect 95 46 102 61
rect 41 45 48 46
rect 41 38 46 45
<< metal1 >>
rect -2 65 106 72
rect -2 64 57 65
rect 56 61 57 64
rect 61 64 77 65
rect 61 61 62 64
rect 76 61 77 64
rect 81 64 97 65
rect 81 61 82 64
rect 96 61 97 64
rect 101 64 106 65
rect 101 61 102 64
rect 12 57 49 58
rect 12 53 13 57
rect 17 54 49 57
rect 53 54 87 58
rect 91 54 102 58
rect 17 53 18 54
rect 2 50 7 51
rect 2 46 3 50
rect 12 50 18 53
rect 66 50 67 51
rect 12 46 13 50
rect 17 46 18 50
rect 22 46 23 50
rect 27 46 43 50
rect 47 46 48 50
rect 54 47 67 50
rect 71 47 72 51
rect 54 46 72 47
rect 2 43 7 46
rect 2 39 3 43
rect 22 43 27 46
rect 22 42 23 43
rect 7 39 23 42
rect 2 38 27 39
rect 32 39 33 43
rect 37 39 38 43
rect 32 38 38 39
rect 54 38 58 46
rect 82 42 86 51
rect 73 38 74 42
rect 78 38 86 42
rect 90 42 94 43
rect 2 26 6 38
rect 32 34 58 38
rect 90 34 94 38
rect 18 30 19 34
rect 23 30 38 34
rect 2 25 50 26
rect 2 22 22 25
rect 26 22 50 25
rect 22 18 26 21
rect 4 14 5 18
rect 9 14 10 18
rect 4 8 10 14
rect 22 13 26 14
rect 39 18 43 19
rect 46 18 50 22
rect 54 25 58 34
rect 63 30 64 34
rect 68 30 94 34
rect 69 25 74 26
rect 98 25 102 54
rect 54 21 59 25
rect 63 21 64 25
rect 73 21 74 25
rect 78 21 79 25
rect 83 21 102 25
rect 69 18 74 21
rect 46 14 69 18
rect 73 14 74 18
rect 90 16 94 17
rect 39 8 43 14
rect 90 8 94 12
rect -2 4 44 8
rect 48 4 51 8
rect 55 4 106 8
rect -2 0 106 4
<< ntransistor >>
rect 11 13 13 26
rect 18 13 20 26
rect 28 13 30 26
rect 35 13 37 26
rect 55 16 57 26
rect 65 6 67 26
rect 75 6 77 26
rect 85 16 87 26
<< ptransistor >>
rect 9 38 11 58
rect 19 38 21 58
rect 29 38 31 58
rect 39 38 41 58
rect 63 46 65 66
rect 73 46 75 66
rect 83 46 85 66
rect 93 46 95 66
<< polycontact >>
rect 49 54 53 58
rect 19 30 23 34
rect 74 38 78 42
rect 90 38 94 42
rect 64 30 68 34
<< ndcontact >>
rect 5 14 9 18
rect 22 21 26 25
rect 22 14 26 18
rect 39 14 43 18
rect 59 21 63 25
rect 69 21 73 25
rect 69 14 73 18
rect 79 21 83 25
rect 90 12 94 16
<< pdcontact >>
rect 57 61 61 65
rect 3 46 7 50
rect 3 39 7 43
rect 13 53 17 57
rect 13 46 17 50
rect 23 46 27 50
rect 23 39 27 43
rect 33 39 37 43
rect 43 46 47 50
rect 67 47 71 51
rect 77 61 81 65
rect 87 54 91 58
rect 97 61 101 65
<< psubstratepcontact >>
rect 44 4 48 8
rect 51 4 55 8
<< psubstratepdiff >>
rect 43 8 56 9
rect 43 4 44 8
rect 48 4 51 8
rect 55 4 56 8
rect 43 3 56 4
<< labels >>
rlabel ptransistor 20 46 20 46 6 bn
rlabel polycontact 51 56 51 56 6 an
rlabel metal1 12 24 12 24 6 z
rlabel pdcontact 4 40 4 40 6 z
rlabel metal1 12 40 12 40 6 z
rlabel metal1 15 52 15 52 6 an
rlabel metal1 20 24 20 24 6 z
rlabel metal1 28 24 28 24 6 z
rlabel metal1 36 24 36 24 6 z
rlabel metal1 28 32 28 32 6 bn
rlabel metal1 20 40 20 40 6 z
rlabel metal1 28 48 28 48 6 z
rlabel metal1 36 48 36 48 6 z
rlabel metal1 52 4 52 4 6 vss
rlabel metal1 60 16 60 16 6 z
rlabel metal1 52 16 52 16 6 z
rlabel metal1 44 24 44 24 6 z
rlabel metal1 45 36 45 36 6 bn
rlabel pdcontact 44 48 44 48 6 z
rlabel metal1 52 68 52 68 6 vdd
rlabel metal1 68 16 68 16 6 z
rlabel metal1 59 23 59 23 6 bn
rlabel metal1 76 32 76 32 6 a
rlabel metal1 68 32 68 32 6 a
rlabel polycontact 76 40 76 40 6 b
rlabel pdcontact 69 48 69 48 6 bn
rlabel metal1 90 23 90 23 6 an
rlabel metal1 84 32 84 32 6 a
rlabel polycontact 92 40 92 40 6 a
rlabel metal1 84 48 84 48 6 b
rlabel metal1 57 56 57 56 6 an
<< end >>
