magic
tech scmos
timestamp 1185039123
<< checkpaint >>
rect -22 -24 182 124
<< ab >>
rect 0 0 160 100
<< pwell >>
rect -2 -4 162 49
<< nwell >>
rect -2 49 162 104
<< polysilicon >>
rect 11 95 13 98
rect 23 95 25 98
rect 47 95 49 98
rect 59 95 61 98
rect 71 95 73 98
rect 83 95 85 98
rect 111 95 113 98
rect 123 95 125 98
rect 135 95 137 98
rect 147 95 149 98
rect 11 53 13 55
rect 7 52 13 53
rect 7 48 8 52
rect 12 48 13 52
rect 7 47 13 48
rect 11 25 13 47
rect 23 53 25 55
rect 47 53 49 55
rect 59 53 61 55
rect 71 53 73 55
rect 83 53 85 55
rect 111 53 113 55
rect 23 52 33 53
rect 23 48 28 52
rect 32 48 33 52
rect 23 47 33 48
rect 47 52 53 53
rect 47 48 48 52
rect 52 48 53 52
rect 47 47 53 48
rect 57 52 63 53
rect 57 48 58 52
rect 62 48 63 52
rect 57 47 63 48
rect 67 52 73 53
rect 67 48 68 52
rect 72 48 73 52
rect 67 47 73 48
rect 77 52 85 53
rect 77 48 78 52
rect 82 51 85 52
rect 107 52 113 53
rect 82 48 83 51
rect 77 47 83 48
rect 107 48 108 52
rect 112 48 113 52
rect 107 47 113 48
rect 123 53 125 55
rect 123 52 129 53
rect 123 48 124 52
rect 128 48 129 52
rect 123 47 129 48
rect 23 25 25 47
rect 51 25 53 47
rect 59 25 61 47
rect 71 25 73 47
rect 79 25 81 47
rect 93 42 99 43
rect 93 38 94 42
rect 98 41 99 42
rect 135 41 137 55
rect 147 41 149 55
rect 98 39 149 41
rect 98 38 99 39
rect 93 37 99 38
rect 111 32 117 33
rect 111 28 112 32
rect 116 28 117 32
rect 111 27 117 28
rect 115 25 117 27
rect 123 32 129 33
rect 123 28 124 32
rect 128 28 129 32
rect 123 27 129 28
rect 123 25 125 27
rect 135 25 137 39
rect 147 25 149 39
rect 11 2 13 5
rect 23 2 25 5
rect 51 2 53 5
rect 59 2 61 5
rect 71 2 73 5
rect 79 2 81 5
rect 115 2 117 5
rect 123 2 125 5
rect 135 2 137 5
rect 147 2 149 5
<< ndiffusion >>
rect 3 12 11 25
rect 3 8 4 12
rect 8 8 11 12
rect 3 5 11 8
rect 13 5 23 25
rect 25 22 33 25
rect 25 18 28 22
rect 32 18 33 22
rect 25 5 33 18
rect 43 12 51 25
rect 43 8 44 12
rect 48 8 51 12
rect 43 5 51 8
rect 53 5 59 25
rect 61 22 71 25
rect 61 18 64 22
rect 68 18 71 22
rect 61 5 71 18
rect 73 5 79 25
rect 81 12 89 25
rect 107 22 115 25
rect 107 18 108 22
rect 112 18 115 22
rect 81 8 84 12
rect 88 8 89 12
rect 81 5 89 8
rect 107 5 115 18
rect 117 5 123 25
rect 125 12 135 25
rect 125 8 128 12
rect 132 8 135 12
rect 125 5 135 8
rect 137 22 147 25
rect 137 18 140 22
rect 144 18 147 22
rect 137 5 147 18
rect 149 22 157 25
rect 149 18 152 22
rect 156 18 157 22
rect 149 12 157 18
rect 149 8 152 12
rect 156 8 157 12
rect 149 5 157 8
<< pdiffusion >>
rect 3 82 11 95
rect 3 78 4 82
rect 8 78 11 82
rect 3 72 11 78
rect 3 68 4 72
rect 8 68 11 72
rect 3 55 11 68
rect 13 72 23 95
rect 13 68 16 72
rect 20 68 23 72
rect 13 55 23 68
rect 25 82 33 95
rect 25 78 28 82
rect 32 78 33 82
rect 25 72 33 78
rect 25 68 28 72
rect 32 68 33 72
rect 25 55 33 68
rect 39 82 47 95
rect 39 78 40 82
rect 44 78 47 82
rect 39 55 47 78
rect 49 72 59 95
rect 49 68 52 72
rect 56 68 59 72
rect 49 55 59 68
rect 61 82 71 95
rect 61 78 64 82
rect 68 78 71 82
rect 61 72 71 78
rect 61 68 64 72
rect 68 68 71 72
rect 61 55 71 68
rect 73 72 83 95
rect 73 68 76 72
rect 80 68 83 72
rect 73 55 83 68
rect 85 82 93 95
rect 85 78 88 82
rect 92 78 93 82
rect 85 55 93 78
rect 103 92 111 95
rect 103 88 104 92
rect 108 88 111 92
rect 103 82 111 88
rect 103 78 104 82
rect 108 78 111 82
rect 103 55 111 78
rect 113 82 123 95
rect 113 78 116 82
rect 120 78 123 82
rect 113 55 123 78
rect 125 92 135 95
rect 125 88 128 92
rect 132 88 135 92
rect 125 82 135 88
rect 125 78 128 82
rect 132 78 135 82
rect 125 55 135 78
rect 137 82 147 95
rect 137 78 140 82
rect 144 78 147 82
rect 137 72 147 78
rect 137 68 140 72
rect 144 68 147 72
rect 137 62 147 68
rect 137 58 140 62
rect 144 58 147 62
rect 137 55 147 58
rect 149 92 157 95
rect 149 88 152 92
rect 156 88 157 92
rect 149 82 157 88
rect 149 78 152 82
rect 156 78 157 82
rect 149 72 157 78
rect 149 68 152 72
rect 156 68 157 72
rect 149 55 157 68
<< metal1 >>
rect -2 92 162 101
rect -2 88 104 92
rect 108 88 128 92
rect 132 88 152 92
rect 156 88 162 92
rect -2 87 162 88
rect 3 82 9 83
rect 27 82 33 83
rect 3 78 4 82
rect 8 78 28 82
rect 32 78 33 82
rect 3 77 9 78
rect 27 77 33 78
rect 39 82 45 83
rect 63 82 69 83
rect 87 82 93 83
rect 39 78 40 82
rect 44 78 64 82
rect 68 78 88 82
rect 92 78 93 82
rect 39 77 45 78
rect 63 77 69 78
rect 87 77 93 78
rect 103 82 109 87
rect 103 78 104 82
rect 108 78 109 82
rect 103 77 109 78
rect 115 82 121 83
rect 115 78 116 82
rect 120 78 121 82
rect 115 77 121 78
rect 127 82 133 87
rect 127 78 128 82
rect 132 78 133 82
rect 127 77 133 78
rect 137 82 145 83
rect 137 78 140 82
rect 144 78 145 82
rect 137 77 145 78
rect 151 82 157 87
rect 151 78 152 82
rect 156 78 157 82
rect 4 73 8 77
rect 28 73 32 77
rect 64 73 68 77
rect 3 72 9 73
rect 3 68 4 72
rect 8 68 9 72
rect 3 67 9 68
rect 15 72 21 73
rect 27 72 33 73
rect 51 72 57 73
rect 15 68 16 72
rect 20 68 22 72
rect 15 67 22 68
rect 27 68 28 72
rect 32 68 52 72
rect 56 68 57 72
rect 27 67 33 68
rect 51 67 57 68
rect 63 72 69 73
rect 63 68 64 72
rect 68 68 69 72
rect 63 67 69 68
rect 75 72 81 73
rect 116 72 120 77
rect 137 73 143 77
rect 137 72 145 73
rect 75 68 76 72
rect 80 68 120 72
rect 75 67 81 68
rect 7 52 13 62
rect 7 48 8 52
rect 12 48 13 52
rect 7 18 13 48
rect 18 22 22 67
rect 27 52 33 62
rect 27 48 28 52
rect 32 48 33 52
rect 27 28 33 48
rect 47 52 53 62
rect 47 48 48 52
rect 52 48 53 52
rect 47 28 53 48
rect 57 52 63 62
rect 57 48 58 52
rect 62 48 63 52
rect 57 28 63 48
rect 67 52 73 62
rect 67 48 68 52
rect 72 48 73 52
rect 67 28 73 48
rect 77 52 83 62
rect 77 48 78 52
rect 82 48 83 52
rect 77 28 83 48
rect 107 52 113 62
rect 127 53 133 72
rect 107 48 108 52
rect 112 48 113 52
rect 93 42 99 43
rect 93 38 94 42
rect 98 38 99 42
rect 93 37 99 38
rect 27 22 33 23
rect 63 22 69 23
rect 94 22 98 37
rect 107 33 113 48
rect 123 52 133 53
rect 123 48 124 52
rect 128 48 133 52
rect 123 47 133 48
rect 127 33 133 47
rect 107 32 117 33
rect 107 28 112 32
rect 116 28 117 32
rect 108 27 117 28
rect 123 32 133 33
rect 123 28 124 32
rect 128 28 133 32
rect 137 68 140 72
rect 144 68 145 72
rect 137 67 145 68
rect 151 72 157 78
rect 151 68 152 72
rect 156 68 157 72
rect 151 67 157 68
rect 137 63 143 67
rect 137 62 145 63
rect 137 58 140 62
rect 144 58 145 62
rect 137 57 145 58
rect 123 27 132 28
rect 137 23 143 57
rect 107 22 113 23
rect 18 18 28 22
rect 32 18 64 22
rect 68 18 108 22
rect 112 18 113 22
rect 27 17 33 18
rect 63 17 69 18
rect 107 17 113 18
rect 137 22 145 23
rect 137 18 140 22
rect 144 18 145 22
rect 137 17 145 18
rect 151 22 157 23
rect 151 18 152 22
rect 156 18 157 22
rect 151 13 157 18
rect -2 12 162 13
rect -2 8 4 12
rect 8 8 44 12
rect 48 8 84 12
rect 88 10 128 12
rect 88 8 96 10
rect -2 6 96 8
rect 100 8 128 10
rect 132 8 152 12
rect 156 8 162 12
rect 100 6 162 8
rect -2 -1 162 6
<< ntransistor >>
rect 11 5 13 25
rect 23 5 25 25
rect 51 5 53 25
rect 59 5 61 25
rect 71 5 73 25
rect 79 5 81 25
rect 115 5 117 25
rect 123 5 125 25
rect 135 5 137 25
rect 147 5 149 25
<< ptransistor >>
rect 11 55 13 95
rect 23 55 25 95
rect 47 55 49 95
rect 59 55 61 95
rect 71 55 73 95
rect 83 55 85 95
rect 111 55 113 95
rect 123 55 125 95
rect 135 55 137 95
rect 147 55 149 95
<< polycontact >>
rect 8 48 12 52
rect 28 48 32 52
rect 48 48 52 52
rect 58 48 62 52
rect 68 48 72 52
rect 78 48 82 52
rect 108 48 112 52
rect 124 48 128 52
rect 94 38 98 42
rect 112 28 116 32
rect 124 28 128 32
<< ndcontact >>
rect 4 8 8 12
rect 28 18 32 22
rect 44 8 48 12
rect 64 18 68 22
rect 108 18 112 22
rect 84 8 88 12
rect 128 8 132 12
rect 140 18 144 22
rect 152 18 156 22
rect 152 8 156 12
<< pdcontact >>
rect 4 78 8 82
rect 4 68 8 72
rect 16 68 20 72
rect 28 78 32 82
rect 28 68 32 72
rect 40 78 44 82
rect 52 68 56 72
rect 64 78 68 82
rect 64 68 68 72
rect 76 68 80 72
rect 88 78 92 82
rect 104 88 108 92
rect 104 78 108 82
rect 116 78 120 82
rect 128 88 132 92
rect 128 78 132 82
rect 140 78 144 82
rect 140 68 144 72
rect 140 58 144 62
rect 152 88 156 92
rect 152 78 156 82
rect 152 68 156 72
<< psubstratepcontact >>
rect 96 6 100 10
<< psubstratepdiff >>
rect 95 10 101 17
rect 95 6 96 10
rect 100 6 101 10
rect 95 5 101 6
<< labels >>
rlabel metal1 10 40 10 40 6 i7
rlabel metal1 10 40 10 40 6 i7
rlabel metal1 30 45 30 45 6 i6
rlabel metal1 30 45 30 45 6 i6
rlabel metal1 50 45 50 45 6 i5
rlabel metal1 60 45 60 45 6 i4
rlabel metal1 60 45 60 45 6 i4
rlabel metal1 50 45 50 45 6 i5
rlabel metal1 80 6 80 6 6 vss
rlabel metal1 80 6 80 6 6 vss
rlabel metal1 80 45 80 45 6 i2
rlabel metal1 70 45 70 45 6 i3
rlabel metal1 70 45 70 45 6 i3
rlabel metal1 80 45 80 45 6 i2
rlabel metal1 80 94 80 94 6 vdd
rlabel metal1 80 94 80 94 6 vdd
rlabel metal1 110 45 110 45 6 i1
rlabel metal1 110 45 110 45 6 i1
rlabel metal1 130 50 130 50 6 i0
rlabel metal1 130 50 130 50 6 i0
rlabel metal1 140 50 140 50 6 q
rlabel metal1 140 50 140 50 6 q
<< end >>
