.subckt nd2v5x1 a b vdd vss z
*   SPICE3 file   created from nd2v5x1.ext -      technology: scmos
m00 z      b      vdd    vdd p w=19u  l=2.3636u ad=76p      pd=27u      as=158p     ps=56u
m01 vdd    a      z      vdd p w=19u  l=2.3636u ad=158p     pd=56u      as=76p      ps=27u
m02 w1     b      z      vss n w=12u  l=2.3636u ad=30p      pd=17u      as=72p      ps=38u
m03 vss    a      w1     vss n w=12u  l=2.3636u ad=144p     pd=48u      as=30p      ps=17u
C0  a      b      0.105f
C1  z      vdd    0.182f
C2  b      vdd    0.020f
C3  vss    z      0.045f
C4  vss    b      0.020f
C5  z      b      0.144f
C6  a      vdd    0.016f
C7  vss    w1     0.004f
C8  vss    a      0.063f
C9  z      a      0.038f
C10 vss    vdd    0.005f
C12 z      vss    0.009f
C13 a      vss    0.024f
C14 b      vss    0.021f
.ends
