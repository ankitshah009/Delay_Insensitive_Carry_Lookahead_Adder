magic
tech scmos
timestamp 1180600706
<< checkpaint >>
rect -22 -22 142 122
<< ab >>
rect 0 0 120 100
<< pwell >>
rect -4 -4 124 48
<< nwell >>
rect -4 48 124 104
<< polysilicon >>
rect 27 94 29 98
rect 39 94 41 98
rect 51 94 53 98
rect 59 94 61 98
rect 71 94 73 98
rect 83 94 85 98
rect 91 94 93 98
rect 15 70 17 74
rect 15 53 17 56
rect 7 52 17 53
rect 7 48 8 52
rect 12 48 17 52
rect 7 47 17 48
rect 15 37 17 47
rect 27 53 29 75
rect 39 73 41 76
rect 33 72 41 73
rect 33 68 34 72
rect 38 68 41 72
rect 33 67 41 68
rect 27 52 33 53
rect 27 48 28 52
rect 32 48 33 52
rect 27 47 33 48
rect 15 25 17 29
rect 27 23 29 47
rect 39 41 41 67
rect 51 63 53 75
rect 47 62 53 63
rect 47 58 48 62
rect 52 58 53 62
rect 47 57 53 58
rect 47 52 53 53
rect 47 48 48 52
rect 52 51 53 52
rect 59 51 61 75
rect 71 73 73 76
rect 83 73 85 76
rect 52 49 61 51
rect 52 48 53 49
rect 47 47 53 48
rect 39 39 53 41
rect 33 32 41 33
rect 33 28 34 32
rect 38 28 41 32
rect 33 27 41 28
rect 39 23 41 27
rect 51 23 53 39
rect 59 23 61 49
rect 69 71 73 73
rect 79 71 85 73
rect 69 33 71 71
rect 79 53 81 71
rect 91 63 93 76
rect 103 69 105 73
rect 85 62 93 63
rect 85 58 86 62
rect 90 58 93 62
rect 85 57 93 58
rect 75 52 81 53
rect 75 48 76 52
rect 80 51 81 52
rect 103 51 105 55
rect 80 49 105 51
rect 80 48 81 49
rect 75 47 81 48
rect 79 39 81 47
rect 65 32 71 33
rect 65 28 66 32
rect 70 28 71 32
rect 65 27 71 28
rect 75 37 81 39
rect 85 42 93 43
rect 85 38 86 42
rect 90 38 93 42
rect 85 37 93 38
rect 103 37 105 49
rect 75 23 77 37
rect 81 32 87 33
rect 81 28 82 32
rect 86 28 87 32
rect 81 27 87 28
rect 71 21 77 23
rect 71 18 73 21
rect 83 19 85 27
rect 91 19 93 37
rect 103 25 105 29
rect 27 7 29 11
rect 39 7 41 11
rect 51 7 53 11
rect 59 7 61 11
rect 71 2 73 6
rect 83 3 85 7
rect 91 3 93 7
<< ndiffusion >>
rect 7 29 15 37
rect 17 34 25 37
rect 17 30 20 34
rect 24 30 25 34
rect 17 29 25 30
rect 7 22 13 29
rect 43 32 49 33
rect 43 28 44 32
rect 48 28 49 32
rect 43 23 49 28
rect 7 18 8 22
rect 12 18 13 22
rect 7 17 13 18
rect 19 22 27 23
rect 19 18 20 22
rect 24 18 27 22
rect 19 11 27 18
rect 29 11 39 23
rect 41 11 51 23
rect 53 11 59 23
rect 61 22 69 23
rect 61 18 64 22
rect 68 18 69 22
rect 95 34 103 37
rect 95 30 96 34
rect 100 30 103 34
rect 95 29 103 30
rect 105 29 113 37
rect 95 22 101 23
rect 95 19 96 22
rect 78 18 83 19
rect 61 11 71 18
rect 63 6 71 11
rect 73 12 83 18
rect 73 8 76 12
rect 80 8 83 12
rect 73 7 83 8
rect 85 7 91 19
rect 93 18 96 19
rect 100 18 101 22
rect 93 7 101 18
rect 107 12 113 29
rect 107 8 108 12
rect 112 8 113 12
rect 107 7 113 8
rect 73 6 80 7
<< pdiffusion >>
rect 7 82 13 83
rect 7 78 8 82
rect 12 78 13 82
rect 7 70 13 78
rect 19 82 27 94
rect 19 78 20 82
rect 24 78 27 82
rect 19 75 27 78
rect 29 76 39 94
rect 41 76 51 94
rect 29 75 34 76
rect 7 56 15 70
rect 17 62 25 70
rect 17 58 20 62
rect 24 58 25 62
rect 17 56 25 58
rect 43 75 51 76
rect 53 75 59 94
rect 61 82 71 94
rect 61 78 64 82
rect 68 78 71 82
rect 61 76 71 78
rect 73 92 83 94
rect 73 88 76 92
rect 80 88 83 92
rect 73 76 83 88
rect 85 76 91 94
rect 93 82 101 94
rect 93 78 96 82
rect 100 78 101 82
rect 93 76 101 78
rect 107 82 113 83
rect 107 78 108 82
rect 112 78 113 82
rect 61 75 66 76
rect 43 72 49 75
rect 43 68 44 72
rect 48 68 49 72
rect 43 67 49 68
rect 107 69 113 78
rect 95 62 103 69
rect 95 58 96 62
rect 100 58 103 62
rect 95 55 103 58
rect 105 55 113 69
<< metal1 >>
rect -2 92 122 100
rect -2 88 76 92
rect 80 88 122 92
rect 8 82 12 88
rect 96 82 100 83
rect 19 78 20 82
rect 24 78 64 82
rect 68 78 69 82
rect 8 77 12 78
rect 8 72 12 73
rect 96 72 100 78
rect 108 82 112 88
rect 108 77 112 78
rect 108 72 112 73
rect 8 68 34 72
rect 38 68 39 72
rect 43 68 44 72
rect 48 68 112 72
rect 8 52 12 68
rect 8 27 12 48
rect 18 58 20 62
rect 24 58 48 62
rect 52 58 53 62
rect 18 34 22 58
rect 28 52 32 53
rect 39 48 48 52
rect 52 48 53 52
rect 28 41 32 48
rect 58 42 62 68
rect 44 38 62 42
rect 68 52 72 63
rect 86 62 90 63
rect 77 58 86 62
rect 95 58 96 62
rect 100 58 102 62
rect 86 52 90 58
rect 68 48 76 52
rect 80 48 81 52
rect 86 48 93 52
rect 18 30 20 34
rect 24 32 25 34
rect 44 32 48 38
rect 68 37 72 48
rect 86 42 90 48
rect 77 38 86 42
rect 86 37 90 38
rect 98 34 102 58
rect 95 32 96 34
rect 24 30 34 32
rect 18 28 34 30
rect 38 28 39 32
rect 65 28 66 32
rect 70 28 82 32
rect 86 30 96 32
rect 100 30 102 34
rect 86 28 102 30
rect 44 27 48 28
rect 8 22 12 23
rect 108 22 112 68
rect 19 18 20 22
rect 24 18 64 22
rect 68 18 69 22
rect 95 18 96 22
rect 100 18 112 22
rect 8 12 12 18
rect 108 17 112 18
rect -2 8 76 12
rect 80 8 108 12
rect 112 8 122 12
rect -2 0 122 8
<< ntransistor >>
rect 15 29 17 37
rect 27 11 29 23
rect 39 11 41 23
rect 51 11 53 23
rect 59 11 61 23
rect 103 29 105 37
rect 71 6 73 18
rect 83 7 85 19
rect 91 7 93 19
<< ptransistor >>
rect 27 75 29 94
rect 39 76 41 94
rect 15 56 17 70
rect 51 75 53 94
rect 59 75 61 94
rect 71 76 73 94
rect 83 76 85 94
rect 91 76 93 94
rect 103 55 105 69
<< polycontact >>
rect 8 48 12 52
rect 34 68 38 72
rect 28 48 32 52
rect 48 58 52 62
rect 48 48 52 52
rect 34 28 38 32
rect 86 58 90 62
rect 76 48 80 52
rect 66 28 70 32
rect 86 38 90 42
rect 82 28 86 32
<< ndcontact >>
rect 20 30 24 34
rect 44 28 48 32
rect 8 18 12 22
rect 20 18 24 22
rect 64 18 68 22
rect 96 30 100 34
rect 76 8 80 12
rect 96 18 100 22
rect 108 8 112 12
<< pdcontact >>
rect 8 78 12 82
rect 20 78 24 82
rect 20 58 24 62
rect 64 78 68 82
rect 76 88 80 92
rect 96 78 100 82
rect 108 78 112 82
rect 44 68 48 72
rect 96 58 100 62
<< labels >>
rlabel polycontact 10 50 10 50 6 cmd1
rlabel polycontact 30 50 30 50 6 i2
rlabel metal1 20 70 20 70 6 cmd1
rlabel metal1 30 70 30 70 6 cmd1
rlabel metal1 60 6 60 6 6 vss
rlabel metal1 50 40 50 40 6 nq
rlabel polycontact 50 50 50 50 6 i1
rlabel metal1 60 50 60 50 6 nq
rlabel metal1 60 60 60 60 6 nq
rlabel metal1 50 70 50 70 6 nq
rlabel metal1 60 70 60 70 6 nq
rlabel metal1 60 94 60 94 6 vdd
rlabel metal1 80 40 80 40 6 i0
rlabel metal1 70 50 70 50 6 cmd0
rlabel metal1 90 50 90 50 6 i0
rlabel metal1 80 60 80 60 6 i0
rlabel metal1 70 70 70 70 6 nq
rlabel metal1 80 70 80 70 6 nq
rlabel metal1 90 70 90 70 6 nq
rlabel metal1 100 20 100 20 6 nq
rlabel metal1 110 45 110 45 6 nq
rlabel metal1 100 70 100 70 6 nq
<< end >>
