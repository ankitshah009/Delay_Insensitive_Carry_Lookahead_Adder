magic
tech scmos
timestamp 1179387521
<< checkpaint >>
rect -22 -25 190 105
<< ab >>
rect 0 0 168 80
<< pwell >>
rect -4 -7 172 36
<< nwell >>
rect -4 36 172 87
<< polysilicon >>
rect 9 70 11 74
rect 16 70 18 74
rect 26 70 28 74
rect 33 70 35 74
rect 43 70 45 74
rect 50 70 52 74
rect 60 70 62 74
rect 67 70 69 74
rect 77 70 79 74
rect 87 70 89 74
rect 117 70 119 74
rect 127 70 129 74
rect 137 70 139 74
rect 147 70 149 74
rect 97 61 99 65
rect 107 61 109 65
rect 157 61 159 65
rect 9 39 11 42
rect 16 39 18 42
rect 26 39 28 42
rect 33 39 35 42
rect 43 39 45 42
rect 5 38 11 39
rect 5 34 6 38
rect 10 34 11 38
rect 5 33 11 34
rect 15 37 28 39
rect 32 38 45 39
rect 15 22 17 37
rect 32 34 33 38
rect 37 37 45 38
rect 50 39 52 42
rect 60 39 62 42
rect 67 39 69 42
rect 77 39 79 42
rect 87 39 89 42
rect 97 39 99 42
rect 50 37 62 39
rect 66 38 72 39
rect 37 34 38 37
rect 32 33 38 34
rect 26 29 28 33
rect 36 29 38 33
rect 46 29 48 33
rect 56 29 58 37
rect 66 34 67 38
rect 71 34 72 38
rect 66 33 72 34
rect 76 38 99 39
rect 76 37 94 38
rect 66 29 68 33
rect 76 29 78 37
rect 88 34 94 37
rect 98 34 99 38
rect 88 33 99 34
rect 107 39 109 42
rect 117 39 119 42
rect 127 39 129 42
rect 137 39 139 42
rect 147 39 149 42
rect 157 39 159 42
rect 107 38 129 39
rect 107 34 122 38
rect 126 34 129 38
rect 107 33 129 34
rect 133 38 159 39
rect 133 34 134 38
rect 138 37 159 38
rect 138 34 139 37
rect 133 33 139 34
rect 88 29 90 33
rect 109 30 111 33
rect 119 30 121 33
rect 11 21 17 22
rect 11 17 12 21
rect 16 17 17 21
rect 11 16 17 17
rect 15 8 17 16
rect 26 15 28 18
rect 36 15 38 18
rect 26 13 38 15
rect 46 8 48 11
rect 56 8 58 11
rect 66 8 68 13
rect 15 6 58 8
rect 76 6 78 10
rect 88 6 90 10
rect 109 6 111 11
rect 119 6 121 11
<< ndiffusion >>
rect 19 28 26 29
rect 19 24 20 28
rect 24 24 26 28
rect 19 23 26 24
rect 21 18 26 23
rect 28 23 36 29
rect 28 19 30 23
rect 34 19 36 23
rect 28 18 36 19
rect 38 28 46 29
rect 38 24 40 28
rect 44 24 46 28
rect 38 18 46 24
rect 41 11 46 18
rect 48 28 56 29
rect 48 24 50 28
rect 54 24 56 28
rect 48 11 56 24
rect 58 28 66 29
rect 58 24 60 28
rect 64 24 66 28
rect 58 13 66 24
rect 68 21 76 29
rect 68 17 70 21
rect 74 17 76 21
rect 68 13 76 17
rect 58 11 63 13
rect 71 10 76 13
rect 78 12 88 29
rect 78 10 81 12
rect 80 8 81 10
rect 85 10 88 12
rect 90 22 95 29
rect 90 21 97 22
rect 90 17 92 21
rect 96 17 97 21
rect 90 16 97 17
rect 90 10 95 16
rect 101 12 109 30
rect 85 8 86 10
rect 80 7 86 8
rect 101 8 102 12
rect 106 11 109 12
rect 111 29 119 30
rect 111 25 113 29
rect 117 25 119 29
rect 111 11 119 25
rect 121 12 129 30
rect 121 11 124 12
rect 106 8 107 11
rect 101 7 107 8
rect 123 8 124 11
rect 128 8 129 12
rect 123 7 129 8
<< pdiffusion >>
rect 4 55 9 70
rect 2 54 9 55
rect 2 50 3 54
rect 7 50 9 54
rect 2 47 9 50
rect 2 43 3 47
rect 7 43 9 47
rect 2 42 9 43
rect 11 42 16 70
rect 18 69 26 70
rect 18 65 20 69
rect 24 65 26 69
rect 18 42 26 65
rect 28 42 33 70
rect 35 62 43 70
rect 35 58 37 62
rect 41 58 43 62
rect 35 47 43 58
rect 35 43 37 47
rect 41 43 43 47
rect 35 42 43 43
rect 45 42 50 70
rect 52 69 60 70
rect 52 65 54 69
rect 58 65 60 69
rect 52 42 60 65
rect 62 42 67 70
rect 69 62 77 70
rect 69 58 71 62
rect 75 58 77 62
rect 69 47 77 58
rect 69 43 71 47
rect 75 43 77 47
rect 69 42 77 43
rect 79 54 87 70
rect 79 50 81 54
rect 85 50 87 54
rect 79 47 87 50
rect 79 43 81 47
rect 85 43 87 47
rect 79 42 87 43
rect 89 61 94 70
rect 112 61 117 70
rect 89 60 97 61
rect 89 56 91 60
rect 95 56 97 60
rect 89 42 97 56
rect 99 54 107 61
rect 99 50 101 54
rect 105 50 107 54
rect 99 47 107 50
rect 99 43 101 47
rect 105 43 107 47
rect 99 42 107 43
rect 109 60 117 61
rect 109 56 111 60
rect 115 56 117 60
rect 109 42 117 56
rect 119 61 127 70
rect 119 57 121 61
rect 125 57 127 61
rect 119 54 127 57
rect 119 50 121 54
rect 125 50 127 54
rect 119 42 127 50
rect 129 69 137 70
rect 129 65 131 69
rect 135 65 137 69
rect 129 62 137 65
rect 129 58 131 62
rect 135 58 137 62
rect 129 42 137 58
rect 139 54 147 70
rect 139 50 141 54
rect 145 50 147 54
rect 139 47 147 50
rect 139 43 141 47
rect 145 43 147 47
rect 139 42 147 43
rect 149 61 154 70
rect 149 60 157 61
rect 149 56 151 60
rect 155 56 157 60
rect 149 42 157 56
rect 159 55 164 61
rect 159 54 166 55
rect 159 50 161 54
rect 165 50 166 54
rect 159 47 166 50
rect 159 43 161 47
rect 165 43 166 47
rect 159 42 166 43
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect 118 78 122 82
rect 126 78 130 82
rect 134 78 138 82
rect 142 78 146 82
rect 150 78 154 82
rect 158 78 162 82
rect 166 78 170 82
rect -2 69 170 78
rect -2 68 20 69
rect 19 65 20 68
rect 24 68 54 69
rect 24 65 25 68
rect 53 65 54 68
rect 58 68 131 69
rect 58 65 59 68
rect 17 58 37 62
rect 41 58 71 62
rect 75 60 95 62
rect 75 58 91 60
rect 17 54 23 58
rect 110 60 116 68
rect 135 68 170 69
rect 131 62 135 65
rect 110 56 111 60
rect 115 56 116 60
rect 121 61 125 62
rect 131 57 135 58
rect 151 60 155 68
rect 91 55 95 56
rect 101 54 105 55
rect 2 50 3 54
rect 7 50 23 54
rect 28 50 81 54
rect 85 50 86 54
rect 2 47 7 50
rect 2 43 3 47
rect 2 41 7 43
rect 28 38 32 50
rect 36 43 37 47
rect 5 34 6 38
rect 10 34 33 38
rect 37 34 38 38
rect 41 30 45 47
rect 19 28 45 30
rect 19 24 20 28
rect 24 26 40 28
rect 24 24 25 26
rect 39 24 40 26
rect 44 24 45 28
rect 49 28 53 50
rect 81 47 86 50
rect 59 43 71 47
rect 75 43 76 47
rect 85 46 86 47
rect 121 54 125 57
rect 151 55 155 56
rect 105 50 121 53
rect 101 49 125 50
rect 141 54 145 55
rect 101 47 105 49
rect 85 43 101 46
rect 141 47 145 50
rect 59 28 63 43
rect 81 42 105 43
rect 113 42 135 46
rect 161 54 165 55
rect 161 47 165 50
rect 145 43 161 46
rect 141 42 165 43
rect 81 38 85 42
rect 113 38 117 42
rect 131 38 135 42
rect 66 34 67 38
rect 71 34 85 38
rect 93 34 94 38
rect 98 34 117 38
rect 121 34 122 38
rect 126 34 127 38
rect 131 34 134 38
rect 138 34 139 38
rect 81 29 85 34
rect 121 30 127 34
rect 49 24 50 28
rect 54 24 55 28
rect 59 24 60 28
rect 64 24 65 28
rect 81 25 113 29
rect 117 25 118 29
rect 121 26 135 30
rect 29 21 30 23
rect 11 17 12 21
rect 16 19 30 21
rect 34 21 35 23
rect 143 21 147 42
rect 34 19 70 21
rect 16 17 70 19
rect 74 17 92 21
rect 96 17 147 21
rect -2 8 81 12
rect 85 8 102 12
rect 106 8 124 12
rect 128 8 170 12
rect -2 2 170 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 122 2
rect 126 -2 130 2
rect 134 -2 138 2
rect 142 -2 146 2
rect 150 -2 154 2
rect 158 -2 162 2
rect 166 -2 170 2
<< ntransistor >>
rect 26 18 28 29
rect 36 18 38 29
rect 46 11 48 29
rect 56 11 58 29
rect 66 13 68 29
rect 76 10 78 29
rect 88 10 90 29
rect 109 11 111 30
rect 119 11 121 30
<< ptransistor >>
rect 9 42 11 70
rect 16 42 18 70
rect 26 42 28 70
rect 33 42 35 70
rect 43 42 45 70
rect 50 42 52 70
rect 60 42 62 70
rect 67 42 69 70
rect 77 42 79 70
rect 87 42 89 70
rect 97 42 99 61
rect 107 42 109 61
rect 117 42 119 70
rect 127 42 129 70
rect 137 42 139 70
rect 147 42 149 70
rect 157 42 159 61
<< polycontact >>
rect 6 34 10 38
rect 33 34 37 38
rect 67 34 71 38
rect 94 34 98 38
rect 122 34 126 38
rect 134 34 138 38
rect 12 17 16 21
<< ndcontact >>
rect 20 24 24 28
rect 30 19 34 23
rect 40 24 44 28
rect 50 24 54 28
rect 60 24 64 28
rect 70 17 74 21
rect 81 8 85 12
rect 92 17 96 21
rect 102 8 106 12
rect 113 25 117 29
rect 124 8 128 12
<< pdcontact >>
rect 3 50 7 54
rect 3 43 7 47
rect 20 65 24 69
rect 37 58 41 62
rect 37 43 41 47
rect 54 65 58 69
rect 71 58 75 62
rect 71 43 75 47
rect 81 50 85 54
rect 81 43 85 47
rect 91 56 95 60
rect 101 50 105 54
rect 101 43 105 47
rect 111 56 115 60
rect 121 57 125 61
rect 121 50 125 54
rect 131 65 135 69
rect 131 58 135 62
rect 141 50 145 54
rect 141 43 145 47
rect 151 56 155 60
rect 161 50 165 54
rect 161 43 165 47
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
rect 90 -2 94 2
rect 98 -2 102 2
rect 106 -2 110 2
rect 114 -2 118 2
rect 122 -2 126 2
rect 130 -2 134 2
rect 138 -2 142 2
rect 146 -2 150 2
rect 154 -2 158 2
rect 162 -2 166 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
rect 90 78 94 82
rect 98 78 102 82
rect 106 78 110 82
rect 114 78 118 82
rect 122 78 126 82
rect 130 78 134 82
rect 138 78 142 82
rect 146 78 150 82
rect 154 78 158 82
rect 162 78 166 82
<< psubstratepdiff >>
rect 0 2 168 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 122 2
rect 126 -2 130 2
rect 134 -2 138 2
rect 142 -2 146 2
rect 150 -2 154 2
rect 158 -2 162 2
rect 166 -2 168 2
rect 0 -3 168 -2
<< nsubstratendiff >>
rect 0 82 168 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect 118 78 122 82
rect 126 78 130 82
rect 134 78 138 82
rect 142 78 146 82
rect 150 78 154 82
rect 158 78 162 82
rect 166 78 168 82
rect 0 77 168 78
<< labels >>
rlabel polycontact 14 19 14 19 6 bn
rlabel polycontact 8 36 8 36 6 an
rlabel ptransistor 34 53 34 53 6 an
rlabel ptransistor 68 53 68 53 6 an
rlabel pdcontact 4 44 4 44 6 z
rlabel metal1 12 52 12 52 6 z
rlabel metal1 28 60 28 60 6 z
rlabel metal1 20 56 20 56 6 z
rlabel metal1 21 36 21 36 6 an
rlabel metal1 51 39 51 39 6 an
rlabel metal1 60 60 60 60 6 z
rlabel metal1 52 60 52 60 6 z
rlabel metal1 44 60 44 60 6 z
rlabel metal1 36 60 36 60 6 z
rlabel metal1 84 6 84 6 6 vss
rlabel metal1 75 36 75 36 6 an
rlabel metal1 83 39 83 39 6 an
rlabel metal1 68 60 68 60 6 z
rlabel metal1 92 60 92 60 6 z
rlabel metal1 84 60 84 60 6 z
rlabel metal1 76 60 76 60 6 z
rlabel metal1 84 74 84 74 6 vdd
rlabel metal1 99 27 99 27 6 an
rlabel metal1 132 28 132 28 6 a
rlabel metal1 124 32 124 32 6 a
rlabel metal1 100 36 100 36 6 b
rlabel metal1 132 44 132 44 6 b
rlabel metal1 124 44 124 44 6 b
rlabel metal1 116 44 116 44 6 b
rlabel metal1 108 36 108 36 6 b
rlabel metal1 123 55 123 55 6 an
rlabel metal1 103 48 103 48 6 an
rlabel metal1 79 19 79 19 6 bn
rlabel metal1 163 48 163 48 6 bn
rlabel metal1 143 48 143 48 6 bn
<< end >>
