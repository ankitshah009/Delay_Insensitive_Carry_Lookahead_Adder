.subckt aoi22v0x1 a1 a2 b1 b2 vdd vss z
*   SPICE3 file   created from aoi22v0x1.ext -      technology: scmos
m00 z      b1     n3     vdd p w=27u  l=2.3636u ad=108p     pd=35u      as=127.5p   ps=51.5u
m01 n3     b2     z      vdd p w=27u  l=2.3636u ad=127.5p   pd=51.5u    as=108p     ps=35u
m02 vdd    a2     n3     vdd p w=27u  l=2.3636u ad=135p     pd=37u      as=127.5p   ps=51.5u
m03 n3     a1     vdd    vdd p w=27u  l=2.3636u ad=127.5p   pd=51.5u    as=135p     ps=37u
m04 w1     b1     vss    vss n w=12u  l=2.3636u ad=36p      pd=18u      as=116p     ps=45u
m05 z      b2     w1     vss n w=12u  l=2.3636u ad=48p      pd=20u      as=36p      ps=18u
m06 w2     a2     z      vss n w=12u  l=2.3636u ad=36p      pd=18u      as=48p      ps=20u
m07 vss    a1     w2     vss n w=12u  l=2.3636u ad=116p     pd=45u      as=36p      ps=18u
C0  vdd    a1     0.021f
C1  vss    a2     0.024f
C2  z      n3     0.213f
C3  vss    b1     0.029f
C4  n3     a1     0.029f
C5  z      a2     0.026f
C6  vdd    b2     0.025f
C7  w2     vss    0.004f
C8  n3     b2     0.089f
C9  a1     a2     0.207f
C10 z      b1     0.292f
C11 a2     b2     0.234f
C12 a1     b1     0.075f
C13 w2     a1     0.011f
C14 vss    z      0.196f
C15 b2     b1     0.187f
C16 vss    a1     0.071f
C17 vdd    n3     0.310f
C18 z      a1     0.070f
C19 vdd    a2     0.067f
C20 vss    b2     0.018f
C21 vdd    b1     0.016f
C22 n3     a2     0.121f
C23 z      b2     0.080f
C24 w1     vss    0.004f
C25 a1     b2     0.048f
C26 n3     b1     0.025f
C27 w1     z      0.013f
C28 a2     b1     0.052f
C29 vdd    z      0.045f
C30 vss    n3     0.003f
C33 z      vss    0.013f
C34 a1     vss    0.029f
C35 a2     vss    0.021f
C36 b2     vss    0.020f
C37 b1     vss    0.024f
.ends
