magic
tech scmos
timestamp 1179387596
<< checkpaint >>
rect -22 -25 102 105
<< ab >>
rect 0 0 80 80
<< pwell >>
rect -4 -7 84 36
<< nwell >>
rect -4 36 84 87
<< polysilicon >>
rect 19 70 21 74
rect 29 70 31 74
rect 36 70 38 74
rect 9 63 11 68
rect 69 58 71 63
rect 52 53 58 54
rect 52 49 53 53
rect 57 49 58 53
rect 9 44 11 47
rect 9 43 15 44
rect 9 39 10 43
rect 14 39 15 43
rect 9 38 15 39
rect 19 39 21 47
rect 19 38 25 39
rect 10 23 12 38
rect 19 34 20 38
rect 24 34 25 38
rect 29 38 31 47
rect 36 44 38 47
rect 52 44 58 49
rect 36 42 58 44
rect 29 37 48 38
rect 29 36 43 37
rect 19 33 25 34
rect 37 33 43 36
rect 47 33 48 37
rect 19 29 21 33
rect 17 26 21 29
rect 37 32 48 33
rect 56 35 58 42
rect 69 39 71 42
rect 65 38 71 39
rect 56 32 59 35
rect 65 34 66 38
rect 70 34 71 38
rect 65 33 71 34
rect 17 23 19 26
rect 27 23 29 28
rect 37 23 39 32
rect 57 29 59 32
rect 69 24 71 33
rect 57 18 59 22
rect 10 11 12 16
rect 17 11 19 16
rect 27 8 29 16
rect 37 12 39 16
rect 69 8 71 17
rect 27 6 71 8
<< ndiffusion >>
rect 50 27 57 29
rect 50 23 51 27
rect 55 23 57 27
rect 2 16 10 23
rect 12 16 17 23
rect 19 22 27 23
rect 19 18 21 22
rect 25 18 27 22
rect 19 16 27 18
rect 29 22 37 23
rect 29 18 31 22
rect 35 18 37 22
rect 29 16 37 18
rect 39 21 46 23
rect 50 22 57 23
rect 59 24 67 29
rect 59 22 69 24
rect 39 17 41 21
rect 45 17 46 21
rect 61 18 62 22
rect 66 18 69 22
rect 61 17 69 18
rect 71 23 78 24
rect 71 19 73 23
rect 77 19 78 23
rect 71 17 78 19
rect 39 16 46 17
rect 2 12 8 16
rect 2 8 3 12
rect 7 8 8 12
rect 2 7 8 8
<< pdiffusion >>
rect 61 72 67 73
rect 14 63 19 70
rect 2 62 9 63
rect 2 58 3 62
rect 7 58 9 62
rect 2 57 9 58
rect 4 47 9 57
rect 11 54 19 63
rect 11 50 13 54
rect 17 50 19 54
rect 11 47 19 50
rect 21 52 29 70
rect 21 48 23 52
rect 27 48 29 52
rect 21 47 29 48
rect 31 47 36 70
rect 38 69 47 70
rect 38 65 40 69
rect 44 65 47 69
rect 38 47 47 65
rect 61 68 62 72
rect 66 68 67 72
rect 61 58 67 68
rect 61 42 69 58
rect 71 55 76 58
rect 71 54 78 55
rect 71 50 73 54
rect 77 50 78 54
rect 71 47 78 50
rect 71 43 73 47
rect 77 43 78 47
rect 71 42 78 43
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect -2 72 82 78
rect -2 69 62 72
rect -2 68 40 69
rect 39 65 40 68
rect 44 68 62 69
rect 66 68 82 72
rect 44 65 45 68
rect 2 58 3 62
rect 7 58 77 62
rect 2 50 13 54
rect 17 50 18 54
rect 23 52 27 53
rect 2 22 6 50
rect 23 46 27 48
rect 10 43 27 46
rect 14 42 27 43
rect 10 30 14 39
rect 31 38 35 58
rect 19 34 20 38
rect 24 34 35 38
rect 42 39 46 55
rect 50 53 62 55
rect 50 49 53 53
rect 57 49 62 53
rect 58 41 62 49
rect 73 54 77 58
rect 73 47 77 50
rect 42 37 54 39
rect 42 33 43 37
rect 47 33 54 37
rect 66 38 70 47
rect 66 31 70 34
rect 10 29 35 30
rect 10 27 55 29
rect 10 26 51 27
rect 31 25 51 26
rect 31 22 35 25
rect 58 25 70 31
rect 51 22 55 23
rect 73 23 77 43
rect 2 18 21 22
rect 25 18 26 22
rect 31 17 35 18
rect 40 17 41 21
rect 45 17 46 21
rect 40 12 46 17
rect 61 18 62 22
rect 66 18 67 22
rect 73 18 77 19
rect 51 12 55 16
rect 61 12 67 18
rect -2 8 3 12
rect 7 8 82 12
rect -2 2 82 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
<< ntransistor >>
rect 10 16 12 23
rect 17 16 19 23
rect 27 16 29 23
rect 37 16 39 23
rect 57 22 59 29
rect 69 17 71 24
<< ptransistor >>
rect 9 47 11 63
rect 19 47 21 70
rect 29 47 31 70
rect 36 47 38 70
rect 69 42 71 58
<< polycontact >>
rect 53 49 57 53
rect 10 39 14 43
rect 20 34 24 38
rect 43 33 47 37
rect 66 34 70 38
<< ndcontact >>
rect 51 23 55 27
rect 21 18 25 22
rect 31 18 35 22
rect 41 17 45 21
rect 62 18 66 22
rect 73 19 77 23
rect 3 8 7 12
<< pdcontact >>
rect 3 58 7 62
rect 13 50 17 54
rect 23 48 27 52
rect 40 65 44 69
rect 62 68 66 72
rect 73 50 77 54
rect 73 43 77 47
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
<< psubstratepdiff >>
rect 0 2 80 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 80 2
rect 0 -3 80 -2
<< nsubstratendiff >>
rect 0 82 80 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 80 82
rect 0 77 80 78
<< labels >>
rlabel polycontact 12 41 12 41 6 an
rlabel polycontact 22 36 22 36 6 bn
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 20 12 20 6 z
rlabel metal1 20 20 20 20 6 z
rlabel metal1 12 36 12 36 6 an
rlabel metal1 25 47 25 47 6 an
rlabel metal1 12 52 12 52 6 z
rlabel metal1 40 6 40 6 6 vss
rlabel metal1 33 23 33 23 6 an
rlabel metal1 27 36 27 36 6 bn
rlabel metal1 44 44 44 44 6 a2
rlabel metal1 40 74 40 74 6 vdd
rlabel ndcontact 53 25 53 25 6 an
rlabel metal1 60 28 60 28 6 b
rlabel metal1 52 36 52 36 6 a2
rlabel metal1 60 48 60 48 6 a1
rlabel metal1 52 52 52 52 6 a1
rlabel polycontact 68 36 68 36 6 b
rlabel metal1 75 40 75 40 6 bn
rlabel metal1 39 60 39 60 6 bn
<< end >>
