.subckt nd3v0x3 a b c vdd vss z
*   SPICE3 file   created from nd3v0x3.ext -      technology: scmos
m00 z      a      vdd    vdd p w=20u  l=2.3636u ad=80p      pd=28u      as=100p     ps=36.6667u
m01 vdd    b      z      vdd p w=20u  l=2.3636u ad=100p     pd=36.6667u as=80p      ps=28u
m02 z      c      vdd    vdd p w=20u  l=2.3636u ad=80p      pd=28u      as=100p     ps=36.6667u
m03 vdd    c      z      vdd p w=20u  l=2.3636u ad=100p     pd=36.6667u as=80p      ps=28u
m04 z      b      vdd    vdd p w=20u  l=2.3636u ad=80p      pd=28u      as=100p     ps=36.6667u
m05 vdd    a      z      vdd p w=20u  l=2.3636u ad=100p     pd=36.6667u as=80p      ps=28u
m06 w1     a      vss    vss n w=20u  l=2.3636u ad=50p      pd=25u      as=149.5p   ps=56u
m07 w2     b      w1     vss n w=20u  l=2.3636u ad=50p      pd=25u      as=50p      ps=25u
m08 z      c      w2     vss n w=20u  l=2.3636u ad=80p      pd=28u      as=50p      ps=25u
m09 w3     c      z      vss n w=20u  l=2.3636u ad=50p      pd=25u      as=80p      ps=28u
m10 w4     b      w3     vss n w=20u  l=2.3636u ad=50p      pd=25u      as=50p      ps=25u
m11 vss    a      w4     vss n w=20u  l=2.3636u ad=149.5p   pd=56u      as=50p      ps=25u
C0  w3     vss    0.005f
C1  b      vdd    0.083f
C2  w1     vss    0.005f
C3  w2     z      0.010f
C4  vss    z      0.279f
C5  w3     a      0.018f
C6  z      c      0.086f
C7  vss    b      0.044f
C8  w1     a      0.007f
C9  z      a      0.457f
C10 c      b      0.355f
C11 vss    vdd    0.005f
C12 w4     vss    0.005f
C13 b      a      0.339f
C14 c      vdd    0.023f
C15 w2     vss    0.005f
C16 a      vdd    0.058f
C17 w1     z      0.010f
C18 w4     a      0.003f
C19 vss    c      0.027f
C20 w2     a      0.007f
C21 z      b      0.329f
C22 vss    a      0.207f
C23 c      a      0.243f
C24 z      vdd    0.522f
C26 z      vss    0.016f
C27 c      vss    0.036f
C28 b      vss    0.046f
C29 a      vss    0.043f
.ends
