.subckt oai211v0x05 a1 a2 b c vdd vss z
*   SPICE3 file   created from oai211v0x05.ext -      technology: scmos
m00 z      c      vdd    vdd p w=9u   l=2.3636u ad=43.4118p pd=21.1765u as=76.7647p ps=31.7647u
m01 vdd    b      z      vdd p w=9u   l=2.3636u ad=76.7647p pd=31.7647u as=43.4118p ps=21.1765u
m02 w1     a1     vdd    vdd p w=16u  l=2.3636u ad=40p      pd=21u      as=136.471p ps=56.4706u
m03 z      a2     w1     vdd p w=16u  l=2.3636u ad=77.1765p pd=37.6471u as=40p      ps=21u
m04 w2     c      z      vss n w=10u  l=2.3636u ad=25p      pd=15u      as=62p      ps=34u
m05 n1     b      w2     vss n w=10u  l=2.3636u ad=47.3333p pd=23.3333u as=25p      ps=15u
m06 vss    a1     n1     vss n w=10u  l=2.3636u ad=78p      pd=32u      as=47.3333p ps=23.3333u
m07 n1     a2     vss    vss n w=10u  l=2.3636u ad=47.3333p pd=23.3333u as=78p      ps=32u
C0  vss    a2     0.011f
C1  n1     vdd    0.003f
C2  z      b      0.142f
C3  b      c      0.163f
C4  z      a2     0.116f
C5  n1     vss    0.173f
C6  b      a1     0.110f
C7  c      a2     0.081f
C8  z      vdd    0.301f
C9  n1     z      0.035f
C10 a2     a1     0.125f
C11 c      vdd    0.038f
C12 n1     c      0.016f
C13 vss    z      0.030f
C14 w2     b      0.009f
C15 a1     vdd    0.016f
C16 vss    c      0.024f
C17 n1     a1     0.056f
C18 z      c      0.142f
C19 w1     a2     0.005f
C20 vss    a1     0.031f
C21 w1     vdd    0.003f
C22 b      a2     0.025f
C23 z      a1     0.041f
C24 c      a1     0.079f
C25 b      vdd    0.010f
C26 n1     b      0.052f
C27 a2     vdd    0.031f
C28 w1     z      0.010f
C29 n1     a2     0.020f
C30 vss    b      0.046f
C31 n1     vss    0.002f
C33 z      vss    0.017f
C34 b      vss    0.026f
C35 c      vss    0.031f
C36 a2     vss    0.028f
C37 a1     vss    0.028f
.ends
