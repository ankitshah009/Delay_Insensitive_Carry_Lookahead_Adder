magic
tech scmos
timestamp 1179385751
<< checkpaint >>
rect -22 -25 190 105
<< ab >>
rect 0 0 168 80
<< pwell >>
rect -4 -7 172 36
<< nwell >>
rect -4 36 172 87
<< polysilicon >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 39 70 41 74
rect 49 70 51 74
rect 59 70 61 74
rect 69 70 71 74
rect 76 70 78 74
rect 89 70 91 74
rect 96 70 98 74
rect 106 70 108 74
rect 113 70 115 74
rect 125 70 127 74
rect 135 70 137 74
rect 145 70 147 74
rect 9 37 11 42
rect 19 37 21 42
rect 29 37 31 42
rect 9 35 31 37
rect 9 30 11 35
rect 19 30 21 35
rect 29 30 31 35
rect 39 39 41 42
rect 49 39 51 42
rect 59 39 61 42
rect 69 39 71 42
rect 76 39 78 42
rect 89 39 91 42
rect 39 38 61 39
rect 39 37 56 38
rect 39 30 41 37
rect 49 34 56 37
rect 60 34 61 38
rect 49 33 61 34
rect 66 38 72 39
rect 66 34 67 38
rect 71 34 72 38
rect 66 33 72 34
rect 76 38 91 39
rect 76 34 82 38
rect 86 34 91 38
rect 76 33 91 34
rect 49 30 51 33
rect 59 30 61 33
rect 69 30 71 33
rect 76 30 78 33
rect 89 30 91 33
rect 96 39 98 42
rect 106 39 108 42
rect 96 38 108 39
rect 96 34 97 38
rect 101 34 108 38
rect 96 33 108 34
rect 96 30 98 33
rect 106 30 108 33
rect 113 39 115 42
rect 125 39 127 42
rect 135 39 137 42
rect 145 39 147 42
rect 113 38 147 39
rect 113 34 114 38
rect 118 37 147 38
rect 118 34 128 37
rect 113 33 128 34
rect 113 30 115 33
rect 126 30 128 33
rect 136 30 138 37
rect 9 11 11 16
rect 19 11 21 16
rect 29 8 31 16
rect 39 12 41 16
rect 49 12 51 16
rect 59 12 61 16
rect 69 8 71 16
rect 76 11 78 16
rect 29 6 71 8
rect 89 11 91 16
rect 96 11 98 16
rect 106 11 108 16
rect 113 11 115 16
rect 126 6 128 10
rect 136 6 138 10
<< ndiffusion >>
rect 2 28 9 30
rect 2 24 3 28
rect 7 24 9 28
rect 2 21 9 24
rect 2 17 3 21
rect 7 17 9 21
rect 2 16 9 17
rect 11 29 19 30
rect 11 25 13 29
rect 17 25 19 29
rect 11 22 19 25
rect 11 18 13 22
rect 17 18 19 22
rect 11 16 19 18
rect 21 21 29 30
rect 21 17 23 21
rect 27 17 29 21
rect 21 16 29 17
rect 31 29 39 30
rect 31 25 33 29
rect 37 25 39 29
rect 31 22 39 25
rect 31 18 33 22
rect 37 18 39 22
rect 31 16 39 18
rect 41 29 49 30
rect 41 25 43 29
rect 47 25 49 29
rect 41 16 49 25
rect 51 22 59 30
rect 51 18 53 22
rect 57 18 59 22
rect 51 16 59 18
rect 61 29 69 30
rect 61 25 63 29
rect 67 25 69 29
rect 61 16 69 25
rect 71 16 76 30
rect 78 16 89 30
rect 91 16 96 30
rect 98 29 106 30
rect 98 25 100 29
rect 104 25 106 29
rect 98 16 106 25
rect 108 16 113 30
rect 115 16 126 30
rect 80 12 87 16
rect 80 8 81 12
rect 85 8 87 12
rect 117 15 126 16
rect 117 11 118 15
rect 122 11 126 15
rect 117 10 126 11
rect 128 29 136 30
rect 128 25 130 29
rect 134 25 136 29
rect 128 22 136 25
rect 128 18 130 22
rect 134 18 136 22
rect 128 10 136 18
rect 138 23 146 30
rect 138 19 140 23
rect 144 19 146 23
rect 138 15 146 19
rect 138 11 140 15
rect 144 11 146 15
rect 138 10 146 11
rect 80 7 87 8
<< pdiffusion >>
rect 2 69 9 70
rect 2 65 3 69
rect 7 65 9 69
rect 2 62 9 65
rect 2 58 3 62
rect 7 58 9 62
rect 2 55 9 58
rect 2 51 3 55
rect 7 51 9 55
rect 2 42 9 51
rect 11 62 19 70
rect 11 58 13 62
rect 17 58 19 62
rect 11 55 19 58
rect 11 51 13 55
rect 17 51 19 55
rect 11 42 19 51
rect 21 69 29 70
rect 21 65 23 69
rect 27 65 29 69
rect 21 62 29 65
rect 21 58 23 62
rect 27 58 29 62
rect 21 42 29 58
rect 31 62 39 70
rect 31 58 33 62
rect 37 58 39 62
rect 31 55 39 58
rect 31 51 33 55
rect 37 51 39 55
rect 31 42 39 51
rect 41 54 49 70
rect 41 50 43 54
rect 47 50 49 54
rect 41 42 49 50
rect 51 62 59 70
rect 51 58 53 62
rect 57 58 59 62
rect 51 42 59 58
rect 61 54 69 70
rect 61 50 63 54
rect 67 50 69 54
rect 61 42 69 50
rect 71 42 76 70
rect 78 69 89 70
rect 78 65 81 69
rect 85 65 89 69
rect 78 42 89 65
rect 91 42 96 70
rect 98 54 106 70
rect 98 50 100 54
rect 104 50 106 54
rect 98 42 106 50
rect 108 42 113 70
rect 115 69 125 70
rect 115 65 118 69
rect 122 65 125 69
rect 115 42 125 65
rect 127 62 135 70
rect 127 58 129 62
rect 133 58 135 62
rect 127 55 135 58
rect 127 51 129 55
rect 133 51 135 55
rect 127 42 135 51
rect 137 69 145 70
rect 137 65 139 69
rect 143 65 145 69
rect 137 62 145 65
rect 137 58 139 62
rect 143 58 145 62
rect 137 42 145 58
rect 147 55 152 70
rect 147 54 154 55
rect 147 50 149 54
rect 153 50 154 54
rect 147 47 154 50
rect 147 43 149 47
rect 153 43 154 47
rect 147 42 154 43
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect 118 78 122 82
rect 126 78 130 82
rect 134 78 138 82
rect 142 78 146 82
rect 150 78 154 82
rect 158 78 162 82
rect 166 78 170 82
rect -2 69 170 78
rect -2 68 3 69
rect 7 68 23 69
rect 3 62 7 65
rect 22 65 23 68
rect 27 68 81 69
rect 27 65 28 68
rect 80 65 81 68
rect 85 68 118 69
rect 85 65 86 68
rect 117 65 118 68
rect 122 68 139 69
rect 122 65 123 68
rect 138 65 139 68
rect 143 68 170 69
rect 143 65 144 68
rect 3 55 7 58
rect 3 50 7 51
rect 13 62 17 63
rect 22 62 28 65
rect 138 62 144 65
rect 22 58 23 62
rect 27 58 28 62
rect 32 58 33 62
rect 37 58 53 62
rect 57 58 129 62
rect 133 58 134 62
rect 138 58 139 62
rect 143 58 144 62
rect 157 59 161 68
rect 13 55 17 58
rect 32 55 37 58
rect 32 54 33 55
rect 17 51 33 54
rect 129 55 134 58
rect 13 50 37 51
rect 42 50 43 54
rect 47 50 63 54
rect 67 50 100 54
rect 104 50 126 54
rect 133 54 134 55
rect 133 51 149 54
rect 129 50 149 51
rect 153 50 154 54
rect 13 29 37 30
rect 3 28 7 29
rect 3 21 7 24
rect 17 26 33 29
rect 13 22 17 25
rect 32 25 33 26
rect 42 29 46 50
rect 57 39 63 46
rect 81 42 118 46
rect 50 38 63 39
rect 50 34 56 38
rect 60 34 63 38
rect 50 33 63 34
rect 67 38 77 39
rect 71 34 77 38
rect 81 38 87 42
rect 114 38 118 42
rect 81 34 82 38
rect 86 34 87 38
rect 91 34 97 38
rect 101 34 103 38
rect 67 33 77 34
rect 73 30 77 33
rect 91 30 95 34
rect 114 33 118 34
rect 42 25 43 29
rect 47 25 63 29
rect 67 25 68 29
rect 73 26 95 30
rect 122 29 126 50
rect 148 47 154 50
rect 148 43 149 47
rect 153 43 154 47
rect 99 25 100 29
rect 104 25 126 29
rect 130 29 135 30
rect 134 25 135 29
rect 32 22 37 25
rect 130 22 135 25
rect 13 17 17 18
rect 23 21 27 22
rect 32 18 33 22
rect 37 18 53 22
rect 57 18 130 22
rect 134 18 135 22
rect 140 23 144 24
rect 3 12 7 17
rect 23 12 27 17
rect 140 15 144 19
rect 117 12 118 15
rect -2 8 81 12
rect 85 11 118 12
rect 122 12 123 15
rect 122 11 140 12
rect 154 12 158 21
rect 144 11 170 12
rect 85 8 170 11
rect -2 2 170 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 122 2
rect 126 -2 130 2
rect 134 -2 138 2
rect 142 -2 146 2
rect 150 -2 154 2
rect 158 -2 162 2
rect 166 -2 170 2
<< ntransistor >>
rect 9 16 11 30
rect 19 16 21 30
rect 29 16 31 30
rect 39 16 41 30
rect 49 16 51 30
rect 59 16 61 30
rect 69 16 71 30
rect 76 16 78 30
rect 89 16 91 30
rect 96 16 98 30
rect 106 16 108 30
rect 113 16 115 30
rect 126 10 128 30
rect 136 10 138 30
<< ptransistor >>
rect 9 42 11 70
rect 19 42 21 70
rect 29 42 31 70
rect 39 42 41 70
rect 49 42 51 70
rect 59 42 61 70
rect 69 42 71 70
rect 76 42 78 70
rect 89 42 91 70
rect 96 42 98 70
rect 106 42 108 70
rect 113 42 115 70
rect 125 42 127 70
rect 135 42 137 70
rect 145 42 147 70
<< polycontact >>
rect 56 34 60 38
rect 67 34 71 38
rect 82 34 86 38
rect 97 34 101 38
rect 114 34 118 38
<< ndcontact >>
rect 3 24 7 28
rect 3 17 7 21
rect 13 25 17 29
rect 13 18 17 22
rect 23 17 27 21
rect 33 25 37 29
rect 33 18 37 22
rect 43 25 47 29
rect 53 18 57 22
rect 63 25 67 29
rect 100 25 104 29
rect 81 8 85 12
rect 118 11 122 15
rect 130 25 134 29
rect 130 18 134 22
rect 140 19 144 23
rect 140 11 144 15
<< pdcontact >>
rect 3 65 7 69
rect 3 58 7 62
rect 3 51 7 55
rect 13 58 17 62
rect 13 51 17 55
rect 23 65 27 69
rect 23 58 27 62
rect 33 58 37 62
rect 33 51 37 55
rect 43 50 47 54
rect 53 58 57 62
rect 63 50 67 54
rect 81 65 85 69
rect 100 50 104 54
rect 118 65 122 69
rect 129 58 133 62
rect 129 51 133 55
rect 139 65 143 69
rect 139 58 143 62
rect 149 50 153 54
rect 149 43 153 47
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
rect 90 -2 94 2
rect 98 -2 102 2
rect 106 -2 110 2
rect 114 -2 118 2
rect 122 -2 126 2
rect 130 -2 134 2
rect 138 -2 142 2
rect 146 -2 150 2
rect 154 -2 158 2
rect 162 -2 166 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
rect 90 78 94 82
rect 98 78 102 82
rect 106 78 110 82
rect 114 78 118 82
rect 122 78 126 82
rect 130 78 134 82
rect 138 78 142 82
rect 146 78 150 82
rect 154 78 158 82
rect 162 78 166 82
<< psubstratepdiff >>
rect 0 2 168 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 122 2
rect 126 -2 130 2
rect 134 -2 138 2
rect 142 -2 146 2
rect 150 -2 154 2
rect 158 -2 162 2
rect 166 -2 168 2
rect 0 -3 168 -2
<< nsubstratendiff >>
rect 0 82 168 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect 118 78 122 82
rect 126 78 130 82
rect 134 78 138 82
rect 142 78 146 82
rect 150 78 154 82
rect 158 78 162 82
rect 166 78 168 82
rect 0 77 168 78
<< labels >>
rlabel metal1 15 23 15 23 6 n3
rlabel metal1 15 56 15 56 6 n1
rlabel metal1 34 24 34 24 6 n3
rlabel metal1 52 36 52 36 6 c
rlabel metal1 60 40 60 40 6 c
rlabel metal1 44 36 44 36 6 z
rlabel metal1 52 52 52 52 6 z
rlabel metal1 60 52 60 52 6 z
rlabel metal1 34 56 34 56 6 n1
rlabel metal1 84 6 84 6 6 vss
rlabel metal1 76 28 76 28 6 b
rlabel metal1 84 28 84 28 6 b
rlabel metal1 92 28 92 28 6 b
rlabel metal1 84 40 84 40 6 a
rlabel metal1 92 44 92 44 6 a
rlabel metal1 76 52 76 52 6 z
rlabel metal1 84 52 84 52 6 z
rlabel metal1 92 52 92 52 6 z
rlabel metal1 68 52 68 52 6 z
rlabel metal1 84 74 84 74 6 vdd
rlabel polycontact 100 36 100 36 6 b
rlabel metal1 100 44 100 44 6 a
rlabel metal1 108 44 108 44 6 a
rlabel polycontact 116 36 116 36 6 a
rlabel metal1 124 36 124 36 6 z
rlabel metal1 108 52 108 52 6 z
rlabel metal1 116 52 116 52 6 z
rlabel metal1 131 56 131 56 6 n1
rlabel metal1 100 52 100 52 6 z
rlabel metal1 83 60 83 60 6 n1
rlabel metal1 132 24 132 24 6 n3
rlabel metal1 83 20 83 20 6 n3
rlabel metal1 151 48 151 48 6 n1
rlabel metal1 141 52 141 52 6 n1
<< end >>
