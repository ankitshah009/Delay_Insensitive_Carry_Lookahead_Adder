.subckt nr3v0x3 a b c vdd vss z
*   SPICE3 file   created from nr3v0x3.ext -      technology: scmos
m00 w1     a      vdd    vdd p w=28u  l=2.3636u ad=84p      pd=34u      as=157.942p ps=53.2816u
m01 w2     b      w1     vdd p w=28u  l=2.3636u ad=84p      pd=34u      as=84p      ps=34u
m02 z      c      w2     vdd p w=28u  l=2.3636u ad=114.447p pd=39.1456u as=84p      ps=34u
m03 w3     c      z      vdd p w=28u  l=2.3636u ad=70p      pd=33u      as=114.447p ps=39.1456u
m04 w4     b      w3     vdd p w=28u  l=2.3636u ad=70p      pd=33u      as=70p      ps=33u
m05 vdd    a      w4     vdd p w=28u  l=2.3636u ad=157.942p pd=53.2816u as=70p      ps=33u
m06 w5     a      vdd    vdd p w=28u  l=2.3636u ad=70p      pd=33u      as=157.942p ps=53.2816u
m07 w6     b      w5     vdd p w=28u  l=2.3636u ad=70p      pd=33u      as=70p      ps=33u
m08 z      c      w6     vdd p w=28u  l=2.3636u ad=114.447p pd=39.1456u as=70p      ps=33u
m09 w7     c      z      vdd p w=19u  l=2.3636u ad=47.5p    pd=24u      as=77.6602p ps=26.5631u
m10 w8     b      w7     vdd p w=19u  l=2.3636u ad=47.5p    pd=24u      as=47.5p    ps=24u
m11 vdd    a      w8     vdd p w=19u  l=2.3636u ad=107.175p pd=36.1553u as=47.5p    ps=24u
m12 vss    a      z      vss n w=19u  l=2.3636u ad=122p     pd=40u      as=91p      ps=35.3333u
m13 z      b      vss    vss n w=19u  l=2.3636u ad=91p      pd=35.3333u as=122p     ps=40u
m14 vss    c      z      vss n w=19u  l=2.3636u ad=122p     pd=40u      as=91p      ps=35.3333u
C0  vdd    c      0.059f
C1  w2     a      0.009f
C2  w4     z      0.010f
C3  vss    b      0.416f
C4  c      b      0.741f
C5  vdd    a      0.162f
C6  w5     vdd    0.005f
C7  b      a      0.518f
C8  w3     vdd    0.005f
C9  z      w1     0.012f
C10 vss    z      0.293f
C11 w2     vdd    0.006f
C12 w4     a      0.007f
C13 z      c      0.145f
C14 w7     z      0.007f
C15 z      a      0.728f
C16 w5     z      0.010f
C17 vss    c      0.109f
C18 vdd    b      0.041f
C19 w1     a      0.009f
C20 vss    a      0.124f
C21 w6     vdd    0.005f
C22 w3     z      0.010f
C23 c      a      0.552f
C24 z      w2     0.012f
C25 w4     vdd    0.005f
C26 z      vdd    0.359f
C27 w3     a      0.007f
C28 w1     vdd    0.006f
C29 z      b      0.248f
C30 w6     z      0.010f
C31 vss    vdd    0.005f
C33 z      vss    0.010f
C35 c      vss    0.072f
C36 b      vss    0.092f
C37 a      vss    0.055f
.ends
