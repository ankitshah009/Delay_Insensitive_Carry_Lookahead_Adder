magic
tech scmos
timestamp 1179385370
<< checkpaint >>
rect -22 -22 118 94
<< ab >>
rect 0 0 96 72
<< pwell >>
rect -4 -4 100 32
<< nwell >>
rect -4 32 100 76
<< polysilicon >>
rect 9 66 11 70
rect 19 66 21 70
rect 29 66 31 70
rect 39 66 41 70
rect 49 66 51 70
rect 59 66 61 70
rect 69 66 71 70
rect 79 66 81 70
rect 9 35 11 38
rect 19 35 21 38
rect 29 35 31 38
rect 9 34 21 35
rect 9 30 10 34
rect 14 30 21 34
rect 9 29 21 30
rect 25 34 31 35
rect 25 30 26 34
rect 30 31 31 34
rect 39 35 41 38
rect 49 35 51 38
rect 59 35 61 38
rect 69 35 71 38
rect 79 35 81 38
rect 39 34 45 35
rect 30 30 35 31
rect 25 29 35 30
rect 39 30 40 34
rect 44 30 45 34
rect 39 29 45 30
rect 49 34 63 35
rect 49 30 50 34
rect 54 30 58 34
rect 62 30 63 34
rect 49 29 63 30
rect 67 34 73 35
rect 67 30 68 34
rect 72 30 73 34
rect 67 29 73 30
rect 77 34 88 35
rect 77 30 83 34
rect 87 30 88 34
rect 77 29 88 30
rect 9 26 11 29
rect 19 26 21 29
rect 33 26 35 29
rect 41 26 43 29
rect 49 26 51 29
rect 61 26 63 29
rect 69 26 71 29
rect 77 26 79 29
rect 9 13 11 18
rect 19 13 21 18
rect 33 3 35 8
rect 41 3 43 8
rect 49 3 51 8
rect 61 3 63 8
rect 69 3 71 8
rect 77 3 79 8
<< ndiffusion >>
rect 2 23 9 26
rect 2 19 3 23
rect 7 19 9 23
rect 2 18 9 19
rect 11 25 19 26
rect 11 21 13 25
rect 17 21 19 25
rect 11 18 19 21
rect 21 18 33 26
rect 23 8 33 18
rect 35 8 41 26
rect 43 8 49 26
rect 51 18 61 26
rect 51 14 54 18
rect 58 14 61 18
rect 51 8 61 14
rect 63 8 69 26
rect 71 8 77 26
rect 79 13 87 26
rect 79 9 81 13
rect 85 9 87 13
rect 79 8 87 9
rect 23 4 25 8
rect 29 4 31 8
rect 23 3 31 4
<< pdiffusion >>
rect 4 60 9 66
rect 2 59 9 60
rect 2 55 3 59
rect 7 55 9 59
rect 2 54 9 55
rect 4 38 9 54
rect 11 50 19 66
rect 11 46 13 50
rect 17 46 19 50
rect 11 43 19 46
rect 11 39 13 43
rect 17 39 19 43
rect 11 38 19 39
rect 21 58 29 66
rect 21 54 23 58
rect 27 54 29 58
rect 21 51 29 54
rect 21 47 23 51
rect 27 47 29 51
rect 21 38 29 47
rect 31 65 39 66
rect 31 61 33 65
rect 37 61 39 65
rect 31 38 39 61
rect 41 58 49 66
rect 41 54 43 58
rect 47 54 49 58
rect 41 51 49 54
rect 41 47 43 51
rect 47 47 49 51
rect 41 38 49 47
rect 51 65 59 66
rect 51 61 53 65
rect 57 61 59 65
rect 51 58 59 61
rect 51 54 53 58
rect 57 54 59 58
rect 51 38 59 54
rect 61 57 69 66
rect 61 53 63 57
rect 67 53 69 57
rect 61 50 69 53
rect 61 46 63 50
rect 67 46 69 50
rect 61 38 69 46
rect 71 65 79 66
rect 71 61 73 65
rect 77 61 79 65
rect 71 58 79 61
rect 71 54 73 58
rect 77 54 79 58
rect 71 38 79 54
rect 81 51 86 66
rect 81 50 88 51
rect 81 46 83 50
rect 87 46 88 50
rect 81 43 88 46
rect 81 39 83 43
rect 87 39 88 43
rect 81 38 88 39
<< metal1 >>
rect -2 65 98 72
rect -2 64 33 65
rect 37 64 53 65
rect 33 60 37 61
rect 52 61 53 64
rect 57 64 73 65
rect 57 61 58 64
rect 2 55 3 59
rect 7 58 27 59
rect 7 55 23 58
rect 23 51 27 54
rect 2 35 6 51
rect 12 46 13 50
rect 17 46 18 50
rect 43 58 47 59
rect 52 58 58 61
rect 72 61 73 64
rect 77 64 98 65
rect 77 61 78 64
rect 72 58 78 61
rect 52 54 53 58
rect 57 54 58 58
rect 63 57 67 58
rect 43 51 47 54
rect 27 47 43 50
rect 72 54 73 58
rect 77 54 78 58
rect 63 50 67 53
rect 47 47 63 50
rect 23 46 63 47
rect 67 46 83 50
rect 87 46 88 50
rect 12 43 18 46
rect 82 43 88 46
rect 12 39 13 43
rect 17 39 22 43
rect 2 34 14 35
rect 2 30 10 34
rect 2 29 14 30
rect 18 25 22 39
rect 39 38 73 42
rect 82 39 83 43
rect 87 39 88 43
rect 3 23 7 24
rect 12 21 13 25
rect 17 21 22 25
rect 26 34 30 35
rect 39 34 45 38
rect 67 34 73 38
rect 83 34 87 35
rect 39 30 40 34
rect 44 30 45 34
rect 49 30 50 34
rect 54 30 58 34
rect 62 30 63 34
rect 67 30 68 34
rect 72 30 79 34
rect 26 26 30 30
rect 83 26 87 30
rect 26 22 87 26
rect 3 8 7 19
rect 18 18 22 21
rect 18 14 54 18
rect 58 14 59 18
rect 66 13 70 22
rect 81 13 85 14
rect 81 8 85 9
rect -2 4 4 8
rect 8 4 12 8
rect 16 4 25 8
rect 29 4 98 8
rect -2 0 98 4
<< ntransistor >>
rect 9 18 11 26
rect 19 18 21 26
rect 33 8 35 26
rect 41 8 43 26
rect 49 8 51 26
rect 61 8 63 26
rect 69 8 71 26
rect 77 8 79 26
<< ptransistor >>
rect 9 38 11 66
rect 19 38 21 66
rect 29 38 31 66
rect 39 38 41 66
rect 49 38 51 66
rect 59 38 61 66
rect 69 38 71 66
rect 79 38 81 66
<< polycontact >>
rect 10 30 14 34
rect 26 30 30 34
rect 40 30 44 34
rect 50 30 54 34
rect 58 30 62 34
rect 68 30 72 34
rect 83 30 87 34
<< ndcontact >>
rect 3 19 7 23
rect 13 21 17 25
rect 54 14 58 18
rect 81 9 85 13
rect 25 4 29 8
<< pdcontact >>
rect 3 55 7 59
rect 13 46 17 50
rect 13 39 17 43
rect 23 54 27 58
rect 23 47 27 51
rect 33 61 37 65
rect 43 54 47 58
rect 43 47 47 51
rect 53 61 57 65
rect 53 54 57 58
rect 63 53 67 57
rect 63 46 67 50
rect 73 61 77 65
rect 73 54 77 58
rect 83 46 87 50
rect 83 39 87 43
<< psubstratepcontact >>
rect 4 4 8 8
rect 12 4 16 8
<< psubstratepdiff >>
rect 3 8 17 9
rect 3 4 4 8
rect 8 4 12 8
rect 16 4 17 8
rect 3 3 17 4
<< labels >>
rlabel polycontact 12 32 12 32 6 b
rlabel metal1 4 40 4 40 6 b
rlabel metal1 28 16 28 16 6 z
rlabel polycontact 28 32 28 32 6 a1
rlabel metal1 20 32 20 32 6 z
rlabel metal1 25 52 25 52 6 n3
rlabel metal1 14 57 14 57 6 n3
rlabel metal1 48 4 48 4 6 vss
rlabel metal1 44 16 44 16 6 z
rlabel metal1 52 16 52 16 6 z
rlabel metal1 36 16 36 16 6 z
rlabel metal1 36 24 36 24 6 a1
rlabel metal1 44 24 44 24 6 a1
rlabel metal1 52 24 52 24 6 a1
rlabel polycontact 52 32 52 32 6 a3
rlabel metal1 44 40 44 40 6 a2
rlabel metal1 52 40 52 40 6 a2
rlabel metal1 45 52 45 52 6 n3
rlabel metal1 48 68 48 68 6 vdd
rlabel metal1 60 24 60 24 6 a1
rlabel metal1 76 24 76 24 6 a1
rlabel metal1 68 20 68 20 6 a1
rlabel metal1 76 32 76 32 6 a2
rlabel polycontact 60 32 60 32 6 a3
rlabel metal1 60 40 60 40 6 a2
rlabel metal1 68 40 68 40 6 a2
rlabel metal1 65 52 65 52 6 n3
rlabel metal1 84 24 84 24 6 a1
rlabel metal1 85 44 85 44 6 n3
rlabel metal1 55 48 55 48 6 n3
<< end >>
