magic
tech scmos
timestamp 1185094768
<< checkpaint >>
rect -22 -22 62 122
<< ab >>
rect 0 0 40 100
<< pwell >>
rect -4 -4 44 48
<< nwell >>
rect -4 48 44 104
<< polysilicon >>
rect 15 94 17 98
rect 23 94 25 98
rect 15 43 17 55
rect 23 52 25 55
rect 23 51 33 52
rect 23 49 28 51
rect 25 47 28 49
rect 32 47 33 51
rect 25 46 33 47
rect 13 42 21 43
rect 13 38 16 42
rect 20 38 21 42
rect 13 37 21 38
rect 13 28 15 37
rect 25 28 27 46
rect 13 12 15 17
rect 25 12 27 17
<< ndiffusion >>
rect 4 22 13 28
rect 4 18 6 22
rect 10 18 13 22
rect 4 17 13 18
rect 15 27 25 28
rect 15 23 18 27
rect 22 23 25 27
rect 15 17 25 23
rect 27 22 36 28
rect 27 18 30 22
rect 34 18 36 22
rect 27 17 36 18
<< pdiffusion >>
rect 10 69 15 94
rect 7 68 15 69
rect 7 64 8 68
rect 12 64 15 68
rect 7 60 15 64
rect 7 56 8 60
rect 12 56 15 60
rect 7 55 15 56
rect 17 55 23 94
rect 25 92 34 94
rect 25 88 28 92
rect 32 88 34 92
rect 25 82 34 88
rect 25 78 28 82
rect 32 78 34 82
rect 25 55 34 78
<< metal1 >>
rect -2 92 42 100
rect -2 88 28 92
rect 32 88 42 92
rect 28 82 32 88
rect 28 77 32 78
rect 8 68 12 73
rect 8 60 12 64
rect 27 62 33 72
rect 17 58 33 62
rect 8 33 12 56
rect 18 43 22 53
rect 27 51 33 58
rect 27 47 28 51
rect 32 47 33 51
rect 16 42 32 43
rect 20 38 32 42
rect 16 37 32 38
rect 8 27 22 33
rect 6 22 10 23
rect 6 12 10 18
rect 18 17 22 23
rect 30 22 34 23
rect 30 12 34 18
rect -2 8 42 12
rect -2 4 8 8
rect 12 4 18 8
rect 22 4 42 8
rect -2 0 42 4
<< ntransistor >>
rect 13 17 15 28
rect 25 17 27 28
<< ptransistor >>
rect 15 55 17 94
rect 23 55 25 94
<< polycontact >>
rect 28 47 32 51
rect 16 38 20 42
<< ndcontact >>
rect 6 18 10 22
rect 18 23 22 27
rect 30 18 34 22
<< pdcontact >>
rect 8 64 12 68
rect 8 56 12 60
rect 28 88 32 92
rect 28 78 32 82
<< psubstratepcontact >>
rect 8 4 12 8
rect 18 4 22 8
<< psubstratepdiff >>
rect 7 8 23 9
rect 7 4 8 8
rect 12 4 18 8
rect 22 4 23 8
rect 7 3 23 4
<< labels >>
rlabel metal1 10 50 10 50 6 z
rlabel psubstratepcontact 20 6 20 6 6 vss
rlabel ndcontact 20 25 20 25 6 z
rlabel metal1 20 45 20 45 6 b
rlabel metal1 20 60 20 60 6 a
rlabel metal1 20 94 20 94 6 vdd
rlabel metal1 30 40 30 40 6 b
rlabel metal1 30 60 30 60 6 a
<< end >>
