magic
tech scmos
timestamp 1179387117
<< checkpaint >>
rect -22 -25 94 105
<< ab >>
rect 0 0 72 80
<< pwell >>
rect -4 -7 76 36
<< nwell >>
rect -4 36 76 87
<< polysilicon >>
rect 22 70 24 74
rect 29 70 31 74
rect 36 70 38 74
rect 46 70 48 74
rect 53 70 55 74
rect 60 70 62 74
rect 9 61 11 65
rect 9 39 11 42
rect 22 41 24 44
rect 19 40 25 41
rect 9 38 15 39
rect 9 34 10 38
rect 14 34 15 38
rect 9 33 15 34
rect 19 36 20 40
rect 24 36 25 40
rect 19 35 25 36
rect 29 35 31 44
rect 36 41 38 44
rect 46 41 48 44
rect 36 40 48 41
rect 36 39 41 40
rect 40 36 41 39
rect 45 39 48 40
rect 45 36 46 39
rect 40 35 46 36
rect 53 35 55 44
rect 60 41 62 44
rect 60 40 70 41
rect 60 39 65 40
rect 64 36 65 39
rect 69 36 70 40
rect 64 35 70 36
rect 9 30 11 33
rect 19 30 21 35
rect 29 34 35 35
rect 29 30 30 34
rect 34 30 35 34
rect 29 29 35 30
rect 40 26 42 35
rect 50 34 56 35
rect 50 30 51 34
rect 55 30 56 34
rect 50 29 56 30
rect 50 26 52 29
rect 9 9 11 14
rect 19 9 21 14
rect 40 6 42 10
rect 50 6 52 10
<< ndiffusion >>
rect 2 29 9 30
rect 2 25 3 29
rect 7 25 9 29
rect 2 22 9 25
rect 2 18 3 22
rect 7 18 9 22
rect 2 17 9 18
rect 4 14 9 17
rect 11 29 19 30
rect 11 25 13 29
rect 17 25 19 29
rect 11 22 19 25
rect 11 18 13 22
rect 17 18 19 22
rect 11 14 19 18
rect 21 26 26 30
rect 21 14 40 26
rect 23 12 40 14
rect 23 8 24 12
rect 28 8 33 12
rect 37 10 40 12
rect 42 21 50 26
rect 42 17 44 21
rect 48 17 50 21
rect 42 10 50 17
rect 52 22 59 26
rect 52 18 54 22
rect 58 18 59 22
rect 52 15 59 18
rect 52 11 54 15
rect 58 11 59 15
rect 52 10 59 11
rect 37 8 38 10
rect 23 7 38 8
<< pdiffusion >>
rect 13 69 22 70
rect 13 65 15 69
rect 19 65 22 69
rect 13 61 22 65
rect 2 60 9 61
rect 2 56 3 60
rect 7 56 9 60
rect 2 53 9 56
rect 2 49 3 53
rect 7 49 9 53
rect 2 48 9 49
rect 4 42 9 48
rect 11 44 22 61
rect 24 44 29 70
rect 31 44 36 70
rect 38 62 46 70
rect 38 58 40 62
rect 44 58 46 62
rect 38 44 46 58
rect 48 44 53 70
rect 55 44 60 70
rect 62 69 70 70
rect 62 65 64 69
rect 68 65 70 69
rect 62 62 70 65
rect 62 58 64 62
rect 68 58 70 62
rect 62 44 70 58
rect 11 42 16 44
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect -2 69 74 78
rect -2 68 15 69
rect 14 65 15 68
rect 19 68 64 69
rect 19 65 20 68
rect 63 65 64 68
rect 68 68 74 69
rect 68 65 69 68
rect 63 62 69 65
rect 2 60 40 62
rect 2 56 3 60
rect 7 58 40 60
rect 44 58 47 62
rect 63 58 64 62
rect 68 58 69 62
rect 2 53 7 56
rect 2 49 3 53
rect 2 48 7 49
rect 10 50 23 54
rect 31 50 70 54
rect 2 29 6 48
rect 10 38 14 50
rect 31 46 35 50
rect 10 33 14 34
rect 18 42 35 46
rect 41 42 55 46
rect 18 40 24 42
rect 18 36 20 40
rect 18 33 24 36
rect 41 40 47 42
rect 45 36 47 40
rect 30 34 34 35
rect 41 34 47 36
rect 65 40 70 50
rect 69 36 70 40
rect 65 35 70 36
rect 51 34 55 35
rect 13 29 17 30
rect 2 25 3 29
rect 7 25 8 29
rect 2 22 8 25
rect 2 18 3 22
rect 7 18 8 22
rect 2 17 8 18
rect 30 26 70 30
rect 13 22 17 25
rect 17 18 44 21
rect 13 17 44 18
rect 48 17 49 21
rect 53 18 54 22
rect 58 18 59 22
rect 53 15 59 18
rect 66 17 70 26
rect 53 12 54 15
rect -2 8 24 12
rect 28 8 33 12
rect 37 11 54 12
rect 58 12 59 15
rect 58 11 74 12
rect 37 8 74 11
rect -2 2 74 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
<< ntransistor >>
rect 9 14 11 30
rect 19 14 21 30
rect 40 10 42 26
rect 50 10 52 26
<< ptransistor >>
rect 9 42 11 61
rect 22 44 24 70
rect 29 44 31 70
rect 36 44 38 70
rect 46 44 48 70
rect 53 44 55 70
rect 60 44 62 70
<< polycontact >>
rect 10 34 14 38
rect 20 36 24 40
rect 41 36 45 40
rect 65 36 69 40
rect 30 30 34 34
rect 51 30 55 34
<< ndcontact >>
rect 3 25 7 29
rect 3 18 7 22
rect 13 25 17 29
rect 13 18 17 22
rect 24 8 28 12
rect 33 8 37 12
rect 44 17 48 21
rect 54 18 58 22
rect 54 11 58 15
<< pdcontact >>
rect 15 65 19 69
rect 3 56 7 60
rect 3 49 7 53
rect 40 58 44 62
rect 64 65 68 69
rect 64 58 68 62
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
<< psubstratepdiff >>
rect 0 2 72 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 72 2
rect 0 -3 72 -2
<< nsubstratendiff >>
rect 0 82 72 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 72 82
rect 0 77 72 78
<< labels >>
rlabel metal1 4 36 4 36 6 z
rlabel metal1 15 23 15 23 6 n3
rlabel metal1 12 40 12 40 6 b
rlabel metal1 20 36 20 36 6 a1
rlabel metal1 20 52 20 52 6 b
rlabel metal1 12 60 12 60 6 z
rlabel metal1 20 60 20 60 6 z
rlabel metal1 36 6 36 6 6 vss
rlabel metal1 36 28 36 28 6 a2
rlabel metal1 28 44 28 44 6 a1
rlabel metal1 36 52 36 52 6 a1
rlabel metal1 28 60 28 60 6 z
rlabel metal1 36 60 36 60 6 z
rlabel metal1 36 74 36 74 6 vdd
rlabel metal1 44 28 44 28 6 a2
rlabel metal1 31 19 31 19 6 n3
rlabel metal1 52 28 52 28 6 a2
rlabel metal1 44 40 44 40 6 a3
rlabel metal1 52 44 52 44 6 a3
rlabel metal1 52 52 52 52 6 a1
rlabel metal1 44 52 44 52 6 a1
rlabel metal1 44 60 44 60 6 z
rlabel metal1 60 28 60 28 6 a2
rlabel metal1 68 20 68 20 6 a2
rlabel metal1 68 44 68 44 6 a1
rlabel metal1 60 52 60 52 6 a1
<< end >>
