magic
tech scmos
timestamp 1182286862
<< checkpaint >>
rect -22 -25 190 105
<< ab >>
rect 0 0 168 80
<< pwell >>
rect -4 -7 172 36
<< nwell >>
rect -4 36 172 87
<< polysilicon >>
rect 9 69 11 74
rect 19 69 21 74
rect 29 72 53 74
rect 29 69 31 72
rect 39 69 41 72
rect 51 55 53 72
rect 62 70 64 74
rect 72 70 74 74
rect 82 70 84 74
rect 92 70 94 74
rect 112 70 114 74
rect 122 70 124 74
rect 132 70 134 74
rect 48 54 54 55
rect 48 50 49 54
rect 53 50 54 54
rect 48 49 54 50
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 39 39 41 42
rect 62 41 64 44
rect 72 41 74 44
rect 143 64 158 65
rect 143 63 153 64
rect 143 60 145 63
rect 152 60 153 63
rect 157 60 158 64
rect 152 59 158 60
rect 153 56 155 59
rect 143 42 145 46
rect 9 38 22 39
rect 9 37 17 38
rect 16 34 17 37
rect 21 34 22 38
rect 29 37 41 39
rect 61 39 74 41
rect 82 39 84 42
rect 92 39 94 42
rect 112 39 114 42
rect 122 39 124 42
rect 61 38 67 39
rect 16 33 22 34
rect 9 28 11 33
rect 16 31 28 33
rect 16 28 18 31
rect 26 28 28 31
rect 33 28 35 37
rect 61 35 62 38
rect 45 30 47 35
rect 55 34 62 35
rect 66 34 67 38
rect 79 38 108 39
rect 79 37 103 38
rect 79 35 81 37
rect 55 33 67 34
rect 55 30 57 33
rect 65 30 67 33
rect 75 33 81 35
rect 102 34 103 37
rect 107 34 108 38
rect 102 33 108 34
rect 112 38 118 39
rect 112 34 113 38
rect 117 34 118 38
rect 112 33 118 34
rect 122 38 128 39
rect 122 34 123 38
rect 127 34 128 38
rect 132 38 134 42
rect 132 37 146 38
rect 132 36 141 37
rect 122 33 128 34
rect 140 33 141 36
rect 145 33 146 37
rect 75 30 77 33
rect 85 32 91 33
rect 85 28 86 32
rect 90 29 91 32
rect 90 28 97 29
rect 85 27 97 28
rect 85 24 87 27
rect 95 24 97 27
rect 113 24 115 33
rect 122 29 124 33
rect 140 32 146 33
rect 140 29 142 32
rect 153 30 155 42
rect 120 27 124 29
rect 120 24 122 27
rect 130 24 132 29
rect 9 8 11 16
rect 16 12 18 16
rect 26 12 28 16
rect 33 8 35 16
rect 9 6 35 8
rect 45 8 47 16
rect 55 12 57 16
rect 65 12 67 16
rect 75 8 77 16
rect 45 6 77 8
rect 85 7 87 12
rect 95 7 97 12
rect 140 12 142 16
rect 113 6 115 11
rect 120 6 122 11
rect 130 8 132 11
rect 153 8 155 19
rect 130 6 155 8
<< ndiffusion >>
rect 37 28 45 30
rect 2 21 9 28
rect 2 17 3 21
rect 7 17 9 21
rect 2 16 9 17
rect 11 16 16 28
rect 18 27 26 28
rect 18 23 20 27
rect 24 23 26 27
rect 18 16 26 23
rect 28 16 33 28
rect 35 16 45 28
rect 47 29 55 30
rect 47 25 49 29
rect 53 25 55 29
rect 47 16 55 25
rect 57 22 65 30
rect 57 18 59 22
rect 63 18 65 22
rect 57 16 65 18
rect 67 29 75 30
rect 67 25 69 29
rect 73 25 75 29
rect 67 22 75 25
rect 67 18 69 22
rect 73 18 75 22
rect 67 16 75 18
rect 77 24 82 30
rect 148 29 153 30
rect 135 24 140 29
rect 77 21 85 24
rect 77 17 79 21
rect 83 17 85 21
rect 77 16 85 17
rect 37 12 43 16
rect 37 8 38 12
rect 42 8 43 12
rect 37 7 43 8
rect 80 12 85 16
rect 87 22 95 24
rect 87 18 89 22
rect 93 18 95 22
rect 87 12 95 18
rect 97 15 113 24
rect 97 12 103 15
rect 99 11 103 12
rect 107 11 113 15
rect 115 11 120 24
rect 122 22 130 24
rect 122 18 124 22
rect 128 18 130 22
rect 122 11 130 18
rect 132 23 140 24
rect 132 19 134 23
rect 138 19 140 23
rect 132 16 140 19
rect 142 22 153 29
rect 142 18 146 22
rect 150 19 153 22
rect 155 29 162 30
rect 155 25 157 29
rect 161 25 162 29
rect 155 24 162 25
rect 155 19 160 24
rect 150 18 151 19
rect 142 16 151 18
rect 132 11 137 16
rect 99 9 111 11
<< pdiffusion >>
rect 4 62 9 69
rect 2 61 9 62
rect 2 57 3 61
rect 7 57 9 61
rect 2 54 9 57
rect 2 50 3 54
rect 7 50 9 54
rect 2 49 9 50
rect 4 42 9 49
rect 11 54 19 69
rect 11 50 13 54
rect 17 50 19 54
rect 11 47 19 50
rect 11 43 13 47
rect 17 43 19 47
rect 11 42 19 43
rect 21 62 29 69
rect 21 58 23 62
rect 27 58 29 62
rect 21 42 29 58
rect 31 47 39 69
rect 31 43 33 47
rect 37 43 39 47
rect 31 42 39 43
rect 41 63 46 69
rect 41 62 49 63
rect 41 58 44 62
rect 48 58 49 62
rect 41 57 49 58
rect 41 42 46 57
rect 160 72 166 73
rect 55 69 62 70
rect 55 65 56 69
rect 60 65 62 69
rect 55 62 62 65
rect 55 58 56 62
rect 60 58 62 62
rect 55 57 62 58
rect 56 44 62 57
rect 64 61 72 70
rect 64 57 66 61
rect 70 57 72 61
rect 64 54 72 57
rect 64 50 66 54
rect 70 50 72 54
rect 64 44 72 50
rect 74 69 82 70
rect 74 65 76 69
rect 80 65 82 69
rect 74 62 82 65
rect 74 58 76 62
rect 80 58 82 62
rect 74 44 82 58
rect 77 42 82 44
rect 84 47 92 70
rect 84 43 86 47
rect 90 43 92 47
rect 84 42 92 43
rect 94 69 101 70
rect 94 65 96 69
rect 100 65 101 69
rect 94 62 101 65
rect 107 63 112 70
rect 94 58 96 62
rect 100 58 101 62
rect 94 42 101 58
rect 105 62 112 63
rect 105 58 106 62
rect 110 58 112 62
rect 105 57 112 58
rect 107 42 112 57
rect 114 55 122 70
rect 114 51 116 55
rect 120 51 122 55
rect 114 42 122 51
rect 124 54 132 70
rect 124 50 126 54
rect 130 50 132 54
rect 124 47 132 50
rect 124 43 126 47
rect 130 43 132 47
rect 124 42 132 43
rect 134 69 141 70
rect 134 65 136 69
rect 140 65 141 69
rect 160 68 161 72
rect 165 68 166 72
rect 134 60 141 65
rect 134 46 143 60
rect 145 56 150 60
rect 160 56 166 68
rect 145 51 153 56
rect 145 47 147 51
rect 151 47 153 51
rect 145 46 153 47
rect 134 42 141 46
rect 148 42 153 46
rect 155 42 166 56
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect 118 78 122 82
rect 126 78 130 82
rect 134 78 138 82
rect 142 78 146 82
rect 150 78 154 82
rect 158 78 162 82
rect 166 78 170 82
rect -2 72 170 78
rect -2 69 161 72
rect -2 68 56 69
rect 55 65 56 68
rect 60 68 76 69
rect 60 65 61 68
rect 55 62 61 65
rect 75 65 76 68
rect 80 68 96 69
rect 80 65 81 68
rect 75 62 81 65
rect 2 61 23 62
rect 2 57 3 61
rect 7 58 23 61
rect 27 58 44 62
rect 48 58 49 62
rect 55 58 56 62
rect 60 58 61 62
rect 66 61 70 62
rect 2 54 7 57
rect 75 58 76 62
rect 80 58 81 62
rect 95 65 96 68
rect 100 68 136 69
rect 100 65 101 68
rect 135 65 136 68
rect 140 68 161 69
rect 165 68 170 72
rect 140 65 141 68
rect 95 62 101 65
rect 95 58 96 62
rect 100 58 101 62
rect 105 58 106 62
rect 110 58 138 62
rect 66 54 70 57
rect 2 50 3 54
rect 2 49 7 50
rect 12 50 13 54
rect 17 50 49 54
rect 53 50 66 54
rect 70 50 99 54
rect 2 30 6 49
rect 12 47 17 50
rect 12 43 13 47
rect 12 42 17 43
rect 32 43 33 47
rect 37 43 38 47
rect 85 46 86 47
rect 32 38 38 43
rect 48 43 86 46
rect 90 43 91 47
rect 48 42 91 43
rect 48 38 52 42
rect 16 34 17 38
rect 21 34 52 38
rect 57 34 62 38
rect 66 34 87 38
rect 2 27 24 30
rect 2 26 20 27
rect 48 29 52 34
rect 81 32 87 34
rect 48 25 49 29
rect 53 25 69 29
rect 73 25 74 29
rect 81 28 86 32
rect 90 28 91 32
rect 81 26 87 28
rect 20 22 24 23
rect 69 22 74 25
rect 95 22 99 50
rect 3 21 7 22
rect 20 18 59 22
rect 63 18 64 22
rect 73 18 74 22
rect 69 17 74 18
rect 79 21 83 22
rect 88 18 89 22
rect 93 18 99 22
rect 103 51 116 55
rect 120 51 121 55
rect 126 54 130 55
rect 103 38 107 51
rect 126 47 130 50
rect 103 22 107 34
rect 113 43 126 46
rect 113 42 130 43
rect 134 46 138 58
rect 152 60 153 64
rect 157 63 158 64
rect 157 60 166 63
rect 152 57 166 60
rect 147 51 151 52
rect 162 49 166 57
rect 147 46 151 47
rect 134 42 166 46
rect 113 38 117 42
rect 134 38 138 42
rect 145 38 158 39
rect 122 34 123 38
rect 127 34 138 38
rect 141 37 158 38
rect 113 30 117 34
rect 145 33 158 37
rect 141 32 151 33
rect 113 26 138 30
rect 145 26 151 32
rect 162 29 166 42
rect 134 23 138 26
rect 156 25 157 29
rect 161 25 166 29
rect 103 18 124 22
rect 128 18 129 22
rect 134 18 138 19
rect 145 18 146 22
rect 150 18 151 22
rect 3 12 7 17
rect 79 12 83 17
rect 102 12 103 15
rect -2 8 38 12
rect 42 11 103 12
rect 107 12 108 15
rect 145 12 151 18
rect 107 11 170 12
rect 42 8 170 11
rect -2 2 170 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 122 2
rect 126 -2 130 2
rect 134 -2 138 2
rect 142 -2 146 2
rect 150 -2 154 2
rect 158 -2 162 2
rect 166 -2 170 2
<< ntransistor >>
rect 9 16 11 28
rect 16 16 18 28
rect 26 16 28 28
rect 33 16 35 28
rect 45 16 47 30
rect 55 16 57 30
rect 65 16 67 30
rect 75 16 77 30
rect 85 12 87 24
rect 95 12 97 24
rect 113 11 115 24
rect 120 11 122 24
rect 130 11 132 24
rect 140 16 142 29
rect 153 19 155 30
<< ptransistor >>
rect 9 42 11 69
rect 19 42 21 69
rect 29 42 31 69
rect 39 42 41 69
rect 62 44 64 70
rect 72 44 74 70
rect 82 42 84 70
rect 92 42 94 70
rect 112 42 114 70
rect 122 42 124 70
rect 132 42 134 70
rect 143 46 145 60
rect 153 42 155 56
<< polycontact >>
rect 49 50 53 54
rect 153 60 157 64
rect 17 34 21 38
rect 62 34 66 38
rect 103 34 107 38
rect 113 34 117 38
rect 123 34 127 38
rect 141 33 145 37
rect 86 28 90 32
<< ndcontact >>
rect 3 17 7 21
rect 20 23 24 27
rect 49 25 53 29
rect 59 18 63 22
rect 69 25 73 29
rect 69 18 73 22
rect 79 17 83 21
rect 38 8 42 12
rect 89 18 93 22
rect 103 11 107 15
rect 124 18 128 22
rect 134 19 138 23
rect 146 18 150 22
rect 157 25 161 29
<< pdcontact >>
rect 3 57 7 61
rect 3 50 7 54
rect 13 50 17 54
rect 13 43 17 47
rect 23 58 27 62
rect 33 43 37 47
rect 44 58 48 62
rect 56 65 60 69
rect 56 58 60 62
rect 66 57 70 61
rect 66 50 70 54
rect 76 65 80 69
rect 76 58 80 62
rect 86 43 90 47
rect 96 65 100 69
rect 96 58 100 62
rect 106 58 110 62
rect 116 51 120 55
rect 126 50 130 54
rect 126 43 130 47
rect 136 65 140 69
rect 161 68 165 72
rect 147 47 151 51
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
rect 58 -2 62 2
rect 66 -2 70 2
rect 74 -2 78 2
rect 82 -2 86 2
rect 90 -2 94 2
rect 98 -2 102 2
rect 106 -2 110 2
rect 114 -2 118 2
rect 122 -2 126 2
rect 130 -2 134 2
rect 138 -2 142 2
rect 146 -2 150 2
rect 154 -2 158 2
rect 162 -2 166 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
rect 58 78 62 82
rect 66 78 70 82
rect 74 78 78 82
rect 82 78 86 82
rect 90 78 94 82
rect 98 78 102 82
rect 106 78 110 82
rect 114 78 118 82
rect 122 78 126 82
rect 130 78 134 82
rect 138 78 142 82
rect 146 78 150 82
rect 154 78 158 82
rect 162 78 166 82
<< psubstratepdiff >>
rect 0 2 168 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
rect 62 -2 66 2
rect 70 -2 74 2
rect 78 -2 82 2
rect 86 -2 90 2
rect 94 -2 98 2
rect 102 -2 106 2
rect 110 -2 114 2
rect 118 -2 122 2
rect 126 -2 130 2
rect 134 -2 138 2
rect 142 -2 146 2
rect 150 -2 154 2
rect 158 -2 162 2
rect 166 -2 168 2
rect 0 -3 168 -2
<< nsubstratendiff >>
rect 0 82 168 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect 62 78 66 82
rect 70 78 74 82
rect 78 78 82 82
rect 86 78 90 82
rect 94 78 98 82
rect 102 78 106 82
rect 110 78 114 82
rect 118 78 122 82
rect 126 78 130 82
rect 134 78 138 82
rect 142 78 146 82
rect 150 78 154 82
rect 158 78 162 82
rect 166 78 168 82
rect 0 77 168 78
<< labels >>
rlabel polysilicon 52 61 52 61 6 cn
rlabel ntransistor 114 22 114 22 6 an
rlabel polycontact 105 36 105 36 6 iz
rlabel polycontact 125 36 125 36 6 bn
rlabel metal1 20 28 20 28 6 z
rlabel metal1 12 28 12 28 6 z
rlabel metal1 28 20 28 20 6 z
rlabel metal1 4 44 4 44 6 z
rlabel metal1 14 48 14 48 6 cn
rlabel metal1 12 60 12 60 6 z
rlabel metal1 20 60 20 60 6 z
rlabel metal1 28 60 28 60 6 z
rlabel metal1 36 20 36 20 6 z
rlabel metal1 44 20 44 20 6 z
rlabel metal1 52 20 52 20 6 z
rlabel ndcontact 60 20 60 20 6 z
rlabel metal1 35 40 35 40 6 zn
rlabel metal1 60 36 60 36 6 c
rlabel metal1 36 60 36 60 6 z
rlabel metal1 44 60 44 60 6 z
rlabel metal1 84 6 84 6 6 vss
rlabel metal1 61 27 61 27 6 zn
rlabel metal1 71 23 71 23 6 zn
rlabel metal1 93 20 93 20 6 cn
rlabel metal1 84 32 84 32 6 c
rlabel metal1 68 36 68 36 6 c
rlabel metal1 69 44 69 44 6 zn
rlabel metal1 76 36 76 36 6 c
rlabel metal1 68 56 68 56 6 cn
rlabel metal1 55 52 55 52 6 cn
rlabel metal1 84 74 84 74 6 vdd
rlabel metal1 116 20 116 20 6 iz
rlabel polycontact 115 36 115 36 6 an
rlabel metal1 128 48 128 48 6 an
rlabel polycontact 105 36 105 36 6 iz
rlabel metal1 112 53 112 53 6 iz
rlabel metal1 136 24 136 24 6 an
rlabel metal1 161 27 161 27 6 bn
rlabel metal1 148 32 148 32 6 a
rlabel metal1 130 36 130 36 6 bn
rlabel metal1 156 36 156 36 6 a
rlabel metal1 149 47 149 47 6 bn
rlabel metal1 121 60 121 60 6 bn
rlabel metal1 156 60 156 60 6 b
rlabel metal1 164 56 164 56 6 b
<< end >>
