.subckt nd3_x2 a b c vdd vss z
*   SPICE3 file   created from nd3_x2.ext -      technology: scmos
m00 vdd    c      z      vdd p w=33u  l=2.3636u ad=198p     pd=56u      as=179p     ps=56u
m01 z      b      vdd    vdd p w=33u  l=2.3636u ad=179p     pd=56u      as=198p     ps=56u
m02 vdd    a      z      vdd p w=33u  l=2.3636u ad=198p     pd=56u      as=179p     ps=56u
m03 w1     c      z      vss n w=33u  l=2.3636u ad=99p      pd=39u      as=183p     ps=82u
m04 w2     b      w1     vss n w=33u  l=2.3636u ad=99p      pd=39u      as=99p      ps=39u
m05 vss    a      w2     vss n w=33u  l=2.3636u ad=264p     pd=82u      as=99p      ps=39u
C0  vss    c      0.022f
C1  vdd    b      0.042f
C2  z      a      0.088f
C3  z      c      0.184f
C4  a      b      0.186f
C5  w2     vss    0.011f
C6  b      c      0.185f
C7  vss    z      0.078f
C8  w1     a      0.013f
C9  w1     c      0.006f
C10 vdd    a      0.008f
C11 vss    b      0.010f
C12 z      b      0.136f
C13 vdd    c      0.019f
C14 a      c      0.168f
C15 w1     vss    0.011f
C16 w2     a      0.013f
C17 w2     c      0.002f
C18 vdd    z      0.201f
C19 vss    a      0.071f
C22 z      vss    0.022f
C23 a      vss    0.021f
C24 b      vss    0.028f
C25 c      vss    0.030f
.ends
