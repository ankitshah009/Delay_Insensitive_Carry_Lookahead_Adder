magic
tech scmos
timestamp 1185094827
<< checkpaint >>
rect -22 -22 82 122
<< ab >>
rect 0 0 60 100
<< pwell >>
rect -4 -4 64 48
<< nwell >>
rect -4 48 64 104
<< metal1 >>
rect -2 96 62 100
rect -2 92 4 96
rect 8 92 13 96
rect 17 92 23 96
rect 27 92 33 96
rect 37 92 43 96
rect 47 92 52 96
rect 56 92 62 96
rect -2 88 62 92
rect -2 8 62 12
rect -2 4 4 8
rect 8 4 13 8
rect 17 4 23 8
rect 27 4 33 8
rect 37 4 43 8
rect 47 4 52 8
rect 56 4 62 8
rect -2 0 62 4
<< psubstratepcontact >>
rect 4 4 8 8
rect 13 4 17 8
rect 23 4 27 8
rect 33 4 37 8
rect 43 4 47 8
rect 52 4 56 8
<< nsubstratencontact >>
rect 4 92 8 96
rect 13 92 17 96
rect 23 92 27 96
rect 33 92 37 96
rect 43 92 47 96
rect 52 92 56 96
<< psubstratepdiff >>
rect 3 8 57 39
rect 3 4 4 8
rect 8 4 13 8
rect 17 4 23 8
rect 27 4 33 8
rect 37 4 43 8
rect 47 4 52 8
rect 56 4 57 8
rect 3 3 57 4
<< nsubstratendiff >>
rect 3 96 57 97
rect 3 92 4 96
rect 8 92 13 96
rect 17 92 23 96
rect 27 92 33 96
rect 37 92 43 96
rect 47 92 52 96
rect 56 92 57 96
rect 3 55 57 92
<< labels >>
rlabel metal1 30 6 30 6 6 vss
rlabel metal1 30 94 30 94 6 vdd
<< end >>
