.subckt noa22_x4 i0 i1 i2 nq vdd vss
*   SPICE3 file   created from noa22_x4.ext -      technology: scmos
m00 w1     i2     vdd    vdd p w=20u  l=2.3636u ad=120p     pd=38.6667u as=148p     ps=44.6667u
m01 w2     i1     w1     vdd p w=20u  l=2.3636u ad=100p     pd=30u      as=120p     ps=38.6667u
m02 w1     i0     w2     vdd p w=20u  l=2.3636u ad=120p     pd=38.6667u as=100p     ps=30u
m03 vdd    w2     w3     vdd p w=20u  l=2.3636u ad=148p     pd=44.6667u as=160p     ps=56u
m04 nq     w3     vdd    vdd p w=40u  l=2.3636u ad=200p     pd=50u      as=296p     ps=89.3333u
m05 vdd    w3     nq     vdd p w=40u  l=2.3636u ad=296p     pd=89.3333u as=200p     ps=50u
m06 w2     i2     vss    vss n w=10u  l=2.3636u ad=50p      pd=20u      as=85.1429p ps=31.4286u
m07 w4     i1     w2     vss n w=10u  l=2.3636u ad=50p      pd=20u      as=50p      ps=20u
m08 vss    i0     w4     vss n w=10u  l=2.3636u ad=85.1429p pd=31.4286u as=50p      ps=20u
m09 vss    w2     w3     vss n w=10u  l=2.3636u ad=85.1429p pd=31.4286u as=80p      ps=36u
m10 nq     w3     vss    vss n w=20u  l=2.3636u ad=100p     pd=30u      as=170.286p ps=62.8571u
m11 vss    w3     nq     vss n w=20u  l=2.3636u ad=170.286p pd=62.8571u as=100p     ps=30u
C0  vss    i2     0.055f
C1  w2     i0     0.173f
C2  w1     i1     0.017f
C3  w2     i2     0.339f
C4  nq     w3     0.132f
C5  vss    vdd    0.005f
C6  w2     vdd    0.183f
C7  i0     i2     0.090f
C8  vss    nq     0.130f
C9  i0     vdd    0.010f
C10 i1     w3     0.069f
C11 nq     w2     0.088f
C12 w4     i0     0.004f
C13 i2     vdd    0.074f
C14 w2     w1     0.218f
C15 nq     i0     0.039f
C16 vss    i1     0.047f
C17 w2     i1     0.346f
C18 w1     i0     0.017f
C19 vss    w3     0.116f
C20 w2     w3     0.349f
C21 nq     vdd    0.231f
C22 w1     i2     0.039f
C23 i0     i1     0.425f
C24 i0     w3     0.142f
C25 w1     vdd    0.230f
C26 i1     i2     0.172f
C27 vss    w2     0.064f
C28 i2     w3     0.034f
C29 i1     vdd    0.011f
C30 nq     w1     0.006f
C31 vss    i0     0.058f
C32 w4     i1     0.016f
C33 w3     vdd    0.031f
C35 nq     vss    0.018f
C36 w2     vss    0.046f
C37 i0     vss    0.040f
C38 i1     vss    0.050f
C39 i2     vss    0.052f
C40 w3     vss    0.069f
.ends
