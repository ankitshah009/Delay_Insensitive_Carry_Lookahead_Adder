magic
tech scmos
timestamp 1179387702
<< checkpaint >>
rect -22 -22 94 94
<< ab >>
rect 0 0 72 72
<< pwell >>
rect -4 -4 76 32
<< nwell >>
rect -4 32 76 76
<< polysilicon >>
rect 9 66 11 70
rect 19 66 21 70
rect 29 66 31 70
rect 40 66 42 70
rect 50 66 52 70
rect 40 49 42 52
rect 50 49 52 52
rect 40 48 63 49
rect 40 47 42 48
rect 41 44 42 47
rect 46 47 63 48
rect 46 44 47 47
rect 41 43 47 44
rect 9 35 11 38
rect 19 35 21 38
rect 29 35 31 38
rect 9 34 15 35
rect 9 30 10 34
rect 14 30 15 34
rect 9 29 15 30
rect 19 34 25 35
rect 19 30 20 34
rect 24 30 25 34
rect 29 32 33 35
rect 19 29 25 30
rect 12 26 14 29
rect 19 26 21 29
rect 31 26 33 32
rect 41 26 43 43
rect 51 34 57 35
rect 51 30 52 34
rect 56 30 57 34
rect 51 29 57 30
rect 51 26 53 29
rect 61 26 63 47
rect 12 2 14 7
rect 19 2 21 7
rect 31 4 33 19
rect 61 14 63 19
rect 41 8 43 12
rect 51 4 53 12
rect 31 2 53 4
<< ndiffusion >>
rect 7 19 12 26
rect 5 18 12 19
rect 5 14 6 18
rect 10 14 12 18
rect 5 13 12 14
rect 7 7 12 13
rect 14 7 19 26
rect 21 19 31 26
rect 33 25 41 26
rect 33 21 35 25
rect 39 21 41 25
rect 33 19 41 21
rect 21 8 29 19
rect 21 7 24 8
rect 23 4 24 7
rect 28 4 29 8
rect 23 3 29 4
rect 36 12 41 19
rect 43 18 51 26
rect 43 14 45 18
rect 49 14 51 18
rect 43 12 51 14
rect 53 25 61 26
rect 53 21 55 25
rect 59 21 61 25
rect 53 19 61 21
rect 63 24 70 26
rect 63 20 65 24
rect 69 20 70 24
rect 63 19 70 20
rect 53 12 58 19
<< pdiffusion >>
rect 4 59 9 66
rect 2 58 9 59
rect 2 54 3 58
rect 7 54 9 58
rect 2 53 9 54
rect 4 38 9 53
rect 11 50 19 66
rect 11 46 13 50
rect 17 46 19 50
rect 11 38 19 46
rect 21 50 29 66
rect 21 46 23 50
rect 27 46 29 50
rect 21 43 29 46
rect 21 39 23 43
rect 27 39 29 43
rect 21 38 29 39
rect 31 65 40 66
rect 31 61 34 65
rect 38 61 40 65
rect 31 52 40 61
rect 42 58 50 66
rect 42 54 44 58
rect 48 54 50 58
rect 42 52 50 54
rect 52 65 59 66
rect 52 61 54 65
rect 58 61 59 65
rect 52 58 59 61
rect 52 54 54 58
rect 58 54 59 58
rect 52 52 59 54
rect 31 38 38 52
<< metal1 >>
rect -2 68 74 72
rect -2 65 64 68
rect -2 64 34 65
rect 33 61 34 64
rect 38 64 54 65
rect 38 61 39 64
rect 53 61 54 64
rect 58 64 64 65
rect 68 64 74 68
rect 58 61 59 64
rect 53 58 59 61
rect 2 54 3 58
rect 7 54 44 58
rect 48 54 49 58
rect 53 54 54 58
rect 58 54 59 58
rect 23 50 27 51
rect 2 46 13 50
rect 17 46 18 50
rect 2 14 6 46
rect 23 43 27 46
rect 10 39 23 42
rect 10 38 27 39
rect 10 34 14 38
rect 31 34 35 54
rect 41 48 55 50
rect 41 44 42 48
rect 46 44 55 48
rect 49 38 55 44
rect 66 34 70 43
rect 19 30 20 34
rect 24 30 48 34
rect 10 26 14 30
rect 10 25 40 26
rect 10 22 35 25
rect 34 21 35 22
rect 39 21 40 25
rect 44 25 48 30
rect 51 30 52 34
rect 56 30 70 34
rect 51 29 70 30
rect 44 21 55 25
rect 59 21 60 25
rect 65 24 69 25
rect 10 14 45 18
rect 49 14 50 18
rect 65 8 69 20
rect -2 4 24 8
rect 28 4 64 8
rect 68 4 74 8
rect -2 0 74 4
<< ntransistor >>
rect 12 7 14 26
rect 19 7 21 26
rect 31 19 33 26
rect 41 12 43 26
rect 51 12 53 26
rect 61 19 63 26
<< ptransistor >>
rect 9 38 11 66
rect 19 38 21 66
rect 29 38 31 66
rect 40 52 42 66
rect 50 52 52 66
<< polycontact >>
rect 42 44 46 48
rect 10 30 14 34
rect 20 30 24 34
rect 52 30 56 34
<< ndcontact >>
rect 6 14 10 18
rect 35 21 39 25
rect 24 4 28 8
rect 45 14 49 18
rect 55 21 59 25
rect 65 20 69 24
<< pdcontact >>
rect 3 54 7 58
rect 13 46 17 50
rect 23 46 27 50
rect 23 39 27 43
rect 34 61 38 65
rect 44 54 48 58
rect 54 61 58 65
rect 54 54 58 58
<< psubstratepcontact >>
rect 64 4 68 8
<< nsubstratencontact >>
rect 64 64 68 68
<< psubstratepdiff >>
rect 63 8 69 9
rect 63 4 64 8
rect 68 4 69 8
rect 63 3 69 4
<< nsubstratendiff >>
rect 63 68 69 69
rect 63 64 64 68
rect 68 64 69 68
rect 63 52 69 64
<< labels >>
rlabel polycontact 12 32 12 32 6 bn
rlabel polycontact 22 32 22 32 6 an
rlabel metal1 12 16 12 16 6 z
rlabel metal1 4 32 4 32 6 z
rlabel polycontact 12 32 12 32 6 bn
rlabel metal1 12 48 12 48 6 z
rlabel metal1 28 16 28 16 6 z
rlabel metal1 20 16 20 16 6 z
rlabel metal1 25 44 25 44 6 bn
rlabel metal1 33 44 33 44 6 an
rlabel metal1 36 4 36 4 6 vss
rlabel metal1 44 16 44 16 6 z
rlabel metal1 36 16 36 16 6 z
rlabel metal1 25 24 25 24 6 bn
rlabel metal1 44 48 44 48 6 a
rlabel metal1 52 44 52 44 6 a
rlabel metal1 25 56 25 56 6 an
rlabel metal1 36 68 36 68 6 vdd
rlabel metal1 52 23 52 23 6 an
rlabel metal1 60 32 60 32 6 b
rlabel metal1 68 36 68 36 6 b
<< end >>
