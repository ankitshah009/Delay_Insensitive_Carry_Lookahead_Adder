.subckt oai31v0x1 a1 a2 a3 b vdd vss z
*   SPICE3 file   created from oai31v0x1.ext -      technology: scmos
m00 vdd    b      z      vdd p w=19u  l=2.3636u ad=130.056p pd=39.0704u as=88.0423p ps=32.1127u
m01 w1     a1     vdd    vdd p w=26u  l=2.3636u ad=65p      pd=31u      as=177.972p ps=53.4648u
m02 w2     a2     w1     vdd p w=26u  l=2.3636u ad=65p      pd=31u      as=65p      ps=31u
m03 z      a3     w2     vdd p w=26u  l=2.3636u ad=120.479p pd=43.9437u as=65p      ps=31u
m04 w3     a3     z      vdd p w=26u  l=2.3636u ad=65p      pd=31u      as=120.479p ps=43.9437u
m05 w4     a2     w3     vdd p w=26u  l=2.3636u ad=65p      pd=31u      as=65p      ps=31u
m06 vdd    a1     w4     vdd p w=26u  l=2.3636u ad=177.972p pd=53.4648u as=65p      ps=31u
m07 n3     b      z      vss n w=16u  l=2.3636u ad=64p      pd=24u      as=106p     ps=46u
m08 vss    a1     n3     vss n w=16u  l=2.3636u ad=157.667p pd=43.3333u as=64p      ps=24u
m09 n3     a3     vss    vss n w=16u  l=2.3636u ad=64p      pd=24u      as=157.667p ps=43.3333u
m10 vss    a2     n3     vss n w=16u  l=2.3636u ad=157.667p pd=43.3333u as=64p      ps=24u
C0  a2     a1     0.243f
C1  a3     vdd    0.027f
C2  w4     a3     0.001f
C3  w2     z      0.010f
C4  n3     a2     0.136f
C5  vss    a1     0.055f
C6  a1     vdd    0.171f
C7  vss    n3     0.294f
C8  n3     vdd    0.003f
C9  w4     a1     0.010f
C10 z      a3     0.043f
C11 w3     vdd    0.005f
C12 w2     a1     0.016f
C13 w1     vdd    0.005f
C14 b      a2     0.024f
C15 z      a1     0.218f
C16 n3     z      0.106f
C17 vss    b      0.016f
C18 a3     a1     0.224f
C19 b      vdd    0.061f
C20 n3     a3     0.022f
C21 vss    a2     0.169f
C22 a2     vdd    0.042f
C23 w1     z      0.010f
C24 n3     a1     0.051f
C25 w3     a3     0.005f
C26 w4     vdd    0.005f
C27 z      b      0.278f
C28 w3     a1     0.010f
C29 w2     vdd    0.005f
C30 b      a3     0.022f
C31 z      a2     0.036f
C32 w1     a1     0.005f
C33 vss    z      0.037f
C34 b      a1     0.213f
C35 a3     a2     0.234f
C36 z      vdd    0.295f
C37 vss    a3     0.021f
C38 n3     b      0.021f
C40 z      vss    0.008f
C41 b      vss    0.015f
C42 a3     vss    0.026f
C43 a2     vss    0.050f
C44 a1     vss    0.034f
.ends
