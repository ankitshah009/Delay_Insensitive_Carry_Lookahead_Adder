.subckt vddtie vdd vss z
*   SPICE3 file   created from vddtie.ext -      technology: scmos
m00 z      w1     vdd    vdd p w=28u  l=2.3636u ad=176p     pd=50u      as=196p     ps=70u
m01 vdd    w2     z      vdd p w=28u  l=2.3636u ad=196p     pd=70u      as=176p     ps=50u
m02 z      w1     w3     vss n w=20u  l=2.3636u ad=136p     pd=42u      as=140p     ps=54u
m03 w4     w2     z      vss n w=20u  l=2.3636u ad=140p     pd=54u      as=136p     ps=42u
C0  z      vdd    0.105f
C1  vss    w2     0.025f
C2  vss    w1     0.025f
C3  w2     z      0.007f
C4  z      w1     0.007f
C5  w2     vdd    0.021f
C6  w1     vdd    0.021f
C7  vss    z      0.045f
C8  w2     w1     0.065f
C10 w2     vss    0.043f
C11 z      vss    0.006f
C12 w1     vss    0.043f
.ends
