.subckt no2_x1 i0 i1 nq vdd vss
*   SPICE3 file   created from no2_x1.ext -      technology: scmos
m00 w1     i1     nq     vdd p w=40u  l=2.3636u ad=120p     pd=46u      as=400p     ps=104u
m01 vdd    i0     w1     vdd p w=40u  l=2.3636u ad=320p     pd=96u      as=120p     ps=46u
m02 nq     i1     vss    vss n w=10u  l=2.3636u ad=50p      pd=20u      as=128p     ps=52u
m03 vss    i0     nq     vss n w=10u  l=2.3636u ad=128p     pd=52u      as=50p      ps=20u
C0  vdd    nq     0.055f
C1  vss    i0     0.055f
C2  w1     i0     0.014f
C3  vdd    i1     0.041f
C4  nq     i1     0.508f
C5  vdd    w1     0.014f
C6  vss    nq     0.138f
C7  vdd    i0     0.082f
C8  vss    i1     0.015f
C9  w1     i1     0.027f
C10 nq     i0     0.166f
C11 i0     i1     0.488f
C14 nq     vss    0.022f
C15 i0     vss    0.037f
C16 i1     vss    0.037f
.ends
