magic
tech scmos
timestamp 1179385288
<< checkpaint >>
rect -22 -25 78 105
<< ab >>
rect 0 0 56 80
<< pwell >>
rect -4 -7 60 36
<< nwell >>
rect -4 36 60 87
<< polysilicon >>
rect 9 66 11 71
rect 19 66 21 71
rect 29 66 31 71
rect 41 61 43 65
rect 9 33 11 50
rect 19 47 21 50
rect 29 47 31 50
rect 16 46 22 47
rect 16 42 17 46
rect 21 42 22 46
rect 16 41 22 42
rect 26 46 32 47
rect 26 42 27 46
rect 31 42 32 46
rect 26 41 32 42
rect 9 32 15 33
rect 9 28 10 32
rect 14 28 15 32
rect 9 27 15 28
rect 13 24 15 27
rect 20 24 22 41
rect 30 24 32 41
rect 41 39 43 45
rect 37 38 43 39
rect 37 34 38 38
rect 42 34 43 38
rect 37 33 43 34
rect 37 24 39 33
rect 13 12 15 17
rect 20 12 22 17
rect 30 12 32 17
rect 37 12 39 17
<< ndiffusion >>
rect 4 17 13 24
rect 15 17 20 24
rect 22 22 30 24
rect 22 18 24 22
rect 28 18 30 22
rect 22 17 30 18
rect 32 17 37 24
rect 39 22 48 24
rect 39 18 42 22
rect 46 18 48 22
rect 39 17 48 18
rect 4 12 11 17
rect 4 8 6 12
rect 10 8 11 12
rect 4 7 11 8
<< pdiffusion >>
rect 33 72 39 73
rect 33 68 34 72
rect 38 68 39 72
rect 33 66 39 68
rect 4 64 9 66
rect 2 63 9 64
rect 2 59 3 63
rect 7 59 9 63
rect 2 58 9 59
rect 4 50 9 58
rect 11 55 19 66
rect 11 51 13 55
rect 17 51 19 55
rect 11 50 19 51
rect 21 63 29 66
rect 21 59 23 63
rect 27 59 29 63
rect 21 56 29 59
rect 21 52 23 56
rect 27 52 29 56
rect 21 50 29 52
rect 31 61 39 66
rect 31 50 41 61
rect 34 45 41 50
rect 43 60 50 61
rect 43 56 45 60
rect 49 56 50 60
rect 43 53 50 56
rect 43 49 45 53
rect 49 49 50 53
rect 43 48 50 49
rect 43 45 48 48
<< metal1 >>
rect -2 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 58 82
rect -2 72 58 78
rect -2 68 34 72
rect 38 68 58 72
rect 2 59 3 63
rect 7 59 23 63
rect 27 60 50 63
rect 27 59 45 60
rect 23 56 27 59
rect 2 51 13 55
rect 17 51 18 55
rect 44 56 45 59
rect 49 56 50 60
rect 23 51 27 52
rect 2 22 6 51
rect 10 46 21 47
rect 34 46 38 55
rect 44 53 50 56
rect 44 49 45 53
rect 49 49 50 53
rect 10 42 17 46
rect 25 42 27 46
rect 31 42 47 46
rect 10 41 21 42
rect 17 38 21 41
rect 17 34 23 38
rect 27 34 38 38
rect 10 32 14 33
rect 14 28 38 30
rect 10 26 38 28
rect 2 18 24 22
rect 28 18 29 22
rect 2 17 29 18
rect 34 17 38 26
rect 42 25 47 38
rect 41 18 42 22
rect 46 18 47 22
rect 41 12 47 18
rect -2 8 6 12
rect 10 8 58 12
rect -2 2 58 8
rect -2 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 58 2
<< ntransistor >>
rect 13 17 15 24
rect 20 17 22 24
rect 30 17 32 24
rect 37 17 39 24
<< ptransistor >>
rect 9 50 11 66
rect 19 50 21 66
rect 29 50 31 66
rect 41 45 43 61
<< polycontact >>
rect 17 42 21 46
rect 27 42 31 46
rect 10 28 14 32
rect 38 34 42 38
<< ndcontact >>
rect 24 18 28 22
rect 42 18 46 22
rect 6 8 10 12
<< pdcontact >>
rect 34 68 38 72
rect 3 59 7 63
rect 13 51 17 55
rect 23 59 27 63
rect 23 52 27 56
rect 45 56 49 60
rect 45 49 49 53
<< psubstratepcontact >>
rect 2 -2 6 2
rect 10 -2 14 2
rect 18 -2 22 2
rect 26 -2 30 2
rect 34 -2 38 2
rect 42 -2 46 2
rect 50 -2 54 2
<< nsubstratencontact >>
rect 2 78 6 82
rect 10 78 14 82
rect 18 78 22 82
rect 26 78 30 82
rect 34 78 38 82
rect 42 78 46 82
rect 50 78 54 82
<< psubstratepdiff >>
rect 0 2 56 3
rect 0 -2 2 2
rect 6 -2 10 2
rect 14 -2 18 2
rect 22 -2 26 2
rect 30 -2 34 2
rect 38 -2 42 2
rect 46 -2 50 2
rect 54 -2 56 2
rect 0 -3 56 -2
<< nsubstratendiff >>
rect 0 82 56 83
rect 0 78 2 82
rect 6 78 10 82
rect 14 78 18 82
rect 22 78 26 82
rect 30 78 34 82
rect 38 78 42 82
rect 46 78 50 82
rect 54 78 56 82
rect 0 77 56 78
<< labels >>
rlabel metal1 4 36 4 36 6 z
rlabel metal1 12 20 12 20 6 z
rlabel metal1 12 44 12 44 6 b2
rlabel metal1 28 6 28 6 6 vss
rlabel metal1 20 20 20 20 6 z
rlabel metal1 20 28 20 28 6 b1
rlabel metal1 28 28 28 28 6 b1
rlabel metal1 20 36 20 36 6 b2
rlabel polycontact 28 44 28 44 6 a2
rlabel metal1 25 57 25 57 6 n3
rlabel metal1 28 74 28 74 6 vdd
rlabel metal1 36 20 36 20 6 b1
rlabel metal1 44 32 44 32 6 a1
rlabel metal1 36 36 36 36 6 a1
rlabel metal1 44 44 44 44 6 a2
rlabel metal1 36 48 36 48 6 a2
rlabel metal1 47 56 47 56 6 n3
rlabel pdcontact 26 61 26 61 6 n3
<< end >>
