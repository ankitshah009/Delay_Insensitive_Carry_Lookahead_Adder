.subckt aoi112v0x05 a b c1 c2 vdd vss z
*   SPICE3 file   created from aoi112v0x05.ext -      technology: scmos
m00 z      c2     n2     vdd p w=28u  l=2.3636u ad=112p     pd=36u      as=125.333p ps=47.3333u
m01 n2     c1     z      vdd p w=28u  l=2.3636u ad=125.333p pd=47.3333u as=112p     ps=36u
m02 w1     b      n2     vdd p w=28u  l=2.3636u ad=84p      pd=34u      as=125.333p ps=47.3333u
m03 vdd    a      w1     vdd p w=28u  l=2.3636u ad=196p     pd=70u      as=84p      ps=34u
m04 w2     c2     z      vss n w=9u   l=2.3636u ad=22.5p    pd=14u      as=45p      ps=25.7143u
m05 vss    c1     w2     vss n w=9u   l=2.3636u ad=97.7143p pd=46.2857u as=22.5p    ps=14u
m06 z      b      vss    vss n w=6u   l=2.3636u ad=30p      pd=17.1429u as=65.1429p ps=30.8571u
m07 vss    a      z      vss n w=6u   l=2.3636u ad=65.1429p pd=30.8571u as=30p      ps=17.1429u
C0  z      vdd    0.025f
C1  a      c1     0.017f
C2  n2     c2     0.123f
C3  vss    z      0.218f
C4  b      c2     0.039f
C5  a      vdd    0.016f
C6  vss    a      0.055f
C7  c1     vdd    0.025f
C8  z      n2     0.054f
C9  vss    c1     0.017f
C10 z      b      0.051f
C11 w1     c1     0.006f
C12 w1     vdd    0.006f
C13 a      b      0.194f
C14 n2     c1     0.060f
C15 z      c2     0.245f
C16 a      c2     0.010f
C17 b      c1     0.182f
C18 n2     vdd    0.181f
C19 w2     z      0.012f
C20 c1     c2     0.107f
C21 b      vdd    0.081f
C22 vss    b      0.028f
C23 c2     vdd    0.035f
C24 z      a      0.064f
C25 vss    c2     0.014f
C26 z      c1     0.142f
C28 z      vss    0.009f
C29 a      vss    0.023f
C30 b      vss    0.027f
C31 c1     vss    0.018f
C32 c2     vss    0.022f
.ends
