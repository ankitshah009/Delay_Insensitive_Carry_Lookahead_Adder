magic
tech scmos
timestamp 1170759780
<< checkpaint >>
rect -22 -26 54 114
<< ab >>
rect 0 0 32 88
<< pwell >>
rect -4 -8 36 40
<< nwell >>
rect -4 40 36 96
<< polysilicon >>
rect 2 77 11 83
rect 9 74 11 77
rect 21 77 30 83
rect 21 74 23 77
rect 9 43 11 46
rect 21 43 23 46
rect 2 42 14 43
rect 2 38 6 42
rect 10 38 14 42
rect 2 37 14 38
rect 18 42 30 43
rect 18 38 22 42
rect 26 38 30 42
rect 18 37 30 38
rect 9 34 11 37
rect 21 34 23 37
rect 9 11 11 14
rect 2 5 11 11
rect 21 11 23 14
rect 21 5 30 11
<< ndiffusion >>
rect 2 26 9 34
rect 2 22 3 26
rect 7 22 9 26
rect 2 19 9 22
rect 2 15 3 19
rect 7 15 9 19
rect 2 14 9 15
rect 11 33 21 34
rect 11 29 14 33
rect 18 29 21 33
rect 11 25 21 29
rect 11 21 14 25
rect 18 21 21 25
rect 11 14 21 21
rect 23 26 30 34
rect 23 22 25 26
rect 29 22 30 26
rect 23 19 30 22
rect 23 15 25 19
rect 29 15 30 19
rect 23 14 30 15
rect 13 2 19 14
<< pdiffusion >>
rect 13 74 19 86
rect 2 73 9 74
rect 2 69 3 73
rect 7 69 9 73
rect 2 46 9 69
rect 11 51 21 74
rect 11 47 14 51
rect 18 47 21 51
rect 11 46 21 47
rect 23 73 30 74
rect 23 69 25 73
rect 29 69 30 73
rect 23 46 30 69
<< metal1 >>
rect -2 86 2 90
rect 10 86 22 90
rect 30 86 34 90
rect 3 82 7 86
rect 3 73 7 78
rect 3 68 7 69
rect 25 82 29 86
rect 25 73 29 78
rect 25 68 29 69
rect 6 59 26 63
rect 6 42 10 59
rect 6 33 10 38
rect 14 51 18 55
rect 14 33 18 47
rect 22 42 26 59
rect 22 33 26 38
rect 3 26 7 27
rect 3 19 7 22
rect 14 25 18 29
rect 14 17 18 21
rect 25 26 29 27
rect 25 19 29 22
rect 3 10 7 15
rect 3 2 7 6
rect 25 10 29 15
rect 25 2 29 6
rect -2 -2 2 2
rect 10 -2 22 2
rect 30 -2 34 2
<< metal2 >>
rect -2 86 6 90
rect 10 86 22 90
rect 26 86 34 90
rect -2 82 34 86
rect -2 78 3 82
rect 7 78 25 82
rect 29 78 34 82
rect -2 76 34 78
rect -2 10 34 12
rect -2 6 3 10
rect 7 6 25 10
rect 29 6 34 10
rect -2 2 34 6
rect -2 -2 6 2
rect 10 -2 22 2
rect 26 -2 34 2
<< ntransistor >>
rect 9 14 11 34
rect 21 14 23 34
<< ptransistor >>
rect 9 46 11 74
rect 21 46 23 74
<< polycontact >>
rect 6 38 10 42
rect 22 38 26 42
<< ndcontact >>
rect 3 22 7 26
rect 3 15 7 19
rect 14 29 18 33
rect 14 21 18 25
rect 25 22 29 26
rect 25 15 29 19
<< pdcontact >>
rect 3 69 7 73
rect 14 47 18 51
rect 25 69 29 73
<< m2contact >>
rect 6 86 10 90
rect 22 86 26 90
rect 3 78 7 82
rect 25 78 29 82
rect 3 6 7 10
rect 25 6 29 10
rect 6 -2 10 2
rect 22 -2 26 2
<< psubstratepcontact >>
rect 2 -2 6 2
rect 26 -2 30 2
<< nsubstratencontact >>
rect 2 86 6 90
rect 26 86 30 90
<< psubstratepdiff >>
rect 0 2 7 3
rect 25 2 32 3
rect 0 -2 2 2
rect 6 -2 7 2
rect 0 -3 7 -2
rect 25 -2 26 2
rect 30 -2 32 2
rect 25 -3 32 -2
<< nsubstratendiff >>
rect 0 90 7 91
rect 0 86 2 90
rect 6 86 7 90
rect 25 90 32 91
rect 25 86 26 90
rect 30 86 32 90
rect 0 85 7 86
rect 25 85 32 86
<< labels >>
rlabel metal1 8 48 8 48 6 a
rlabel metal1 16 36 16 36 6 z
rlabel metal1 24 48 24 48 6 a
rlabel metal2 16 6 16 6 6 vss
rlabel metal2 16 6 16 6 6 vss
rlabel metal2 16 82 16 82 6 vdd
<< end >>
