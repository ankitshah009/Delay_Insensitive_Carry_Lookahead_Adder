.subckt xor2v0x2 a b vdd vss z
*   SPICE3 file   created from xor2v0x2.ext -      technology: scmos
m00 bn     an     z      vdd p w=28u  l=2.3636u ad=112p     pd=36u      as=138.857p ps=56.5714u
m01 z      an     bn     vdd p w=28u  l=2.3636u ad=138.857p pd=56.5714u as=112p     ps=36u
m02 an     bn     z      vdd p w=21u  l=2.3636u ad=84p      pd=29u      as=104.143p ps=42.4286u
m03 z      bn     an     vdd p w=21u  l=2.3636u ad=104.143p pd=42.4286u as=84p      ps=29u
m04 bn     b      vdd    vdd p w=28u  l=2.3636u ad=112p     pd=36u      as=149.429p ps=56.5714u
m05 vdd    b      bn     vdd p w=28u  l=2.3636u ad=149.429p pd=56.5714u as=112p     ps=36u
m06 an     a      vdd    vdd p w=21u  l=2.3636u ad=84p      pd=29u      as=112.071p ps=42.4286u
m07 vdd    a      an     vdd p w=21u  l=2.3636u ad=112.071p pd=42.4286u as=84p      ps=29u
m08 w1     bn     vss    vss n w=12u  l=2.3636u ad=30p      pd=17u      as=97.8p    ps=39.2u
m09 z      an     w1     vss n w=12u  l=2.3636u ad=56.5714p pd=25.7143u as=30p      ps=17u
m10 w2     an     z      vss n w=12u  l=2.3636u ad=30p      pd=17u      as=56.5714p ps=25.7143u
m11 vss    bn     w2     vss n w=12u  l=2.3636u ad=97.8p    pd=39.2u    as=30p      ps=17u
m12 an     b      z      vss n w=18u  l=2.3636u ad=72p      pd=26u      as=84.8571p ps=38.5714u
m13 vss    a      an     vss n w=18u  l=2.3636u ad=146.7p   pd=58.8u    as=72p      ps=26u
m14 bn     b      vss    vss n w=9u   l=2.3636u ad=36p      pd=17u      as=73.35p   ps=29.4u
m15 vss    b      bn     vss n w=9u   l=2.3636u ad=73.35p   pd=29.4u    as=36p      ps=17u
C0  bn     an     0.744f
C1  vdd    an     0.135f
C2  vss    a      0.023f
C3  w2     z      0.010f
C4  vss    z      0.321f
C5  a      bn     0.243f
C6  bn     z      0.485f
C7  a      vdd    0.032f
C8  vss    b      0.071f
C9  bn     b      0.133f
C10 z      vdd    0.287f
C11 a      an     0.038f
C12 vdd    b      0.035f
C13 z      an     0.295f
C14 b      an     0.301f
C15 w1     z      0.005f
C16 vss    bn     0.252f
C17 vss    an     0.133f
C18 bn     vdd    0.438f
C19 a      b      0.136f
C21 a      vss    0.036f
C22 bn     vss    0.075f
C23 z      vss    0.016f
C25 b      vss    0.044f
C26 an     vss    0.056f
.ends
